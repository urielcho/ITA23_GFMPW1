module ita54 (clk,
    vdd,
    vss,
    segm,
    sel);
 input clk;
 input vdd;
 input vss;
 output [13:0] segm;
 output [11:0] sel;

 wire net26;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire \dut54.count[0] ;
 wire \dut54.count[1] ;
 wire \dut54.count[2] ;
 wire \dut54.count[3] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__189__CLK (.I(clknet_1_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__193__CLK (.I(clknet_1_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__195__CLK (.I(clknet_1_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__196__CLK (.I(clknet_1_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__199__CLK (.I(clknet_1_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__200__CLK (.I(clknet_1_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__201__CLK (.I(clknet_1_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__204__CLK (.I(clknet_1_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__205__CLK (.I(clknet_1_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__206__CLK (.I(clknet_1_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__207__CLK (.I(clknet_1_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__210__CLK (.I(clknet_1_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_180 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_211 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_213 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_245 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_213 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_285 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_75 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_210 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_56 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_63 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_74 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_84 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_91 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _094_ (.I(\dut54.count[2] ),
    .Z(_049_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _095_ (.I(_049_),
    .Z(_050_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _096_ (.I(\dut54.count[0] ),
    .Z(_051_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _097_ (.I(\dut54.count[1] ),
    .Z(_052_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _098_ (.I(_052_),
    .Z(_053_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _099_ (.A1(_051_),
    .A2(_053_),
    .ZN(_054_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _100_ (.I(\dut54.count[3] ),
    .ZN(_055_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _101_ (.A1(_055_),
    .A2(_049_),
    .Z(_056_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _102_ (.A1(_050_),
    .A2(_054_),
    .B(_056_),
    .ZN(_057_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _103_ (.I(\dut54.count[3] ),
    .Z(_058_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _104_ (.I(_058_),
    .Z(_059_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _105_ (.I(_059_),
    .Z(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _106_ (.I(\dut54.count[2] ),
    .ZN(_061_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _107_ (.I(_061_),
    .Z(_062_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _108_ (.A1(_059_),
    .A2(_062_),
    .ZN(_063_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _109_ (.I(\dut54.count[0] ),
    .ZN(_011_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _110_ (.A1(_011_),
    .A2(_053_),
    .Z(_064_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _111_ (.A1(net22),
    .A2(_060_),
    .B1(_063_),
    .B2(_064_),
    .ZN(_065_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _112_ (.A1(_057_),
    .A2(_065_),
    .ZN(_010_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _113_ (.A1(\dut54.count[0] ),
    .A2(\dut54.count[1] ),
    .Z(_066_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _114_ (.I(_066_),
    .Z(_012_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _115_ (.I(_054_),
    .Z(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _116_ (.A1(_050_),
    .A2(_067_),
    .ZN(_068_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _117_ (.A1(\dut54.count[3] ),
    .A2(\dut54.count[2] ),
    .ZN(_069_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _118_ (.A1(_051_),
    .A2(_052_),
    .A3(_069_),
    .ZN(_070_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _119_ (.I(_070_),
    .Z(_071_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _120_ (.A1(_068_),
    .A2(_071_),
    .ZN(_013_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _121_ (.I(_055_),
    .Z(_072_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _122_ (.A1(_072_),
    .A2(_050_),
    .ZN(_073_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _123_ (.A1(_060_),
    .A2(_054_),
    .ZN(_074_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _124_ (.A1(_073_),
    .A2(_067_),
    .B(_074_),
    .ZN(_014_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _125_ (.I(_069_),
    .Z(_075_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _126_ (.A1(_064_),
    .A2(_075_),
    .ZN(_076_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _127_ (.A1(_072_),
    .A2(_062_),
    .ZN(_077_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _128_ (.A1(_053_),
    .A2(_077_),
    .B(net18),
    .ZN(_078_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _129_ (.A1(_051_),
    .A2(_052_),
    .A3(_058_),
    .ZN(_079_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _130_ (.A1(_056_),
    .A2(_079_),
    .ZN(_080_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _131_ (.A1(\dut54.count[0] ),
    .A2(\dut54.count[1] ),
    .ZN(_081_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _132_ (.A1(_055_),
    .A2(_049_),
    .A3(_081_),
    .ZN(_082_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _133_ (.I(_082_),
    .Z(_083_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _134_ (.A1(_070_),
    .A2(_083_),
    .ZN(_084_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _135_ (.A1(_076_),
    .A2(_078_),
    .B(_080_),
    .C(_084_),
    .ZN(_015_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _136_ (.A1(_055_),
    .A2(_061_),
    .ZN(_085_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _137_ (.I(_085_),
    .Z(_086_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _138_ (.A1(net23),
    .A2(_086_),
    .ZN(_087_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _139_ (.A1(_073_),
    .A2(_067_),
    .B(_087_),
    .ZN(_016_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _140_ (.A1(_011_),
    .A2(_052_),
    .ZN(_088_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _141_ (.I(_085_),
    .Z(_089_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _142_ (.A1(_088_),
    .A2(_075_),
    .B1(_089_),
    .B2(net17),
    .ZN(_090_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _143_ (.I(_090_),
    .ZN(_017_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _144_ (.A1(_012_),
    .A2(_069_),
    .ZN(_091_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _145_ (.A1(_070_),
    .A2(_082_),
    .A3(_091_),
    .ZN(_092_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _146_ (.I(_081_),
    .Z(_093_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _147_ (.A1(_075_),
    .A2(_093_),
    .B(net14),
    .ZN(_023_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _148_ (.A1(_080_),
    .A2(_092_),
    .A3(_023_),
    .ZN(_018_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _149_ (.A1(_063_),
    .A2(_088_),
    .Z(_024_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _150_ (.A1(net8),
    .A2(_085_),
    .ZN(_025_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _151_ (.A1(_060_),
    .A2(_092_),
    .A3(_024_),
    .B(_025_),
    .ZN(_019_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _152_ (.I(net1),
    .ZN(_026_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _153_ (.I(_058_),
    .Z(_027_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _154_ (.A1(_050_),
    .A2(_064_),
    .B(_027_),
    .ZN(_028_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _155_ (.A1(_026_),
    .A2(_060_),
    .B1(_028_),
    .B2(_091_),
    .C(_057_),
    .ZN(_020_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _156_ (.A1(net7),
    .A2(_089_),
    .ZN(_029_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _157_ (.A1(_083_),
    .A2(_029_),
    .ZN(_021_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _158_ (.A1(net9),
    .A2(_079_),
    .B(_077_),
    .ZN(_030_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _159_ (.A1(_071_),
    .A2(_030_),
    .B(_080_),
    .ZN(_022_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _160_ (.A1(net6),
    .A2(_089_),
    .ZN(_031_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _161_ (.A1(_071_),
    .A2(_031_),
    .ZN(_000_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _162_ (.A1(_072_),
    .A2(_049_),
    .ZN(_032_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _163_ (.A1(_032_),
    .A2(_064_),
    .B1(_086_),
    .B2(net15),
    .ZN(_033_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _164_ (.I(_033_),
    .ZN(_001_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _165_ (.A1(_058_),
    .A2(_061_),
    .ZN(_034_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _166_ (.A1(net16),
    .A2(_086_),
    .ZN(_035_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _167_ (.A1(_034_),
    .A2(_067_),
    .B(_035_),
    .ZN(_002_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _168_ (.A1(_059_),
    .A2(_062_),
    .A3(_081_),
    .ZN(_036_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _169_ (.A1(net10),
    .A2(_089_),
    .ZN(_037_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _170_ (.A1(_036_),
    .A2(_037_),
    .ZN(_003_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _171_ (.A1(net11),
    .A2(_027_),
    .B1(_088_),
    .B2(_075_),
    .ZN(_038_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _172_ (.A1(_034_),
    .A2(_093_),
    .ZN(_039_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _173_ (.A1(_036_),
    .A2(_038_),
    .B(_039_),
    .ZN(_004_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _174_ (.A1(_070_),
    .A2(_083_),
    .A3(_091_),
    .Z(_040_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _175_ (.A1(net13),
    .A2(_027_),
    .B1(_032_),
    .B2(_093_),
    .ZN(_041_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _176_ (.A1(_040_),
    .A2(_041_),
    .B(_039_),
    .ZN(_005_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _177_ (.A1(net3),
    .A2(_059_),
    .ZN(_042_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _178_ (.A1(_071_),
    .A2(_083_),
    .A3(_036_),
    .A4(_042_),
    .Z(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _179_ (.A1(_039_),
    .A2(_043_),
    .ZN(_006_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _180_ (.A1(_062_),
    .A2(_093_),
    .B(net4),
    .C(_072_),
    .ZN(_044_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _181_ (.A1(_084_),
    .A2(_024_),
    .A3(_039_),
    .A4(_044_),
    .ZN(_045_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _182_ (.I(_045_),
    .Z(_007_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _183_ (.A1(_063_),
    .A2(_088_),
    .B1(_086_),
    .B2(net21),
    .ZN(_046_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _184_ (.I(_046_),
    .ZN(_008_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _185_ (.A1(net25),
    .A2(_027_),
    .A3(_036_),
    .ZN(_047_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _186_ (.A1(_051_),
    .A2(_032_),
    .ZN(_048_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _187_ (.A1(_053_),
    .A2(_032_),
    .B1(_047_),
    .B2(_048_),
    .ZN(_009_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _188_ (.D(_010_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net22),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _189_ (.D(_011_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\dut54.count[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _190_ (.D(_012_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\dut54.count[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _191_ (.D(_013_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\dut54.count[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _192_ (.D(_014_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\dut54.count[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _193_ (.D(_015_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net18),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _194_ (.D(_016_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net23),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _195_ (.D(_017_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net17),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _196_ (.D(_018_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net14),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _197_ (.D(_019_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net8),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _198_ (.D(_020_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _199_ (.D(_021_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net7),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _200_ (.D(_022_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net9),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _201_ (.D(_000_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net6),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _202_ (.D(_001_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net15),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _203_ (.D(_002_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net16),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _204_ (.D(_003_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net10),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _205_ (.D(_004_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net11),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _206_ (.D(_005_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net13),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _207_ (.D(_006_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _208_ (.D(_007_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _209_ (.D(_008_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net21),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _210_ (.D(_009_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net25),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _212_ (.I(net8),
    .Z(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _213_ (.I(net13),
    .Z(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _214_ (.I(net3),
    .Z(net2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _215_ (.I(net6),
    .Z(net19),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _216_ (.I(net7),
    .Z(net20),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _217_ (.I(net10),
    .Z(net24),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita54_26 (.ZN(net26),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1 (.I(net1),
    .Z(segm[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output10 (.I(net10),
    .Z(segm[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output11 (.I(net11),
    .Z(segm[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output12 (.I(net12),
    .Z(segm[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output13 (.I(net13),
    .Z(segm[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output14 (.I(net14),
    .Z(sel[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output15 (.I(net15),
    .Z(sel[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output16 (.I(net16),
    .Z(sel[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output17 (.I(net17),
    .Z(sel[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output18 (.I(net18),
    .Z(sel[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output19 (.I(net19),
    .Z(sel[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output2 (.I(net2),
    .Z(segm[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output20 (.I(net20),
    .Z(sel[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output21 (.I(net21),
    .Z(sel[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output22 (.I(net22),
    .Z(sel[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output23 (.I(net23),
    .Z(sel[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output24 (.I(net24),
    .Z(sel[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output25 (.I(net25),
    .Z(sel[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output3 (.I(net3),
    .Z(segm[12]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output4 (.I(net4),
    .Z(segm[13]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output5 (.I(net5),
    .Z(segm[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output6 (.I(net6),
    .Z(segm[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output7 (.I(net7),
    .Z(segm[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output8 (.I(net8),
    .Z(segm[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output9 (.I(net9),
    .Z(segm[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 assign segm[0] = net26;
endmodule
