magic
tech gf180mcuD
magscale 1 5
timestamp 1699642671
<< obsm1 >>
rect 672 1538 20328 19238
<< metal2 >>
rect 11424 20600 11480 21000
rect 12432 20600 12488 21000
rect 8400 0 8456 400
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 10080 0 10136 400
rect 10416 0 10472 400
rect 10752 0 10808 400
rect 11088 0 11144 400
rect 11424 0 11480 400
rect 11760 0 11816 400
rect 12432 0 12488 400
rect 12768 0 12824 400
<< obsm2 >>
rect 854 20570 11394 20600
rect 11510 20570 12402 20600
rect 12518 20570 20146 20600
rect 854 430 20146 20570
rect 854 400 8370 430
rect 8486 400 8706 430
rect 8822 400 9042 430
rect 9158 400 10050 430
rect 10166 400 10386 430
rect 10502 400 10722 430
rect 10838 400 11058 430
rect 11174 400 11394 430
rect 11510 400 11730 430
rect 11846 400 12402 430
rect 12518 400 12738 430
rect 12854 400 20146 430
<< metal3 >>
rect 0 18144 400 18200
rect 20600 18144 21000 18200
rect 20600 17808 21000 17864
rect 0 13104 400 13160
rect 0 12432 400 12488
rect 20600 12432 21000 12488
rect 0 12096 400 12152
rect 0 11424 400 11480
rect 20600 11424 21000 11480
rect 0 10416 400 10472
rect 20600 10416 21000 10472
rect 20600 9744 21000 9800
rect 20600 9072 21000 9128
rect 0 8736 400 8792
<< obsm3 >>
rect 400 18230 20600 19222
rect 430 18114 20570 18230
rect 400 17894 20600 18114
rect 400 17778 20570 17894
rect 400 13190 20600 17778
rect 430 13074 20600 13190
rect 400 12518 20600 13074
rect 430 12402 20570 12518
rect 400 12182 20600 12402
rect 430 12066 20600 12182
rect 400 11510 20600 12066
rect 430 11394 20570 11510
rect 400 10502 20600 11394
rect 430 10386 20570 10502
rect 400 9830 20600 10386
rect 400 9714 20570 9830
rect 400 9158 20600 9714
rect 400 9042 20570 9158
rect 400 8822 20600 9042
rect 430 8706 20600 8822
rect 400 1554 20600 8706
<< metal4 >>
rect 2224 1538 2384 19238
rect 9904 1538 10064 19238
rect 17584 1538 17744 19238
<< obsm4 >>
rect 10374 8241 10402 8503
<< labels >>
rlabel metal3 s 0 13104 400 13160 6 clk
port 1 nsew signal input
rlabel metal3 s 20600 18144 21000 18200 6 segm[0]
port 2 nsew signal output
rlabel metal2 s 8400 0 8456 400 6 segm[10]
port 3 nsew signal output
rlabel metal2 s 11760 0 11816 400 6 segm[11]
port 4 nsew signal output
rlabel metal2 s 11088 0 11144 400 6 segm[12]
port 5 nsew signal output
rlabel metal2 s 10416 0 10472 400 6 segm[13]
port 6 nsew signal output
rlabel metal2 s 10752 0 10808 400 6 segm[1]
port 7 nsew signal output
rlabel metal3 s 20600 17808 21000 17864 6 segm[2]
port 8 nsew signal output
rlabel metal2 s 12432 0 12488 400 6 segm[3]
port 9 nsew signal output
rlabel metal3 s 0 18144 400 18200 6 segm[4]
port 10 nsew signal output
rlabel metal2 s 11424 0 11480 400 6 segm[5]
port 11 nsew signal output
rlabel metal3 s 0 12432 400 12488 6 segm[6]
port 12 nsew signal output
rlabel metal3 s 0 12096 400 12152 6 segm[7]
port 13 nsew signal output
rlabel metal2 s 9072 0 9128 400 6 segm[8]
port 14 nsew signal output
rlabel metal2 s 8736 0 8792 400 6 segm[9]
port 15 nsew signal output
rlabel metal3 s 20600 12432 21000 12488 6 sel[0]
port 16 nsew signal output
rlabel metal3 s 20600 9744 21000 9800 6 sel[10]
port 17 nsew signal output
rlabel metal3 s 20600 10416 21000 10472 6 sel[11]
port 18 nsew signal output
rlabel metal3 s 0 11424 400 11480 6 sel[1]
port 19 nsew signal output
rlabel metal2 s 12768 0 12824 400 6 sel[2]
port 20 nsew signal output
rlabel metal2 s 11424 20600 11480 21000 6 sel[3]
port 21 nsew signal output
rlabel metal2 s 10080 0 10136 400 6 sel[4]
port 22 nsew signal output
rlabel metal3 s 0 10416 400 10472 6 sel[5]
port 23 nsew signal output
rlabel metal3 s 0 8736 400 8792 6 sel[6]
port 24 nsew signal output
rlabel metal2 s 12432 20600 12488 21000 6 sel[7]
port 25 nsew signal output
rlabel metal3 s 20600 9072 21000 9128 6 sel[8]
port 26 nsew signal output
rlabel metal3 s 20600 11424 21000 11480 6 sel[9]
port 27 nsew signal output
rlabel metal4 s 2224 1538 2384 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 19238 6 vss
port 29 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 21000 21000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 450232
string GDS_FILE /home/urielcho/Proyectos_caravel/ITA23_GFMPW1b/openlane/ita45/runs/23_11_10_12_55/results/signoff/ita45.magic.gds
string GDS_START 152716
<< end >>

