magic
tech gf180mcuD
magscale 1 10
timestamp 1699642983
<< metal1 >>
rect 18834 38558 18846 38610
rect 18898 38607 18910 38610
rect 19954 38607 19966 38610
rect 18898 38561 19966 38607
rect 18898 38558 18910 38561
rect 19954 38558 19966 38561
rect 20018 38558 20030 38610
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 18062 38274 18114 38286
rect 18062 38210 18114 38222
rect 22430 38274 22482 38286
rect 22430 38210 22482 38222
rect 26126 38274 26178 38286
rect 26126 38210 26178 38222
rect 29374 38274 29426 38286
rect 29374 38210 29426 38222
rect 17042 37998 17054 38050
rect 17106 37998 17118 38050
rect 21410 37998 21422 38050
rect 21474 37998 21486 38050
rect 25218 37998 25230 38050
rect 25282 37998 25294 38050
rect 28578 37998 28590 38050
rect 28642 37998 28654 38050
rect 19966 37938 20018 37950
rect 19966 37874 20018 37886
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 18398 37490 18450 37502
rect 18398 37426 18450 37438
rect 21422 37490 21474 37502
rect 21422 37426 21474 37438
rect 17378 37214 17390 37266
rect 17442 37214 17454 37266
rect 20402 37214 20414 37266
rect 20466 37214 20478 37266
rect 28242 37214 28254 37266
rect 28306 37214 28318 37266
rect 26014 37154 26066 37166
rect 26014 37090 26066 37102
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 1710 36370 1762 36382
rect 1710 36306 1762 36318
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 15710 28642 15762 28654
rect 15710 28578 15762 28590
rect 15822 28642 15874 28654
rect 15822 28578 15874 28590
rect 16158 28642 16210 28654
rect 16158 28578 16210 28590
rect 16382 28642 16434 28654
rect 16382 28578 16434 28590
rect 17278 28642 17330 28654
rect 17278 28578 17330 28590
rect 16718 28530 16770 28542
rect 16718 28466 16770 28478
rect 19518 28530 19570 28542
rect 19518 28466 19570 28478
rect 19630 28530 19682 28542
rect 19630 28466 19682 28478
rect 20526 28530 20578 28542
rect 20526 28466 20578 28478
rect 20638 28530 20690 28542
rect 20638 28466 20690 28478
rect 15934 28418 15986 28430
rect 15934 28354 15986 28366
rect 16606 28418 16658 28430
rect 16606 28354 16658 28366
rect 19294 28418 19346 28430
rect 19294 28354 19346 28366
rect 20862 28418 20914 28430
rect 20862 28354 20914 28366
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 18846 27970 18898 27982
rect 14578 27918 14590 27970
rect 14642 27918 14654 27970
rect 18846 27906 18898 27918
rect 18958 27970 19010 27982
rect 18958 27906 19010 27918
rect 18622 27858 18674 27870
rect 13794 27806 13806 27858
rect 13858 27806 13870 27858
rect 22194 27806 22206 27858
rect 22258 27806 22270 27858
rect 18622 27794 18674 27806
rect 17614 27746 17666 27758
rect 22766 27746 22818 27758
rect 16706 27694 16718 27746
rect 16770 27694 16782 27746
rect 19282 27694 19294 27746
rect 19346 27694 19358 27746
rect 21410 27694 21422 27746
rect 21474 27694 21486 27746
rect 17614 27682 17666 27694
rect 22766 27682 22818 27694
rect 25454 27746 25506 27758
rect 25454 27682 25506 27694
rect 25902 27746 25954 27758
rect 25902 27682 25954 27694
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 21422 27298 21474 27310
rect 21422 27234 21474 27246
rect 16370 27134 16382 27186
rect 16434 27134 16446 27186
rect 18162 27134 18174 27186
rect 18226 27134 18238 27186
rect 20290 27134 20302 27186
rect 20354 27134 20366 27186
rect 24994 27134 25006 27186
rect 25058 27134 25070 27186
rect 28242 27134 28254 27186
rect 28306 27134 28318 27186
rect 16606 27074 16658 27086
rect 13570 27022 13582 27074
rect 13634 27022 13646 27074
rect 16606 27010 16658 27022
rect 16942 27074 16994 27086
rect 21310 27074 21362 27086
rect 17490 27022 17502 27074
rect 17554 27022 17566 27074
rect 22194 27022 22206 27074
rect 22258 27022 22270 27074
rect 25442 27022 25454 27074
rect 25506 27022 25518 27074
rect 16942 27010 16994 27022
rect 21310 27010 21362 27022
rect 16830 26962 16882 26974
rect 14242 26910 14254 26962
rect 14306 26910 14318 26962
rect 16830 26898 16882 26910
rect 20750 26962 20802 26974
rect 22866 26910 22878 26962
rect 22930 26910 22942 26962
rect 26114 26910 26126 26962
rect 26178 26910 26190 26962
rect 20750 26898 20802 26910
rect 21422 26850 21474 26862
rect 21422 26786 21474 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 14814 26514 14866 26526
rect 14814 26450 14866 26462
rect 16606 26514 16658 26526
rect 21870 26514 21922 26526
rect 17602 26462 17614 26514
rect 17666 26462 17678 26514
rect 16606 26450 16658 26462
rect 21870 26450 21922 26462
rect 23102 26514 23154 26526
rect 26450 26462 26462 26514
rect 26514 26462 26526 26514
rect 23102 26450 23154 26462
rect 14926 26402 14978 26414
rect 14926 26338 14978 26350
rect 24222 26402 24274 26414
rect 24222 26338 24274 26350
rect 25566 26402 25618 26414
rect 25566 26338 25618 26350
rect 17950 26290 18002 26302
rect 22990 26290 23042 26302
rect 18610 26238 18622 26290
rect 18674 26238 18686 26290
rect 17950 26226 18002 26238
rect 22990 26226 23042 26238
rect 23214 26290 23266 26302
rect 23214 26226 23266 26238
rect 23550 26290 23602 26302
rect 23550 26226 23602 26238
rect 23886 26290 23938 26302
rect 23886 26226 23938 26238
rect 23998 26290 24050 26302
rect 23998 26226 24050 26238
rect 24446 26290 24498 26302
rect 24446 26226 24498 26238
rect 25118 26290 25170 26302
rect 25118 26226 25170 26238
rect 25678 26290 25730 26302
rect 26226 26238 26238 26290
rect 26290 26238 26302 26290
rect 25678 26226 25730 26238
rect 25342 26178 25394 26190
rect 19282 26126 19294 26178
rect 19346 26126 19358 26178
rect 21410 26126 21422 26178
rect 21474 26126 21486 26178
rect 25342 26114 25394 26126
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 24894 25730 24946 25742
rect 24894 25666 24946 25678
rect 24782 25618 24834 25630
rect 24782 25554 24834 25566
rect 24546 25454 24558 25506
rect 24610 25454 24622 25506
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 19406 24946 19458 24958
rect 19406 24882 19458 24894
rect 19742 24946 19794 24958
rect 19742 24882 19794 24894
rect 20078 24946 20130 24958
rect 20078 24882 20130 24894
rect 21982 24946 22034 24958
rect 21982 24882 22034 24894
rect 20302 24834 20354 24846
rect 20302 24770 20354 24782
rect 14366 24722 14418 24734
rect 4274 24670 4286 24722
rect 4338 24670 4350 24722
rect 13794 24670 13806 24722
rect 13858 24670 13870 24722
rect 14366 24658 14418 24670
rect 17390 24722 17442 24734
rect 17390 24658 17442 24670
rect 17614 24722 17666 24734
rect 17614 24658 17666 24670
rect 17838 24722 17890 24734
rect 17838 24658 17890 24670
rect 19294 24722 19346 24734
rect 19294 24658 19346 24670
rect 19518 24722 19570 24734
rect 19518 24658 19570 24670
rect 20414 24722 20466 24734
rect 20414 24658 20466 24670
rect 21422 24722 21474 24734
rect 21422 24658 21474 24670
rect 17502 24610 17554 24622
rect 10994 24558 11006 24610
rect 11058 24558 11070 24610
rect 13122 24558 13134 24610
rect 13186 24558 13198 24610
rect 17502 24546 17554 24558
rect 1934 24498 1986 24510
rect 1934 24434 1986 24446
rect 21646 24498 21698 24510
rect 21646 24434 21698 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 12798 24162 12850 24174
rect 12798 24098 12850 24110
rect 1934 24050 1986 24062
rect 18510 24050 18562 24062
rect 40014 24050 40066 24062
rect 15922 23998 15934 24050
rect 15986 23998 15998 24050
rect 18050 23998 18062 24050
rect 18114 23998 18126 24050
rect 19842 23998 19854 24050
rect 19906 23998 19918 24050
rect 28578 23998 28590 24050
rect 28642 23998 28654 24050
rect 1934 23986 1986 23998
rect 18510 23986 18562 23998
rect 40014 23986 40066 23998
rect 12910 23938 12962 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 12910 23874 12962 23886
rect 14030 23938 14082 23950
rect 15138 23886 15150 23938
rect 15202 23886 15214 23938
rect 20290 23886 20302 23938
rect 20354 23886 20366 23938
rect 21298 23886 21310 23938
rect 21362 23886 21374 23938
rect 25666 23886 25678 23938
rect 25730 23886 25742 23938
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 14030 23874 14082 23886
rect 12798 23826 12850 23838
rect 12798 23762 12850 23774
rect 13470 23826 13522 23838
rect 13470 23762 13522 23774
rect 13582 23826 13634 23838
rect 13582 23762 13634 23774
rect 14366 23826 14418 23838
rect 14366 23762 14418 23774
rect 14590 23826 14642 23838
rect 14590 23762 14642 23774
rect 19518 23826 19570 23838
rect 19518 23762 19570 23774
rect 19742 23826 19794 23838
rect 21634 23774 21646 23826
rect 21698 23774 21710 23826
rect 22194 23774 22206 23826
rect 22258 23774 22270 23826
rect 26450 23774 26462 23826
rect 26514 23774 26526 23826
rect 19742 23762 19794 23774
rect 13806 23714 13858 23726
rect 13806 23650 13858 23662
rect 14142 23714 14194 23726
rect 19182 23714 19234 23726
rect 25342 23714 25394 23726
rect 18834 23662 18846 23714
rect 18898 23662 18910 23714
rect 20514 23662 20526 23714
rect 20578 23662 20590 23714
rect 21858 23662 21870 23714
rect 21922 23662 21934 23714
rect 14142 23650 14194 23662
rect 19182 23650 19234 23662
rect 25342 23650 25394 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 14590 23378 14642 23390
rect 14590 23314 14642 23326
rect 14814 23378 14866 23390
rect 26462 23378 26514 23390
rect 15810 23326 15822 23378
rect 15874 23326 15886 23378
rect 14814 23314 14866 23326
rect 26462 23314 26514 23326
rect 27022 23378 27074 23390
rect 27022 23314 27074 23326
rect 25454 23266 25506 23278
rect 13122 23214 13134 23266
rect 13186 23214 13198 23266
rect 22082 23214 22094 23266
rect 22146 23214 22158 23266
rect 25454 23202 25506 23214
rect 14366 23154 14418 23166
rect 13794 23102 13806 23154
rect 13858 23102 13870 23154
rect 14366 23090 14418 23102
rect 14478 23154 14530 23166
rect 14478 23090 14530 23102
rect 14702 23154 14754 23166
rect 14702 23090 14754 23102
rect 16158 23154 16210 23166
rect 16158 23090 16210 23102
rect 16382 23154 16434 23166
rect 25342 23154 25394 23166
rect 18274 23102 18286 23154
rect 18338 23102 18350 23154
rect 20066 23102 20078 23154
rect 20130 23102 20142 23154
rect 16382 23090 16434 23102
rect 25342 23090 25394 23102
rect 25678 23154 25730 23166
rect 25678 23090 25730 23102
rect 26014 23154 26066 23166
rect 26014 23090 26066 23102
rect 26238 23154 26290 23166
rect 26238 23090 26290 23102
rect 26686 23154 26738 23166
rect 26686 23090 26738 23102
rect 26910 23154 26962 23166
rect 26910 23090 26962 23102
rect 17950 23042 18002 23054
rect 10994 22990 11006 23042
rect 11058 22990 11070 23042
rect 17950 22978 18002 22990
rect 18846 23042 18898 23054
rect 18846 22978 18898 22990
rect 17726 22930 17778 22942
rect 17378 22878 17390 22930
rect 17442 22878 17454 22930
rect 17726 22866 17778 22878
rect 18622 22930 18674 22942
rect 18622 22866 18674 22878
rect 27022 22930 27074 22942
rect 27022 22866 27074 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 14142 22482 14194 22494
rect 14142 22418 14194 22430
rect 20414 22482 20466 22494
rect 40014 22482 40066 22494
rect 21746 22430 21758 22482
rect 21810 22430 21822 22482
rect 28242 22430 28254 22482
rect 28306 22430 28318 22482
rect 20414 22418 20466 22430
rect 40014 22418 40066 22430
rect 20190 22370 20242 22382
rect 23886 22370 23938 22382
rect 18610 22318 18622 22370
rect 18674 22318 18686 22370
rect 22082 22318 22094 22370
rect 22146 22318 22158 22370
rect 25330 22318 25342 22370
rect 25394 22318 25406 22370
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 20190 22306 20242 22318
rect 23886 22306 23938 22318
rect 18062 22258 18114 22270
rect 21310 22258 21362 22270
rect 19506 22206 19518 22258
rect 19570 22206 19582 22258
rect 20066 22206 20078 22258
rect 20130 22206 20142 22258
rect 18062 22194 18114 22206
rect 21310 22194 21362 22206
rect 23102 22258 23154 22270
rect 26114 22206 26126 22258
rect 26178 22206 26190 22258
rect 23102 22194 23154 22206
rect 18174 22146 18226 22158
rect 21534 22146 21586 22158
rect 18834 22094 18846 22146
rect 18898 22094 18910 22146
rect 18174 22082 18226 22094
rect 21534 22082 21586 22094
rect 21758 22146 21810 22158
rect 21758 22082 21810 22094
rect 22206 22146 22258 22158
rect 22206 22082 22258 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 19966 21810 20018 21822
rect 21634 21758 21646 21810
rect 21698 21758 21710 21810
rect 23762 21758 23774 21810
rect 23826 21758 23838 21810
rect 19966 21746 20018 21758
rect 25678 21698 25730 21710
rect 17714 21646 17726 21698
rect 17778 21646 17790 21698
rect 18610 21646 18622 21698
rect 18674 21646 18686 21698
rect 19506 21646 19518 21698
rect 19570 21646 19582 21698
rect 20962 21646 20974 21698
rect 21026 21646 21038 21698
rect 21746 21646 21758 21698
rect 21810 21646 21822 21698
rect 22978 21646 22990 21698
rect 23042 21646 23054 21698
rect 23538 21646 23550 21698
rect 23602 21646 23614 21698
rect 24658 21646 24670 21698
rect 24722 21646 24734 21698
rect 25678 21634 25730 21646
rect 25902 21698 25954 21710
rect 25902 21634 25954 21646
rect 26238 21698 26290 21710
rect 26238 21634 26290 21646
rect 24334 21586 24386 21598
rect 17490 21534 17502 21586
rect 17554 21534 17566 21586
rect 18386 21534 18398 21586
rect 18450 21534 18462 21586
rect 19394 21534 19406 21586
rect 19458 21534 19470 21586
rect 20850 21534 20862 21586
rect 20914 21534 20926 21586
rect 22866 21534 22878 21586
rect 22930 21534 22942 21586
rect 24334 21522 24386 21534
rect 25342 21586 25394 21598
rect 25342 21522 25394 21534
rect 25454 21586 25506 21598
rect 25454 21522 25506 21534
rect 26350 21586 26402 21598
rect 28142 21586 28194 21598
rect 27682 21534 27694 21586
rect 27746 21534 27758 21586
rect 28354 21534 28366 21586
rect 28418 21534 28430 21586
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 26350 21522 26402 21534
rect 28142 21522 28194 21534
rect 20526 21474 20578 21486
rect 20526 21410 20578 21422
rect 25566 21474 25618 21486
rect 25566 21410 25618 21422
rect 26686 21474 26738 21486
rect 26686 21410 26738 21422
rect 19518 21362 19570 21374
rect 19518 21298 19570 21310
rect 26574 21362 26626 21374
rect 26574 21298 26626 21310
rect 27134 21362 27186 21374
rect 27134 21298 27186 21310
rect 27246 21362 27298 21374
rect 27246 21298 27298 21310
rect 27470 21362 27522 21374
rect 27470 21298 27522 21310
rect 28030 21362 28082 21374
rect 28030 21298 28082 21310
rect 40014 21362 40066 21374
rect 40014 21298 40066 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 18846 21026 18898 21038
rect 18846 20962 18898 20974
rect 19182 21026 19234 21038
rect 19182 20962 19234 20974
rect 17054 20914 17106 20926
rect 23326 20914 23378 20926
rect 20178 20862 20190 20914
rect 20242 20862 20254 20914
rect 17054 20850 17106 20862
rect 23326 20850 23378 20862
rect 25342 20914 25394 20926
rect 26450 20862 26462 20914
rect 26514 20862 26526 20914
rect 28578 20862 28590 20914
rect 28642 20862 28654 20914
rect 25342 20850 25394 20862
rect 14814 20802 14866 20814
rect 16494 20802 16546 20814
rect 15026 20750 15038 20802
rect 15090 20750 15102 20802
rect 14814 20738 14866 20750
rect 16494 20738 16546 20750
rect 17390 20802 17442 20814
rect 17390 20738 17442 20750
rect 17950 20802 18002 20814
rect 17950 20738 18002 20750
rect 18174 20802 18226 20814
rect 21758 20802 21810 20814
rect 24558 20802 24610 20814
rect 19282 20750 19294 20802
rect 19346 20750 19358 20802
rect 19842 20750 19854 20802
rect 19906 20750 19918 20802
rect 22194 20750 22206 20802
rect 22258 20750 22270 20802
rect 23090 20750 23102 20802
rect 23154 20750 23166 20802
rect 23650 20750 23662 20802
rect 23714 20750 23726 20802
rect 24210 20750 24222 20802
rect 24274 20750 24286 20802
rect 25666 20750 25678 20802
rect 25730 20750 25742 20802
rect 18174 20738 18226 20750
rect 21758 20738 21810 20750
rect 24558 20738 24610 20750
rect 15710 20690 15762 20702
rect 22754 20638 22766 20690
rect 22818 20638 22830 20690
rect 24882 20638 24894 20690
rect 24946 20638 24958 20690
rect 15710 20626 15762 20638
rect 18510 20578 18562 20590
rect 18510 20514 18562 20526
rect 18734 20578 18786 20590
rect 18734 20514 18786 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 24558 20242 24610 20254
rect 24558 20178 24610 20190
rect 24782 20242 24834 20254
rect 24782 20178 24834 20190
rect 26014 20242 26066 20254
rect 26014 20178 26066 20190
rect 15710 20130 15762 20142
rect 15710 20066 15762 20078
rect 17390 20130 17442 20142
rect 17390 20066 17442 20078
rect 24446 20130 24498 20142
rect 24446 20066 24498 20078
rect 25230 20130 25282 20142
rect 25230 20066 25282 20078
rect 18510 20018 18562 20030
rect 12114 19966 12126 20018
rect 12178 19966 12190 20018
rect 15474 19966 15486 20018
rect 15538 19966 15550 20018
rect 19730 19966 19742 20018
rect 19794 19966 19806 20018
rect 18510 19954 18562 19966
rect 16270 19906 16322 19918
rect 12898 19854 12910 19906
rect 12962 19854 12974 19906
rect 15026 19854 15038 19906
rect 15090 19854 15102 19906
rect 16270 19842 16322 19854
rect 17950 19906 18002 19918
rect 22306 19854 22318 19906
rect 22370 19854 22382 19906
rect 25442 19854 25454 19906
rect 25506 19854 25518 19906
rect 17950 19842 18002 19854
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 15262 19458 15314 19470
rect 15262 19394 15314 19406
rect 27246 19458 27298 19470
rect 27246 19394 27298 19406
rect 15486 19346 15538 19358
rect 15486 19282 15538 19294
rect 18622 19346 18674 19358
rect 18622 19282 18674 19294
rect 19294 19346 19346 19358
rect 20290 19294 20302 19346
rect 20354 19294 20366 19346
rect 24658 19294 24670 19346
rect 24722 19294 24734 19346
rect 19294 19282 19346 19294
rect 18734 19234 18786 19246
rect 19406 19234 19458 19246
rect 26574 19234 26626 19246
rect 27358 19234 27410 19246
rect 17266 19182 17278 19234
rect 17330 19182 17342 19234
rect 17938 19182 17950 19234
rect 18002 19182 18014 19234
rect 18386 19182 18398 19234
rect 18450 19182 18462 19234
rect 19058 19182 19070 19234
rect 19122 19182 19134 19234
rect 23538 19182 23550 19234
rect 23602 19182 23614 19234
rect 23986 19182 23998 19234
rect 24050 19182 24062 19234
rect 26338 19182 26350 19234
rect 26402 19182 26414 19234
rect 26898 19182 26910 19234
rect 26962 19182 26974 19234
rect 27570 19182 27582 19234
rect 27634 19182 27646 19234
rect 18734 19170 18786 19182
rect 19406 19170 19458 19182
rect 26574 19170 26626 19182
rect 27358 19170 27410 19182
rect 23102 19122 23154 19134
rect 17042 19070 17054 19122
rect 17106 19070 17118 19122
rect 17714 19070 17726 19122
rect 17778 19070 17790 19122
rect 23102 19058 23154 19070
rect 24558 19122 24610 19134
rect 24558 19058 24610 19070
rect 26126 19122 26178 19134
rect 26126 19058 26178 19070
rect 20750 19010 20802 19022
rect 14914 18958 14926 19010
rect 14978 18958 14990 19010
rect 20750 18946 20802 18958
rect 26238 19010 26290 19022
rect 26238 18946 26290 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 21086 18674 21138 18686
rect 21086 18610 21138 18622
rect 17726 18562 17778 18574
rect 17726 18498 17778 18510
rect 17838 18562 17890 18574
rect 18162 18510 18174 18562
rect 18226 18510 18238 18562
rect 19506 18510 19518 18562
rect 19570 18510 19582 18562
rect 22418 18510 22430 18562
rect 22482 18510 22494 18562
rect 22978 18510 22990 18562
rect 23042 18510 23054 18562
rect 26338 18510 26350 18562
rect 26402 18510 26414 18562
rect 17838 18498 17890 18510
rect 18510 18450 18562 18462
rect 19854 18450 19906 18462
rect 21198 18450 21250 18462
rect 11666 18398 11678 18450
rect 11730 18398 11742 18450
rect 19170 18398 19182 18450
rect 19234 18398 19246 18450
rect 20290 18398 20302 18450
rect 20354 18398 20366 18450
rect 18510 18386 18562 18398
rect 19854 18386 19906 18398
rect 21198 18386 21250 18398
rect 21758 18450 21810 18462
rect 21758 18386 21810 18398
rect 23102 18450 23154 18462
rect 23102 18386 23154 18398
rect 24110 18450 24162 18462
rect 24110 18386 24162 18398
rect 24446 18450 24498 18462
rect 25554 18398 25566 18450
rect 25618 18398 25630 18450
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 24446 18386 24498 18398
rect 14926 18338 14978 18350
rect 12338 18286 12350 18338
rect 12402 18286 12414 18338
rect 14466 18286 14478 18338
rect 14530 18286 14542 18338
rect 14926 18274 14978 18286
rect 20750 18338 20802 18350
rect 20750 18274 20802 18286
rect 23326 18338 23378 18350
rect 28466 18286 28478 18338
rect 28530 18286 28542 18338
rect 23326 18274 23378 18286
rect 17726 18226 17778 18238
rect 17726 18162 17778 18174
rect 18846 18226 18898 18238
rect 18846 18162 18898 18174
rect 19182 18226 19234 18238
rect 19182 18162 19234 18174
rect 23886 18226 23938 18238
rect 23886 18162 23938 18174
rect 24558 18226 24610 18238
rect 24558 18162 24610 18174
rect 24670 18226 24722 18238
rect 24670 18162 24722 18174
rect 40014 18226 40066 18238
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 14478 17890 14530 17902
rect 14478 17826 14530 17838
rect 1934 17778 1986 17790
rect 18510 17778 18562 17790
rect 9986 17726 9998 17778
rect 10050 17726 10062 17778
rect 1934 17714 1986 17726
rect 18510 17714 18562 17726
rect 40014 17778 40066 17790
rect 40014 17714 40066 17726
rect 13582 17666 13634 17678
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 12786 17614 12798 17666
rect 12850 17614 12862 17666
rect 13582 17602 13634 17614
rect 14254 17666 14306 17678
rect 14254 17602 14306 17614
rect 14814 17666 14866 17678
rect 14814 17602 14866 17614
rect 17390 17666 17442 17678
rect 17390 17602 17442 17614
rect 17726 17666 17778 17678
rect 17726 17602 17778 17614
rect 17950 17666 18002 17678
rect 17950 17602 18002 17614
rect 18398 17666 18450 17678
rect 19518 17666 19570 17678
rect 18946 17614 18958 17666
rect 19010 17614 19022 17666
rect 19730 17614 19742 17666
rect 19794 17614 19806 17666
rect 23314 17614 23326 17666
rect 23378 17614 23390 17666
rect 23762 17614 23774 17666
rect 23826 17614 23838 17666
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 18398 17602 18450 17614
rect 19518 17602 19570 17614
rect 15038 17554 15090 17566
rect 12114 17502 12126 17554
rect 12178 17502 12190 17554
rect 15038 17490 15090 17502
rect 17166 17554 17218 17566
rect 17166 17490 17218 17502
rect 17502 17554 17554 17566
rect 17502 17490 17554 17502
rect 18622 17554 18674 17566
rect 24334 17554 24386 17566
rect 21858 17502 21870 17554
rect 21922 17502 21934 17554
rect 18622 17490 18674 17502
rect 24334 17490 24386 17502
rect 25902 17554 25954 17566
rect 25902 17490 25954 17502
rect 14142 17442 14194 17454
rect 14142 17378 14194 17390
rect 15486 17442 15538 17454
rect 15486 17378 15538 17390
rect 19630 17442 19682 17454
rect 19630 17378 19682 17390
rect 25006 17442 25058 17454
rect 25006 17378 25058 17390
rect 26238 17442 26290 17454
rect 26238 17378 26290 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 16494 17106 16546 17118
rect 16494 17042 16546 17054
rect 16830 17106 16882 17118
rect 16830 17042 16882 17054
rect 23886 17106 23938 17118
rect 23886 17042 23938 17054
rect 24670 17106 24722 17118
rect 24670 17042 24722 17054
rect 25342 17106 25394 17118
rect 25342 17042 25394 17054
rect 16270 16994 16322 17006
rect 16270 16930 16322 16942
rect 17390 16994 17442 17006
rect 17390 16930 17442 16942
rect 17950 16994 18002 17006
rect 18498 16942 18510 16994
rect 18562 16942 18574 16994
rect 24210 16942 24222 16994
rect 24274 16942 24286 16994
rect 26450 16942 26462 16994
rect 26514 16942 26526 16994
rect 17950 16930 18002 16942
rect 16158 16882 16210 16894
rect 4274 16830 4286 16882
rect 4338 16830 4350 16882
rect 15698 16830 15710 16882
rect 15762 16830 15774 16882
rect 16158 16818 16210 16830
rect 17726 16882 17778 16894
rect 22306 16830 22318 16882
rect 22370 16830 22382 16882
rect 25666 16830 25678 16882
rect 25730 16830 25742 16882
rect 17726 16818 17778 16830
rect 1934 16770 1986 16782
rect 17838 16770 17890 16782
rect 12786 16718 12798 16770
rect 12850 16718 12862 16770
rect 14914 16718 14926 16770
rect 14978 16718 14990 16770
rect 28578 16718 28590 16770
rect 28642 16718 28654 16770
rect 1934 16706 1986 16718
rect 17838 16706 17890 16718
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 13694 16322 13746 16334
rect 13694 16258 13746 16270
rect 19070 16322 19122 16334
rect 25454 16322 25506 16334
rect 23090 16270 23102 16322
rect 23154 16319 23166 16322
rect 23314 16319 23326 16322
rect 23154 16273 23326 16319
rect 23154 16270 23166 16273
rect 23314 16270 23326 16273
rect 23378 16270 23390 16322
rect 25778 16270 25790 16322
rect 25842 16270 25854 16322
rect 19070 16258 19122 16270
rect 25454 16258 25506 16270
rect 1934 16210 1986 16222
rect 1934 16146 1986 16158
rect 19294 16210 19346 16222
rect 19294 16146 19346 16158
rect 25230 16210 25282 16222
rect 25230 16146 25282 16158
rect 14030 16098 14082 16110
rect 4274 16046 4286 16098
rect 4338 16046 4350 16098
rect 14030 16034 14082 16046
rect 14478 16098 14530 16110
rect 14478 16034 14530 16046
rect 14702 16098 14754 16110
rect 14702 16034 14754 16046
rect 14926 16098 14978 16110
rect 14926 16034 14978 16046
rect 17166 16098 17218 16110
rect 17166 16034 17218 16046
rect 18958 16098 19010 16110
rect 18958 16034 19010 16046
rect 19518 16098 19570 16110
rect 19518 16034 19570 16046
rect 20526 16098 20578 16110
rect 20526 16034 20578 16046
rect 21198 16098 21250 16110
rect 21198 16034 21250 16046
rect 21870 16098 21922 16110
rect 23326 16098 23378 16110
rect 22642 16046 22654 16098
rect 22706 16046 22718 16098
rect 21870 16034 21922 16046
rect 23326 16034 23378 16046
rect 23886 16098 23938 16110
rect 23886 16034 23938 16046
rect 24222 16098 24274 16110
rect 24222 16034 24274 16046
rect 13694 15986 13746 15998
rect 13694 15922 13746 15934
rect 13806 15986 13858 15998
rect 13806 15922 13858 15934
rect 15150 15986 15202 15998
rect 15150 15922 15202 15934
rect 15262 15986 15314 15998
rect 18622 15986 18674 15998
rect 16818 15934 16830 15986
rect 16882 15934 16894 15986
rect 15262 15922 15314 15934
rect 18622 15922 18674 15934
rect 21646 15986 21698 15998
rect 23998 15986 24050 15998
rect 22866 15934 22878 15986
rect 22930 15934 22942 15986
rect 21646 15922 21698 15934
rect 23998 15922 24050 15934
rect 14590 15874 14642 15886
rect 20638 15874 20690 15886
rect 18946 15822 18958 15874
rect 19010 15822 19022 15874
rect 14590 15810 14642 15822
rect 20638 15810 20690 15822
rect 20862 15874 20914 15886
rect 20862 15810 20914 15822
rect 21534 15874 21586 15886
rect 21534 15810 21586 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 14590 15538 14642 15550
rect 14590 15474 14642 15486
rect 21422 15538 21474 15550
rect 21422 15474 21474 15486
rect 22542 15538 22594 15550
rect 22542 15474 22594 15486
rect 25678 15538 25730 15550
rect 25678 15474 25730 15486
rect 18174 15426 18226 15438
rect 13346 15374 13358 15426
rect 13410 15374 13422 15426
rect 18174 15362 18226 15374
rect 21982 15426 22034 15438
rect 21982 15362 22034 15374
rect 25230 15426 25282 15438
rect 25230 15362 25282 15374
rect 26126 15426 26178 15438
rect 26126 15362 26178 15374
rect 21198 15314 21250 15326
rect 22206 15314 22258 15326
rect 14130 15262 14142 15314
rect 14194 15262 14206 15314
rect 20962 15262 20974 15314
rect 21026 15262 21038 15314
rect 21634 15262 21646 15314
rect 21698 15262 21710 15314
rect 21198 15250 21250 15262
rect 22206 15250 22258 15262
rect 22430 15314 22482 15326
rect 22430 15250 22482 15262
rect 25566 15314 25618 15326
rect 25566 15250 25618 15262
rect 25790 15314 25842 15326
rect 26450 15262 26462 15314
rect 26514 15262 26526 15314
rect 25790 15250 25842 15262
rect 21310 15202 21362 15214
rect 11218 15150 11230 15202
rect 11282 15150 11294 15202
rect 21310 15138 21362 15150
rect 22318 15202 22370 15214
rect 22318 15138 22370 15150
rect 26238 15202 26290 15214
rect 26238 15138 26290 15150
rect 18062 15090 18114 15102
rect 18062 15026 18114 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 22654 14754 22706 14766
rect 22654 14690 22706 14702
rect 23438 14754 23490 14766
rect 23438 14690 23490 14702
rect 19518 14642 19570 14654
rect 16930 14590 16942 14642
rect 16994 14590 17006 14642
rect 19058 14590 19070 14642
rect 19122 14590 19134 14642
rect 19518 14578 19570 14590
rect 24334 14642 24386 14654
rect 25442 14590 25454 14642
rect 25506 14590 25518 14642
rect 27570 14590 27582 14642
rect 27634 14590 27646 14642
rect 24334 14578 24386 14590
rect 15598 14530 15650 14542
rect 23214 14530 23266 14542
rect 16146 14478 16158 14530
rect 16210 14478 16222 14530
rect 22530 14478 22542 14530
rect 22594 14478 22606 14530
rect 22754 14478 22766 14530
rect 22818 14478 22830 14530
rect 23538 14478 23550 14530
rect 23602 14478 23614 14530
rect 24658 14478 24670 14530
rect 24722 14478 24734 14530
rect 15598 14466 15650 14478
rect 23214 14466 23266 14478
rect 15710 14306 15762 14318
rect 15710 14242 15762 14254
rect 15934 14306 15986 14318
rect 15934 14242 15986 14254
rect 22990 14306 23042 14318
rect 22990 14242 23042 14254
rect 23774 14306 23826 14318
rect 23774 14242 23826 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 20974 13970 21026 13982
rect 20974 13906 21026 13918
rect 21422 13970 21474 13982
rect 21422 13906 21474 13918
rect 17390 13858 17442 13870
rect 17390 13794 17442 13806
rect 19406 13858 19458 13870
rect 19406 13794 19458 13806
rect 19518 13858 19570 13870
rect 19518 13794 19570 13806
rect 19742 13858 19794 13870
rect 19742 13794 19794 13806
rect 20302 13858 20354 13870
rect 22530 13806 22542 13858
rect 22594 13806 22606 13858
rect 25218 13806 25230 13858
rect 25282 13806 25294 13858
rect 20302 13794 20354 13806
rect 17614 13746 17666 13758
rect 13570 13694 13582 13746
rect 13634 13694 13646 13746
rect 17614 13682 17666 13694
rect 17950 13746 18002 13758
rect 17950 13682 18002 13694
rect 18174 13746 18226 13758
rect 18174 13682 18226 13694
rect 19854 13746 19906 13758
rect 19854 13682 19906 13694
rect 20414 13746 20466 13758
rect 25566 13746 25618 13758
rect 21858 13694 21870 13746
rect 21922 13694 21934 13746
rect 20414 13682 20466 13694
rect 25566 13682 25618 13694
rect 20078 13634 20130 13646
rect 14354 13582 14366 13634
rect 14418 13582 14430 13634
rect 16482 13582 16494 13634
rect 16546 13582 16558 13634
rect 24658 13582 24670 13634
rect 24722 13582 24734 13634
rect 20078 13570 20130 13582
rect 17502 13522 17554 13534
rect 17502 13458 17554 13470
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 16718 13074 16770 13086
rect 20626 13022 20638 13074
rect 20690 13022 20702 13074
rect 22082 13022 22094 13074
rect 22146 13022 22158 13074
rect 24210 13022 24222 13074
rect 24274 13022 24286 13074
rect 16718 13010 16770 13022
rect 17714 12910 17726 12962
rect 17778 12910 17790 12962
rect 21410 12910 21422 12962
rect 21474 12910 21486 12962
rect 18498 12798 18510 12850
rect 18562 12798 18574 12850
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 21086 12402 21138 12414
rect 21086 12338 21138 12350
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 26126 5234 26178 5246
rect 26126 5170 26178 5182
rect 25330 5070 25342 5122
rect 25394 5070 25406 5122
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 19058 4286 19070 4338
rect 19122 4286 19134 4338
rect 25218 4286 25230 4338
rect 25282 4286 25294 4338
rect 20078 4114 20130 4126
rect 20078 4050 20130 4062
rect 26238 4114 26290 4126
rect 26238 4050 26290 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 29374 3666 29426 3678
rect 29374 3602 29426 3614
rect 16930 3502 16942 3554
rect 16994 3502 17006 3554
rect 20738 3502 20750 3554
rect 20802 3502 20814 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 18498 3390 18510 3442
rect 18562 3390 18574 3442
rect 21758 3330 21810 3342
rect 21758 3266 21810 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 18846 38558 18898 38610
rect 19966 38558 20018 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 18062 38222 18114 38274
rect 22430 38222 22482 38274
rect 26126 38222 26178 38274
rect 29374 38222 29426 38274
rect 17054 37998 17106 38050
rect 21422 37998 21474 38050
rect 25230 37998 25282 38050
rect 28590 37998 28642 38050
rect 19966 37886 20018 37938
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 18398 37438 18450 37490
rect 21422 37438 21474 37490
rect 17390 37214 17442 37266
rect 20414 37214 20466 37266
rect 28254 37214 28306 37266
rect 26014 37102 26066 37154
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 1710 36318 1762 36370
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 15710 28590 15762 28642
rect 15822 28590 15874 28642
rect 16158 28590 16210 28642
rect 16382 28590 16434 28642
rect 17278 28590 17330 28642
rect 16718 28478 16770 28530
rect 19518 28478 19570 28530
rect 19630 28478 19682 28530
rect 20526 28478 20578 28530
rect 20638 28478 20690 28530
rect 15934 28366 15986 28418
rect 16606 28366 16658 28418
rect 19294 28366 19346 28418
rect 20862 28366 20914 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 14590 27918 14642 27970
rect 18846 27918 18898 27970
rect 18958 27918 19010 27970
rect 13806 27806 13858 27858
rect 18622 27806 18674 27858
rect 22206 27806 22258 27858
rect 16718 27694 16770 27746
rect 17614 27694 17666 27746
rect 19294 27694 19346 27746
rect 21422 27694 21474 27746
rect 22766 27694 22818 27746
rect 25454 27694 25506 27746
rect 25902 27694 25954 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 21422 27246 21474 27298
rect 16382 27134 16434 27186
rect 18174 27134 18226 27186
rect 20302 27134 20354 27186
rect 25006 27134 25058 27186
rect 28254 27134 28306 27186
rect 13582 27022 13634 27074
rect 16606 27022 16658 27074
rect 16942 27022 16994 27074
rect 17502 27022 17554 27074
rect 21310 27022 21362 27074
rect 22206 27022 22258 27074
rect 25454 27022 25506 27074
rect 14254 26910 14306 26962
rect 16830 26910 16882 26962
rect 20750 26910 20802 26962
rect 22878 26910 22930 26962
rect 26126 26910 26178 26962
rect 21422 26798 21474 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 14814 26462 14866 26514
rect 16606 26462 16658 26514
rect 17614 26462 17666 26514
rect 21870 26462 21922 26514
rect 23102 26462 23154 26514
rect 26462 26462 26514 26514
rect 14926 26350 14978 26402
rect 24222 26350 24274 26402
rect 25566 26350 25618 26402
rect 17950 26238 18002 26290
rect 18622 26238 18674 26290
rect 22990 26238 23042 26290
rect 23214 26238 23266 26290
rect 23550 26238 23602 26290
rect 23886 26238 23938 26290
rect 23998 26238 24050 26290
rect 24446 26238 24498 26290
rect 25118 26238 25170 26290
rect 25678 26238 25730 26290
rect 26238 26238 26290 26290
rect 19294 26126 19346 26178
rect 21422 26126 21474 26178
rect 25342 26126 25394 26178
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 24894 25678 24946 25730
rect 24782 25566 24834 25618
rect 24558 25454 24610 25506
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 19406 24894 19458 24946
rect 19742 24894 19794 24946
rect 20078 24894 20130 24946
rect 21982 24894 22034 24946
rect 20302 24782 20354 24834
rect 4286 24670 4338 24722
rect 13806 24670 13858 24722
rect 14366 24670 14418 24722
rect 17390 24670 17442 24722
rect 17614 24670 17666 24722
rect 17838 24670 17890 24722
rect 19294 24670 19346 24722
rect 19518 24670 19570 24722
rect 20414 24670 20466 24722
rect 21422 24670 21474 24722
rect 11006 24558 11058 24610
rect 13134 24558 13186 24610
rect 17502 24558 17554 24610
rect 1934 24446 1986 24498
rect 21646 24446 21698 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 12798 24110 12850 24162
rect 1934 23998 1986 24050
rect 15934 23998 15986 24050
rect 18062 23998 18114 24050
rect 18510 23998 18562 24050
rect 19854 23998 19906 24050
rect 28590 23998 28642 24050
rect 40014 23998 40066 24050
rect 4286 23886 4338 23938
rect 12910 23886 12962 23938
rect 14030 23886 14082 23938
rect 15150 23886 15202 23938
rect 20302 23886 20354 23938
rect 21310 23886 21362 23938
rect 25678 23886 25730 23938
rect 37662 23886 37714 23938
rect 12798 23774 12850 23826
rect 13470 23774 13522 23826
rect 13582 23774 13634 23826
rect 14366 23774 14418 23826
rect 14590 23774 14642 23826
rect 19518 23774 19570 23826
rect 19742 23774 19794 23826
rect 21646 23774 21698 23826
rect 22206 23774 22258 23826
rect 26462 23774 26514 23826
rect 13806 23662 13858 23714
rect 14142 23662 14194 23714
rect 18846 23662 18898 23714
rect 19182 23662 19234 23714
rect 20526 23662 20578 23714
rect 21870 23662 21922 23714
rect 25342 23662 25394 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 14590 23326 14642 23378
rect 14814 23326 14866 23378
rect 15822 23326 15874 23378
rect 26462 23326 26514 23378
rect 27022 23326 27074 23378
rect 13134 23214 13186 23266
rect 22094 23214 22146 23266
rect 25454 23214 25506 23266
rect 13806 23102 13858 23154
rect 14366 23102 14418 23154
rect 14478 23102 14530 23154
rect 14702 23102 14754 23154
rect 16158 23102 16210 23154
rect 16382 23102 16434 23154
rect 18286 23102 18338 23154
rect 20078 23102 20130 23154
rect 25342 23102 25394 23154
rect 25678 23102 25730 23154
rect 26014 23102 26066 23154
rect 26238 23102 26290 23154
rect 26686 23102 26738 23154
rect 26910 23102 26962 23154
rect 11006 22990 11058 23042
rect 17950 22990 18002 23042
rect 18846 22990 18898 23042
rect 17390 22878 17442 22930
rect 17726 22878 17778 22930
rect 18622 22878 18674 22930
rect 27022 22878 27074 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 14142 22430 14194 22482
rect 20414 22430 20466 22482
rect 21758 22430 21810 22482
rect 28254 22430 28306 22482
rect 40014 22430 40066 22482
rect 18622 22318 18674 22370
rect 20190 22318 20242 22370
rect 22094 22318 22146 22370
rect 23886 22318 23938 22370
rect 25342 22318 25394 22370
rect 37662 22318 37714 22370
rect 18062 22206 18114 22258
rect 19518 22206 19570 22258
rect 20078 22206 20130 22258
rect 21310 22206 21362 22258
rect 23102 22206 23154 22258
rect 26126 22206 26178 22258
rect 18174 22094 18226 22146
rect 18846 22094 18898 22146
rect 21534 22094 21586 22146
rect 21758 22094 21810 22146
rect 22206 22094 22258 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 19966 21758 20018 21810
rect 21646 21758 21698 21810
rect 23774 21758 23826 21810
rect 17726 21646 17778 21698
rect 18622 21646 18674 21698
rect 19518 21646 19570 21698
rect 20974 21646 21026 21698
rect 21758 21646 21810 21698
rect 22990 21646 23042 21698
rect 23550 21646 23602 21698
rect 24670 21646 24722 21698
rect 25678 21646 25730 21698
rect 25902 21646 25954 21698
rect 26238 21646 26290 21698
rect 17502 21534 17554 21586
rect 18398 21534 18450 21586
rect 19406 21534 19458 21586
rect 20862 21534 20914 21586
rect 22878 21534 22930 21586
rect 24334 21534 24386 21586
rect 25342 21534 25394 21586
rect 25454 21534 25506 21586
rect 26350 21534 26402 21586
rect 27694 21534 27746 21586
rect 28142 21534 28194 21586
rect 28366 21534 28418 21586
rect 37662 21534 37714 21586
rect 20526 21422 20578 21474
rect 25566 21422 25618 21474
rect 26686 21422 26738 21474
rect 19518 21310 19570 21362
rect 26574 21310 26626 21362
rect 27134 21310 27186 21362
rect 27246 21310 27298 21362
rect 27470 21310 27522 21362
rect 28030 21310 28082 21362
rect 40014 21310 40066 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 18846 20974 18898 21026
rect 19182 20974 19234 21026
rect 17054 20862 17106 20914
rect 20190 20862 20242 20914
rect 23326 20862 23378 20914
rect 25342 20862 25394 20914
rect 26462 20862 26514 20914
rect 28590 20862 28642 20914
rect 14814 20750 14866 20802
rect 15038 20750 15090 20802
rect 16494 20750 16546 20802
rect 17390 20750 17442 20802
rect 17950 20750 18002 20802
rect 18174 20750 18226 20802
rect 19294 20750 19346 20802
rect 19854 20750 19906 20802
rect 21758 20750 21810 20802
rect 22206 20750 22258 20802
rect 23102 20750 23154 20802
rect 23662 20750 23714 20802
rect 24222 20750 24274 20802
rect 24558 20750 24610 20802
rect 25678 20750 25730 20802
rect 15710 20638 15762 20690
rect 22766 20638 22818 20690
rect 24894 20638 24946 20690
rect 18510 20526 18562 20578
rect 18734 20526 18786 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 24558 20190 24610 20242
rect 24782 20190 24834 20242
rect 26014 20190 26066 20242
rect 15710 20078 15762 20130
rect 17390 20078 17442 20130
rect 24446 20078 24498 20130
rect 25230 20078 25282 20130
rect 12126 19966 12178 20018
rect 15486 19966 15538 20018
rect 18510 19966 18562 20018
rect 19742 19966 19794 20018
rect 12910 19854 12962 19906
rect 15038 19854 15090 19906
rect 16270 19854 16322 19906
rect 17950 19854 18002 19906
rect 22318 19854 22370 19906
rect 25454 19854 25506 19906
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 15262 19406 15314 19458
rect 27246 19406 27298 19458
rect 15486 19294 15538 19346
rect 18622 19294 18674 19346
rect 19294 19294 19346 19346
rect 20302 19294 20354 19346
rect 24670 19294 24722 19346
rect 17278 19182 17330 19234
rect 17950 19182 18002 19234
rect 18398 19182 18450 19234
rect 18734 19182 18786 19234
rect 19070 19182 19122 19234
rect 19406 19182 19458 19234
rect 23550 19182 23602 19234
rect 23998 19182 24050 19234
rect 26350 19182 26402 19234
rect 26574 19182 26626 19234
rect 26910 19182 26962 19234
rect 27358 19182 27410 19234
rect 27582 19182 27634 19234
rect 17054 19070 17106 19122
rect 17726 19070 17778 19122
rect 23102 19070 23154 19122
rect 24558 19070 24610 19122
rect 26126 19070 26178 19122
rect 14926 18958 14978 19010
rect 20750 18958 20802 19010
rect 26238 18958 26290 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 21086 18622 21138 18674
rect 17726 18510 17778 18562
rect 17838 18510 17890 18562
rect 18174 18510 18226 18562
rect 19518 18510 19570 18562
rect 22430 18510 22482 18562
rect 22990 18510 23042 18562
rect 26350 18510 26402 18562
rect 11678 18398 11730 18450
rect 18510 18398 18562 18450
rect 19182 18398 19234 18450
rect 19854 18398 19906 18450
rect 20302 18398 20354 18450
rect 21198 18398 21250 18450
rect 21758 18398 21810 18450
rect 23102 18398 23154 18450
rect 24110 18398 24162 18450
rect 24446 18398 24498 18450
rect 25566 18398 25618 18450
rect 37662 18398 37714 18450
rect 12350 18286 12402 18338
rect 14478 18286 14530 18338
rect 14926 18286 14978 18338
rect 20750 18286 20802 18338
rect 23326 18286 23378 18338
rect 28478 18286 28530 18338
rect 17726 18174 17778 18226
rect 18846 18174 18898 18226
rect 19182 18174 19234 18226
rect 23886 18174 23938 18226
rect 24558 18174 24610 18226
rect 24670 18174 24722 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 14478 17838 14530 17890
rect 1934 17726 1986 17778
rect 9998 17726 10050 17778
rect 18510 17726 18562 17778
rect 40014 17726 40066 17778
rect 4286 17614 4338 17666
rect 12798 17614 12850 17666
rect 13582 17614 13634 17666
rect 14254 17614 14306 17666
rect 14814 17614 14866 17666
rect 17390 17614 17442 17666
rect 17726 17614 17778 17666
rect 17950 17614 18002 17666
rect 18398 17614 18450 17666
rect 18958 17614 19010 17666
rect 19518 17614 19570 17666
rect 19742 17614 19794 17666
rect 23326 17614 23378 17666
rect 23774 17614 23826 17666
rect 37662 17614 37714 17666
rect 12126 17502 12178 17554
rect 15038 17502 15090 17554
rect 17166 17502 17218 17554
rect 17502 17502 17554 17554
rect 18622 17502 18674 17554
rect 21870 17502 21922 17554
rect 24334 17502 24386 17554
rect 25902 17502 25954 17554
rect 14142 17390 14194 17442
rect 15486 17390 15538 17442
rect 19630 17390 19682 17442
rect 25006 17390 25058 17442
rect 26238 17390 26290 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 16494 17054 16546 17106
rect 16830 17054 16882 17106
rect 23886 17054 23938 17106
rect 24670 17054 24722 17106
rect 25342 17054 25394 17106
rect 16270 16942 16322 16994
rect 17390 16942 17442 16994
rect 17950 16942 18002 16994
rect 18510 16942 18562 16994
rect 24222 16942 24274 16994
rect 26462 16942 26514 16994
rect 4286 16830 4338 16882
rect 15710 16830 15762 16882
rect 16158 16830 16210 16882
rect 17726 16830 17778 16882
rect 22318 16830 22370 16882
rect 25678 16830 25730 16882
rect 1934 16718 1986 16770
rect 12798 16718 12850 16770
rect 14926 16718 14978 16770
rect 17838 16718 17890 16770
rect 28590 16718 28642 16770
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 13694 16270 13746 16322
rect 19070 16270 19122 16322
rect 23102 16270 23154 16322
rect 23326 16270 23378 16322
rect 25454 16270 25506 16322
rect 25790 16270 25842 16322
rect 1934 16158 1986 16210
rect 19294 16158 19346 16210
rect 25230 16158 25282 16210
rect 4286 16046 4338 16098
rect 14030 16046 14082 16098
rect 14478 16046 14530 16098
rect 14702 16046 14754 16098
rect 14926 16046 14978 16098
rect 17166 16046 17218 16098
rect 18958 16046 19010 16098
rect 19518 16046 19570 16098
rect 20526 16046 20578 16098
rect 21198 16046 21250 16098
rect 21870 16046 21922 16098
rect 22654 16046 22706 16098
rect 23326 16046 23378 16098
rect 23886 16046 23938 16098
rect 24222 16046 24274 16098
rect 13694 15934 13746 15986
rect 13806 15934 13858 15986
rect 15150 15934 15202 15986
rect 15262 15934 15314 15986
rect 16830 15934 16882 15986
rect 18622 15934 18674 15986
rect 21646 15934 21698 15986
rect 22878 15934 22930 15986
rect 23998 15934 24050 15986
rect 14590 15822 14642 15874
rect 18958 15822 19010 15874
rect 20638 15822 20690 15874
rect 20862 15822 20914 15874
rect 21534 15822 21586 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 14590 15486 14642 15538
rect 21422 15486 21474 15538
rect 22542 15486 22594 15538
rect 25678 15486 25730 15538
rect 13358 15374 13410 15426
rect 18174 15374 18226 15426
rect 21982 15374 22034 15426
rect 25230 15374 25282 15426
rect 26126 15374 26178 15426
rect 14142 15262 14194 15314
rect 20974 15262 21026 15314
rect 21198 15262 21250 15314
rect 21646 15262 21698 15314
rect 22206 15262 22258 15314
rect 22430 15262 22482 15314
rect 25566 15262 25618 15314
rect 25790 15262 25842 15314
rect 26462 15262 26514 15314
rect 11230 15150 11282 15202
rect 21310 15150 21362 15202
rect 22318 15150 22370 15202
rect 26238 15150 26290 15202
rect 18062 15038 18114 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 22654 14702 22706 14754
rect 23438 14702 23490 14754
rect 16942 14590 16994 14642
rect 19070 14590 19122 14642
rect 19518 14590 19570 14642
rect 24334 14590 24386 14642
rect 25454 14590 25506 14642
rect 27582 14590 27634 14642
rect 15598 14478 15650 14530
rect 16158 14478 16210 14530
rect 22542 14478 22594 14530
rect 22766 14478 22818 14530
rect 23214 14478 23266 14530
rect 23550 14478 23602 14530
rect 24670 14478 24722 14530
rect 15710 14254 15762 14306
rect 15934 14254 15986 14306
rect 22990 14254 23042 14306
rect 23774 14254 23826 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 20974 13918 21026 13970
rect 21422 13918 21474 13970
rect 17390 13806 17442 13858
rect 19406 13806 19458 13858
rect 19518 13806 19570 13858
rect 19742 13806 19794 13858
rect 20302 13806 20354 13858
rect 22542 13806 22594 13858
rect 25230 13806 25282 13858
rect 13582 13694 13634 13746
rect 17614 13694 17666 13746
rect 17950 13694 18002 13746
rect 18174 13694 18226 13746
rect 19854 13694 19906 13746
rect 20414 13694 20466 13746
rect 21870 13694 21922 13746
rect 25566 13694 25618 13746
rect 14366 13582 14418 13634
rect 16494 13582 16546 13634
rect 20078 13582 20130 13634
rect 24670 13582 24722 13634
rect 17502 13470 17554 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 16718 13022 16770 13074
rect 20638 13022 20690 13074
rect 22094 13022 22146 13074
rect 24222 13022 24274 13074
rect 17726 12910 17778 12962
rect 21422 12910 21474 12962
rect 18510 12798 18562 12850
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 21086 12350 21138 12402
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 26126 5182 26178 5234
rect 25342 5070 25394 5122
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 19070 4286 19122 4338
rect 25230 4286 25282 4338
rect 20078 4062 20130 4114
rect 26238 4062 26290 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 25566 3614 25618 3666
rect 29374 3614 29426 3666
rect 16942 3502 16994 3554
rect 20750 3502 20802 3554
rect 24558 3502 24610 3554
rect 28590 3502 28642 3554
rect 18510 3390 18562 3442
rect 21758 3278 21810 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 16128 41200 16240 42000
rect 16800 41200 16912 42000
rect 18816 41200 18928 42000
rect 20160 41200 20272 42000
rect 22176 41200 22288 42000
rect 24864 41200 24976 42000
rect 25536 41200 25648 42000
rect 26208 41200 26320 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 16156 37492 16212 41200
rect 16828 38276 16884 41200
rect 18844 38610 18900 41200
rect 18844 38558 18846 38610
rect 18898 38558 18900 38610
rect 18844 38546 18900 38558
rect 19964 38610 20020 38622
rect 19964 38558 19966 38610
rect 20018 38558 20020 38610
rect 16828 38210 16884 38220
rect 18060 38276 18116 38286
rect 18060 38182 18116 38220
rect 16156 37426 16212 37436
rect 17052 38050 17108 38062
rect 17052 37998 17054 38050
rect 17106 37998 17108 38050
rect 15820 37268 15876 37278
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 1708 36372 1764 36382
rect 1708 36278 1764 36316
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 15708 28756 15764 28766
rect 14588 28644 14644 28654
rect 4172 28308 4228 28318
rect 1932 24500 1988 24510
rect 1932 24406 1988 24444
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 1932 23538 1988 23548
rect 4172 20020 4228 28252
rect 14588 27970 14644 28588
rect 15708 28642 15764 28700
rect 15708 28590 15710 28642
rect 15762 28590 15764 28642
rect 15708 28578 15764 28590
rect 15820 28644 15876 37212
rect 17052 31948 17108 37998
rect 19964 37938 20020 38558
rect 19964 37886 19966 37938
rect 20018 37886 20020 37938
rect 19964 37874 20020 37886
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 18396 37492 18452 37502
rect 18396 37398 18452 37436
rect 20188 37492 20244 41200
rect 22204 38276 22260 41200
rect 24892 38612 24948 41200
rect 24892 38546 24948 38556
rect 22428 38276 22484 38286
rect 22204 38274 22484 38276
rect 22204 38222 22430 38274
rect 22482 38222 22484 38274
rect 22204 38220 22484 38222
rect 22428 38210 22484 38220
rect 21420 38052 21476 38062
rect 20188 37426 20244 37436
rect 20636 38050 21476 38052
rect 20636 37998 21422 38050
rect 21474 37998 21476 38050
rect 20636 37996 21476 37998
rect 17388 37268 17444 37278
rect 17388 37174 17444 37212
rect 20412 37266 20468 37278
rect 20412 37214 20414 37266
rect 20466 37214 20468 37266
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20412 31948 20468 37214
rect 16828 31892 17108 31948
rect 20300 31892 20468 31948
rect 15820 28642 16100 28644
rect 15820 28590 15822 28642
rect 15874 28590 16100 28642
rect 15820 28588 16100 28590
rect 15820 28578 15876 28588
rect 14588 27918 14590 27970
rect 14642 27918 14644 27970
rect 14588 27906 14644 27918
rect 14924 28420 14980 28430
rect 13804 27858 13860 27870
rect 13804 27806 13806 27858
rect 13858 27806 13860 27858
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 13580 27076 13636 27086
rect 13804 27076 13860 27806
rect 13580 27074 13860 27076
rect 13580 27022 13582 27074
rect 13634 27022 13860 27074
rect 13580 27020 13860 27022
rect 13580 27010 13636 27020
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4284 24724 4340 24734
rect 4284 24630 4340 24668
rect 10780 24724 10836 24734
rect 13692 24724 13748 27020
rect 14252 26964 14308 26974
rect 14252 26962 14868 26964
rect 14252 26910 14254 26962
rect 14306 26910 14868 26962
rect 14252 26908 14868 26910
rect 14252 26898 14308 26908
rect 14812 26514 14868 26908
rect 14812 26462 14814 26514
rect 14866 26462 14868 26514
rect 14812 26450 14868 26462
rect 14924 26402 14980 28364
rect 15932 28420 15988 28430
rect 15932 28326 15988 28364
rect 16044 28308 16100 28588
rect 16156 28642 16212 28654
rect 16156 28590 16158 28642
rect 16210 28590 16212 28642
rect 16156 28532 16212 28590
rect 16380 28644 16436 28654
rect 16380 28550 16436 28588
rect 16156 28466 16212 28476
rect 16716 28530 16772 28542
rect 16716 28478 16718 28530
rect 16770 28478 16772 28530
rect 16604 28420 16660 28430
rect 16492 28418 16660 28420
rect 16492 28366 16606 28418
rect 16658 28366 16660 28418
rect 16492 28364 16660 28366
rect 16044 28252 16436 28308
rect 16380 27186 16436 28252
rect 16380 27134 16382 27186
rect 16434 27134 16436 27186
rect 16380 27122 16436 27134
rect 16492 26908 16548 28364
rect 16604 28354 16660 28364
rect 16716 27972 16772 28478
rect 16604 27916 16772 27972
rect 16604 27074 16660 27916
rect 16716 27748 16772 27758
rect 16828 27748 16884 31892
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 17276 28644 17332 28654
rect 17276 28550 17332 28588
rect 19516 28532 19572 28542
rect 19516 28438 19572 28476
rect 19628 28530 19684 28542
rect 19628 28478 19630 28530
rect 19682 28478 19684 28530
rect 16716 27746 16884 27748
rect 16716 27694 16718 27746
rect 16770 27694 16884 27746
rect 16716 27692 16884 27694
rect 16716 27682 16772 27692
rect 16604 27022 16606 27074
rect 16658 27022 16660 27074
rect 16604 27010 16660 27022
rect 14924 26350 14926 26402
rect 14978 26350 14980 26402
rect 14924 26338 14980 26350
rect 16156 26852 16548 26908
rect 16828 26962 16884 27692
rect 16940 28420 16996 28430
rect 19292 28420 19348 28430
rect 16940 27076 16996 28364
rect 18956 28418 19348 28420
rect 18956 28366 19294 28418
rect 19346 28366 19348 28418
rect 18956 28364 19348 28366
rect 18844 27970 18900 27982
rect 18844 27918 18846 27970
rect 18898 27918 18900 27970
rect 18620 27860 18676 27870
rect 18172 27858 18676 27860
rect 18172 27806 18622 27858
rect 18674 27806 18676 27858
rect 18172 27804 18676 27806
rect 17612 27748 17668 27758
rect 16940 26982 16996 27020
rect 17500 27746 17668 27748
rect 17500 27694 17614 27746
rect 17666 27694 17668 27746
rect 17500 27692 17668 27694
rect 17500 27074 17556 27692
rect 17612 27682 17668 27692
rect 18172 27186 18228 27804
rect 18620 27794 18676 27804
rect 18172 27134 18174 27186
rect 18226 27134 18228 27186
rect 18172 27122 18228 27134
rect 17500 27022 17502 27074
rect 17554 27022 17556 27074
rect 16828 26910 16830 26962
rect 16882 26910 16884 26962
rect 16828 26898 16884 26910
rect 16604 26852 16660 26862
rect 15148 25284 15204 25294
rect 13804 24724 13860 24734
rect 14364 24724 14420 24734
rect 10836 24668 10948 24724
rect 10780 24658 10836 24668
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4284 23940 4340 23950
rect 4284 23846 4340 23884
rect 10892 23828 10948 24668
rect 13692 24722 14420 24724
rect 13692 24670 13806 24722
rect 13858 24670 14366 24722
rect 14418 24670 14420 24722
rect 13692 24668 14420 24670
rect 11004 24610 11060 24622
rect 11004 24558 11006 24610
rect 11058 24558 11060 24610
rect 11004 23940 11060 24558
rect 13132 24612 13188 24622
rect 13132 24610 13300 24612
rect 13132 24558 13134 24610
rect 13186 24558 13300 24610
rect 13132 24556 13300 24558
rect 13132 24546 13188 24556
rect 12796 24162 12852 24174
rect 12796 24110 12798 24162
rect 12850 24110 12852 24162
rect 12796 24052 12852 24110
rect 12796 23986 12852 23996
rect 11004 23874 11060 23884
rect 12908 23940 12964 23950
rect 12908 23938 13076 23940
rect 12908 23886 12910 23938
rect 12962 23886 13076 23938
rect 12908 23884 13076 23886
rect 12908 23874 12964 23884
rect 10892 23044 10948 23772
rect 12796 23828 12852 23838
rect 12796 23734 12852 23772
rect 13020 23828 13076 23884
rect 13020 23762 13076 23772
rect 13132 23716 13188 23726
rect 13132 23266 13188 23660
rect 13244 23380 13300 24556
rect 13580 23940 13636 23950
rect 13468 23828 13524 23838
rect 13468 23734 13524 23772
rect 13580 23826 13636 23884
rect 13580 23774 13582 23826
rect 13634 23774 13636 23826
rect 13580 23762 13636 23774
rect 13244 23314 13300 23324
rect 13692 23604 13748 24668
rect 13804 24658 13860 24668
rect 14364 24658 14420 24668
rect 14028 24052 14084 24062
rect 14028 23938 14084 23996
rect 14028 23886 14030 23938
rect 14082 23886 14084 23938
rect 14028 23874 14084 23886
rect 15148 23938 15204 25228
rect 15932 24612 15988 24622
rect 15932 24050 15988 24556
rect 15932 23998 15934 24050
rect 15986 23998 15988 24050
rect 15932 23986 15988 23998
rect 16156 24052 16212 26852
rect 16604 26514 16660 26796
rect 17500 26852 17556 27022
rect 17500 26786 17556 26796
rect 17612 27076 17668 27086
rect 16604 26462 16606 26514
rect 16658 26462 16660 26514
rect 16604 26450 16660 26462
rect 17612 26514 17668 27020
rect 17612 26462 17614 26514
rect 17666 26462 17668 26514
rect 17612 26450 17668 26462
rect 18620 26852 18676 26862
rect 17948 26292 18004 26302
rect 17948 26290 18452 26292
rect 17948 26238 17950 26290
rect 18002 26238 18452 26290
rect 17948 26236 18452 26238
rect 17948 26226 18004 26236
rect 15148 23886 15150 23938
rect 15202 23886 15204 23938
rect 14364 23826 14420 23838
rect 14364 23774 14366 23826
rect 14418 23774 14420 23826
rect 13804 23716 13860 23726
rect 14140 23716 14196 23726
rect 13804 23714 14084 23716
rect 13804 23662 13806 23714
rect 13858 23662 14084 23714
rect 13804 23660 14084 23662
rect 13804 23650 13860 23660
rect 13132 23214 13134 23266
rect 13186 23214 13188 23266
rect 13132 23202 13188 23214
rect 13692 23156 13748 23548
rect 14028 23268 14084 23660
rect 14140 23622 14196 23660
rect 14364 23716 14420 23774
rect 14588 23828 14644 23838
rect 14588 23826 14868 23828
rect 14588 23774 14590 23826
rect 14642 23774 14868 23826
rect 14588 23772 14868 23774
rect 14588 23762 14644 23772
rect 14420 23660 14532 23716
rect 14364 23650 14420 23660
rect 14476 23380 14532 23660
rect 14364 23324 14532 23380
rect 14588 23380 14644 23390
rect 14028 23212 14308 23268
rect 13804 23156 13860 23166
rect 13692 23154 14196 23156
rect 13692 23102 13806 23154
rect 13858 23102 14196 23154
rect 13692 23100 14196 23102
rect 13804 23090 13860 23100
rect 11004 23044 11060 23054
rect 10892 23042 11060 23044
rect 10892 22990 11006 23042
rect 11058 22990 11060 23042
rect 10892 22988 11060 22990
rect 11004 22978 11060 22988
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 14140 22482 14196 23100
rect 14252 22932 14308 23212
rect 14364 23154 14420 23324
rect 14588 23286 14644 23324
rect 14812 23380 14868 23772
rect 15148 23604 15204 23886
rect 15148 23538 15204 23548
rect 14812 23286 14868 23324
rect 15820 23380 15876 23390
rect 15820 23286 15876 23324
rect 14364 23102 14366 23154
rect 14418 23102 14420 23154
rect 14364 23090 14420 23102
rect 14476 23154 14532 23166
rect 14476 23102 14478 23154
rect 14530 23102 14532 23154
rect 14476 22932 14532 23102
rect 14252 22876 14532 22932
rect 14700 23154 14756 23166
rect 14700 23102 14702 23154
rect 14754 23102 14756 23154
rect 14140 22430 14142 22482
rect 14194 22430 14196 22482
rect 14140 22418 14196 22430
rect 14700 22484 14756 23102
rect 16156 23154 16212 23996
rect 17388 24722 17444 24734
rect 17388 24670 17390 24722
rect 17442 24670 17444 24722
rect 17052 23716 17108 23726
rect 17108 23660 17220 23716
rect 17052 23650 17108 23660
rect 16156 23102 16158 23154
rect 16210 23102 16212 23154
rect 16156 23090 16212 23102
rect 16380 23156 16436 23166
rect 16380 23062 16436 23100
rect 14700 22418 14756 22428
rect 17052 22820 17108 22830
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 17052 20914 17108 22764
rect 17052 20862 17054 20914
rect 17106 20862 17108 20914
rect 17052 20850 17108 20862
rect 14476 20804 14532 20814
rect 12124 20020 12180 20030
rect 4172 19954 4228 19964
rect 11788 20018 12180 20020
rect 11788 19966 12126 20018
rect 12178 19966 12180 20018
rect 11788 19964 12180 19966
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 11676 18452 11732 18462
rect 11788 18452 11844 19964
rect 12124 19954 12180 19964
rect 12908 19908 12964 19918
rect 12908 19814 12964 19852
rect 11676 18450 11788 18452
rect 11676 18398 11678 18450
rect 11730 18398 11788 18450
rect 11676 18396 11788 18398
rect 11676 18386 11732 18396
rect 11788 18358 11844 18396
rect 12796 18452 12852 18462
rect 12348 18340 12404 18350
rect 12348 18246 12404 18284
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1932 17780 1988 17790
rect 1932 17686 1988 17724
rect 9996 17778 10052 17790
rect 9996 17726 9998 17778
rect 10050 17726 10052 17778
rect 4284 17668 4340 17678
rect 4284 17574 4340 17612
rect 9996 17668 10052 17726
rect 1932 16884 1988 16894
rect 1932 16770 1988 16828
rect 4284 16884 4340 16894
rect 4284 16790 4340 16828
rect 1932 16718 1934 16770
rect 1986 16718 1988 16770
rect 1932 16706 1988 16718
rect 9996 16772 10052 17612
rect 12796 17668 12852 18396
rect 14476 18338 14532 20748
rect 14812 20802 14868 20814
rect 14812 20750 14814 20802
rect 14866 20750 14868 20802
rect 14812 20188 14868 20750
rect 15036 20804 15092 20814
rect 15036 20710 15092 20748
rect 16492 20804 16548 20814
rect 16492 20710 16548 20748
rect 15708 20692 15764 20702
rect 15484 20690 15764 20692
rect 15484 20638 15710 20690
rect 15762 20638 15764 20690
rect 15484 20636 15764 20638
rect 14812 20132 15092 20188
rect 15036 19906 15092 20076
rect 15484 20018 15540 20636
rect 15708 20626 15764 20636
rect 15484 19966 15486 20018
rect 15538 19966 15540 20018
rect 15484 19954 15540 19966
rect 15708 20130 15764 20142
rect 15708 20078 15710 20130
rect 15762 20078 15764 20130
rect 15036 19854 15038 19906
rect 15090 19854 15092 19906
rect 15036 19842 15092 19854
rect 15260 19908 15316 19918
rect 15260 19458 15316 19852
rect 15708 19908 15764 20078
rect 15708 19842 15764 19852
rect 16268 19908 16324 19918
rect 16268 19906 16772 19908
rect 16268 19854 16270 19906
rect 16322 19854 16772 19906
rect 16268 19852 16772 19854
rect 16268 19842 16324 19852
rect 15260 19406 15262 19458
rect 15314 19406 15316 19458
rect 15260 19394 15316 19406
rect 15484 19460 15540 19470
rect 15484 19346 15540 19404
rect 15484 19294 15486 19346
rect 15538 19294 15540 19346
rect 15484 19282 15540 19294
rect 14924 19012 14980 19022
rect 14476 18286 14478 18338
rect 14530 18286 14532 18338
rect 14476 18274 14532 18286
rect 14588 19010 14980 19012
rect 14588 18958 14926 19010
rect 14978 18958 14980 19010
rect 14588 18956 14980 18958
rect 14476 17892 14532 17902
rect 14588 17892 14644 18956
rect 14924 18946 14980 18956
rect 14476 17890 14644 17892
rect 14476 17838 14478 17890
rect 14530 17838 14644 17890
rect 14476 17836 14644 17838
rect 14812 18788 14868 18798
rect 12796 17574 12852 17612
rect 13580 17668 13636 17678
rect 13580 17574 13636 17612
rect 14252 17666 14308 17678
rect 14252 17614 14254 17666
rect 14306 17614 14308 17666
rect 12124 17554 12180 17566
rect 12124 17502 12126 17554
rect 12178 17502 12180 17554
rect 12124 17444 12180 17502
rect 14252 17556 14308 17614
rect 14252 17490 14308 17500
rect 14364 17668 14420 17678
rect 12124 17378 12180 17388
rect 14140 17444 14196 17454
rect 14140 17350 14196 17388
rect 9996 16706 10052 16716
rect 12796 16884 12852 16894
rect 12796 16770 12852 16828
rect 12796 16718 12798 16770
rect 12850 16718 12852 16770
rect 12796 16706 12852 16718
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 13692 16324 13748 16334
rect 13692 16322 14084 16324
rect 13692 16270 13694 16322
rect 13746 16270 14084 16322
rect 13692 16268 14084 16270
rect 13692 16258 13748 16268
rect 1932 16210 1988 16222
rect 1932 16158 1934 16210
rect 1986 16158 1988 16210
rect 1932 15540 1988 16158
rect 4284 16100 4340 16110
rect 4284 16006 4340 16044
rect 11228 16100 11284 16110
rect 1932 15474 1988 15484
rect 11228 15202 11284 16044
rect 13692 16100 13748 16110
rect 13692 15986 13748 16044
rect 14028 16098 14084 16268
rect 14028 16046 14030 16098
rect 14082 16046 14084 16098
rect 14028 16034 14084 16046
rect 13692 15934 13694 15986
rect 13746 15934 13748 15986
rect 13692 15922 13748 15934
rect 13804 15988 13860 15998
rect 13804 15894 13860 15932
rect 13356 15876 13412 15886
rect 13356 15426 13412 15820
rect 14364 15652 14420 17612
rect 14476 16098 14532 17836
rect 14812 17666 14868 18732
rect 14812 17614 14814 17666
rect 14866 17614 14868 17666
rect 14812 17602 14868 17614
rect 14924 18340 14980 18350
rect 14924 17668 14980 18284
rect 14924 17602 14980 17612
rect 16716 18340 16772 19852
rect 17052 19124 17108 19134
rect 17164 19124 17220 23660
rect 17388 22932 17444 24670
rect 17612 24722 17668 24734
rect 17612 24670 17614 24722
rect 17666 24670 17668 24722
rect 17500 24612 17556 24622
rect 17500 24518 17556 24556
rect 17612 23716 17668 24670
rect 17612 23650 17668 23660
rect 17836 24722 17892 24734
rect 17836 24670 17838 24722
rect 17890 24670 17892 24722
rect 17836 23156 17892 24670
rect 17836 23090 17892 23100
rect 18060 24050 18116 24062
rect 18060 23998 18062 24050
rect 18114 23998 18116 24050
rect 17948 23042 18004 23054
rect 17948 22990 17950 23042
rect 18002 22990 18004 23042
rect 17388 22838 17444 22876
rect 17724 22930 17780 22942
rect 17724 22878 17726 22930
rect 17778 22878 17780 22930
rect 17724 21698 17780 22878
rect 17948 22820 18004 22990
rect 17948 22754 18004 22764
rect 18060 22258 18116 23998
rect 18396 23604 18452 26236
rect 18620 26290 18676 26796
rect 18620 26238 18622 26290
rect 18674 26238 18676 26290
rect 18508 24052 18564 24062
rect 18620 24052 18676 26238
rect 18844 24948 18900 27918
rect 18956 27970 19012 28364
rect 19292 28354 19348 28364
rect 19628 28420 19684 28478
rect 19628 28354 19684 28364
rect 20300 28532 20356 31892
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 18956 27918 18958 27970
rect 19010 27918 19012 27970
rect 18956 27906 19012 27918
rect 19292 27748 19348 27758
rect 19292 27654 19348 27692
rect 20300 27186 20356 28476
rect 20524 28532 20580 28542
rect 20524 28438 20580 28476
rect 20636 28530 20692 37996
rect 21420 37986 21476 37996
rect 25228 38050 25284 38062
rect 25228 37998 25230 38050
rect 25282 37998 25284 38050
rect 21420 37492 21476 37502
rect 21420 37398 21476 37436
rect 22204 28644 22260 28654
rect 22260 28588 22372 28644
rect 22204 28578 22260 28588
rect 20636 28478 20638 28530
rect 20690 28478 20692 28530
rect 20636 27748 20692 28478
rect 20860 28420 20916 28430
rect 20860 28418 21364 28420
rect 20860 28366 20862 28418
rect 20914 28366 21364 28418
rect 20860 28364 21364 28366
rect 20860 28354 20916 28364
rect 20636 27682 20692 27692
rect 20300 27134 20302 27186
rect 20354 27134 20356 27186
rect 20300 27122 20356 27134
rect 21308 27074 21364 28364
rect 22204 27858 22260 27870
rect 22204 27806 22206 27858
rect 22258 27806 22260 27858
rect 21420 27746 21476 27758
rect 21420 27694 21422 27746
rect 21474 27694 21476 27746
rect 21420 27298 21476 27694
rect 21420 27246 21422 27298
rect 21474 27246 21476 27298
rect 21420 27234 21476 27246
rect 22204 27748 22260 27806
rect 22204 27076 22260 27692
rect 21308 27022 21310 27074
rect 21362 27022 21364 27074
rect 21308 27010 21364 27022
rect 21868 27074 22260 27076
rect 21868 27022 22206 27074
rect 22258 27022 22260 27074
rect 21868 27020 22260 27022
rect 20748 26964 20804 26974
rect 20748 26870 20804 26908
rect 21868 26964 21924 27020
rect 22204 27010 22260 27020
rect 21420 26852 21476 26862
rect 21196 26850 21476 26852
rect 21196 26798 21422 26850
rect 21474 26798 21476 26850
rect 21196 26796 21476 26798
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19292 26180 19348 26190
rect 19292 26178 19460 26180
rect 19292 26126 19294 26178
rect 19346 26126 19460 26178
rect 19292 26124 19460 26126
rect 19292 26114 19348 26124
rect 18844 24882 18900 24892
rect 19404 24946 19460 26124
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19404 24894 19406 24946
rect 19458 24894 19460 24946
rect 19404 24882 19460 24894
rect 19740 24948 19796 24958
rect 20076 24948 20132 24958
rect 19796 24946 20132 24948
rect 19796 24894 20078 24946
rect 20130 24894 20132 24946
rect 19796 24892 20132 24894
rect 19740 24854 19796 24892
rect 20076 24882 20132 24892
rect 20300 24834 20356 24846
rect 20300 24782 20302 24834
rect 20354 24782 20356 24834
rect 18508 24050 18676 24052
rect 18508 23998 18510 24050
rect 18562 23998 18676 24050
rect 18508 23996 18676 23998
rect 19292 24724 19348 24734
rect 18508 23986 18564 23996
rect 19292 23940 19348 24668
rect 19516 24722 19572 24734
rect 19516 24670 19518 24722
rect 19570 24670 19572 24722
rect 19516 24164 19572 24670
rect 20300 24724 20356 24782
rect 20300 24658 20356 24668
rect 20412 24722 20468 24734
rect 20412 24670 20414 24722
rect 20466 24670 20468 24722
rect 19852 24276 19908 24286
rect 19516 24098 19572 24108
rect 19740 24220 19852 24276
rect 19068 23884 19348 23940
rect 18844 23716 18900 23726
rect 18900 23660 19012 23716
rect 18844 23622 18900 23660
rect 18396 23548 18564 23604
rect 18284 23156 18340 23166
rect 18284 23062 18340 23100
rect 18060 22206 18062 22258
rect 18114 22206 18116 22258
rect 18060 22036 18116 22206
rect 18060 21970 18116 21980
rect 18172 22146 18228 22158
rect 18172 22094 18174 22146
rect 18226 22094 18228 22146
rect 17724 21646 17726 21698
rect 17778 21646 17780 21698
rect 17500 21586 17556 21598
rect 17500 21534 17502 21586
rect 17554 21534 17556 21586
rect 17388 20804 17444 20814
rect 17388 20710 17444 20748
rect 17388 20132 17444 20142
rect 17500 20132 17556 21534
rect 17724 20804 17780 21646
rect 18172 21588 18228 22094
rect 18396 21588 18452 21598
rect 18172 21586 18452 21588
rect 18172 21534 18398 21586
rect 18450 21534 18452 21586
rect 18172 21532 18452 21534
rect 18060 21364 18116 21374
rect 17724 20738 17780 20748
rect 17948 20802 18004 20814
rect 17948 20750 17950 20802
rect 18002 20750 18004 20802
rect 17724 20580 17780 20590
rect 17444 20076 17556 20132
rect 17612 20132 17668 20142
rect 17388 20038 17444 20076
rect 17612 19796 17668 20076
rect 17500 19740 17668 19796
rect 17052 19122 17220 19124
rect 17052 19070 17054 19122
rect 17106 19070 17220 19122
rect 17052 19068 17220 19070
rect 17276 19234 17332 19246
rect 17276 19182 17278 19234
rect 17330 19182 17332 19234
rect 17052 18788 17108 19068
rect 17052 18722 17108 18732
rect 15036 17554 15092 17566
rect 15036 17502 15038 17554
rect 15090 17502 15092 17554
rect 14700 17444 14756 17454
rect 14700 16884 14756 17388
rect 14700 16828 14980 16884
rect 14924 16770 14980 16828
rect 14924 16718 14926 16770
rect 14978 16718 14980 16770
rect 14924 16706 14980 16718
rect 14476 16046 14478 16098
rect 14530 16046 14532 16098
rect 14476 16034 14532 16046
rect 14700 16660 14756 16670
rect 14700 16098 14756 16604
rect 14700 16046 14702 16098
rect 14754 16046 14756 16098
rect 14700 16034 14756 16046
rect 14924 16100 14980 16110
rect 15036 16100 15092 17502
rect 15484 17556 15540 17566
rect 15484 17442 15540 17500
rect 15484 17390 15486 17442
rect 15538 17390 15540 17442
rect 15484 17332 15540 17390
rect 15484 17266 15540 17276
rect 16492 17556 16548 17566
rect 15708 17108 15764 17118
rect 15708 16882 15764 17052
rect 16492 17106 16548 17500
rect 16492 17054 16494 17106
rect 16546 17054 16548 17106
rect 16492 17042 16548 17054
rect 16716 17108 16772 18284
rect 17276 18116 17332 19182
rect 17500 18564 17556 19740
rect 17612 19572 17668 19582
rect 17612 18788 17668 19516
rect 17724 19124 17780 20524
rect 17948 20132 18004 20750
rect 17948 20066 18004 20076
rect 17948 19906 18004 19918
rect 17948 19854 17950 19906
rect 18002 19854 18004 19906
rect 17948 19572 18004 19854
rect 17948 19506 18004 19516
rect 17724 19030 17780 19068
rect 17948 19234 18004 19246
rect 17948 19182 17950 19234
rect 18002 19182 18004 19234
rect 17948 19012 18004 19182
rect 18060 19124 18116 21308
rect 18396 21140 18452 21532
rect 18396 21074 18452 21084
rect 18172 20802 18228 20814
rect 18172 20750 18174 20802
rect 18226 20750 18228 20802
rect 18172 19908 18228 20750
rect 18508 20804 18564 23548
rect 18844 23044 18900 23054
rect 18732 23042 18900 23044
rect 18732 22990 18846 23042
rect 18898 22990 18900 23042
rect 18732 22988 18900 22990
rect 18620 22930 18676 22942
rect 18620 22878 18622 22930
rect 18674 22878 18676 22930
rect 18620 22596 18676 22878
rect 18620 22530 18676 22540
rect 18620 22370 18676 22382
rect 18620 22318 18622 22370
rect 18674 22318 18676 22370
rect 18620 22036 18676 22318
rect 18620 21970 18676 21980
rect 18620 21700 18676 21710
rect 18732 21700 18788 22988
rect 18844 22978 18900 22988
rect 18844 22148 18900 22158
rect 18844 22054 18900 22092
rect 18620 21698 18788 21700
rect 18620 21646 18622 21698
rect 18674 21646 18788 21698
rect 18620 21644 18788 21646
rect 18620 21634 18676 21644
rect 18508 20748 18676 20804
rect 18508 20580 18564 20590
rect 18508 20486 18564 20524
rect 18620 20356 18676 20748
rect 18620 20290 18676 20300
rect 18732 20578 18788 21644
rect 18844 21588 18900 21598
rect 18844 21026 18900 21532
rect 18844 20974 18846 21026
rect 18898 20974 18900 21026
rect 18844 20962 18900 20974
rect 18956 20804 19012 23660
rect 19068 22932 19124 23884
rect 19516 23826 19572 23838
rect 19740 23828 19796 24220
rect 19852 24210 19908 24220
rect 19852 24050 19908 24062
rect 19852 23998 19854 24050
rect 19906 23998 19908 24050
rect 19852 23940 19908 23998
rect 19852 23874 19908 23884
rect 20300 23938 20356 23950
rect 20300 23886 20302 23938
rect 20354 23886 20356 23938
rect 19516 23774 19518 23826
rect 19570 23774 19572 23826
rect 19180 23716 19236 23726
rect 19516 23716 19572 23774
rect 19180 23714 19516 23716
rect 19180 23662 19182 23714
rect 19234 23662 19516 23714
rect 19180 23660 19516 23662
rect 19180 23650 19236 23660
rect 19516 23650 19572 23660
rect 19628 23826 19796 23828
rect 19628 23774 19742 23826
rect 19794 23774 19796 23826
rect 19628 23772 19796 23774
rect 19068 22866 19124 22876
rect 19628 22484 19684 23772
rect 19740 23762 19796 23772
rect 20300 23828 20356 23886
rect 20412 23940 20468 24670
rect 20412 23874 20468 23884
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20076 23156 20132 23166
rect 20076 23062 20132 23100
rect 19404 22428 19684 22484
rect 20076 22932 20132 22942
rect 20076 22484 20132 22876
rect 20076 22428 20244 22484
rect 19404 22148 19460 22428
rect 20188 22370 20244 22428
rect 20188 22318 20190 22370
rect 20242 22318 20244 22370
rect 20188 22306 20244 22318
rect 19516 22260 19572 22270
rect 19516 22166 19572 22204
rect 20076 22258 20132 22270
rect 20076 22206 20078 22258
rect 20130 22206 20132 22258
rect 20076 22148 20132 22206
rect 20300 22260 20356 23772
rect 20524 23716 20580 23726
rect 20412 22708 20468 22718
rect 20412 22482 20468 22652
rect 20412 22430 20414 22482
rect 20466 22430 20468 22482
rect 20412 22418 20468 22430
rect 20524 22260 20580 23660
rect 21196 22708 21252 26796
rect 21420 26786 21476 26796
rect 21868 26514 21924 26908
rect 22316 26908 22372 28588
rect 25228 28420 25284 37998
rect 25564 37156 25620 41200
rect 26124 38612 26180 38622
rect 26124 38274 26180 38556
rect 26124 38222 26126 38274
rect 26178 38222 26180 38274
rect 26124 38210 26180 38222
rect 26236 38276 26292 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 26236 38210 26292 38220
rect 29372 38276 29428 38286
rect 29372 38182 29428 38220
rect 28588 38050 28644 38062
rect 28588 37998 28590 38050
rect 28642 37998 28644 38050
rect 28252 37266 28308 37278
rect 28252 37214 28254 37266
rect 28306 37214 28308 37266
rect 26012 37156 26068 37166
rect 25564 37154 26068 37156
rect 25564 37102 26014 37154
rect 26066 37102 26068 37154
rect 25564 37100 26068 37102
rect 26012 37090 26068 37100
rect 25004 28364 25284 28420
rect 22764 27748 22820 27758
rect 22764 27654 22820 27692
rect 24220 27188 24276 27198
rect 22876 26964 22932 26974
rect 22876 26962 23156 26964
rect 22876 26910 22878 26962
rect 22930 26910 23156 26962
rect 22876 26908 23156 26910
rect 22316 26852 22484 26908
rect 22876 26898 22932 26908
rect 21868 26462 21870 26514
rect 21922 26462 21924 26514
rect 21868 26450 21924 26462
rect 21420 26180 21476 26190
rect 21420 26178 21588 26180
rect 21420 26126 21422 26178
rect 21474 26126 21588 26178
rect 21420 26124 21588 26126
rect 21420 26114 21476 26124
rect 21420 24722 21476 24734
rect 21420 24670 21422 24722
rect 21474 24670 21476 24722
rect 21420 24276 21476 24670
rect 21420 24210 21476 24220
rect 21532 24500 21588 26124
rect 21980 25396 22036 25406
rect 21980 24946 22036 25340
rect 21980 24894 21982 24946
rect 22034 24894 22036 24946
rect 21980 24882 22036 24894
rect 22092 25284 22148 25294
rect 21644 24500 21700 24510
rect 21532 24498 21700 24500
rect 21532 24446 21646 24498
rect 21698 24446 21700 24498
rect 21532 24444 21700 24446
rect 21308 23940 21364 23950
rect 21308 23846 21364 23884
rect 21420 23828 21476 23838
rect 21532 23828 21588 24444
rect 21644 24434 21700 24444
rect 21868 24052 21924 24062
rect 21476 23772 21588 23828
rect 21644 23826 21700 23838
rect 21644 23774 21646 23826
rect 21698 23774 21700 23826
rect 21420 23762 21476 23772
rect 21196 22642 21252 22652
rect 21420 22820 21476 22830
rect 21644 22820 21700 23774
rect 21868 23714 21924 23996
rect 21868 23662 21870 23714
rect 21922 23662 21924 23714
rect 21868 23650 21924 23662
rect 22092 23492 22148 25228
rect 22204 23828 22260 23838
rect 22204 23734 22260 23772
rect 22092 23266 22148 23436
rect 22428 23380 22484 26852
rect 23100 26514 23156 26908
rect 23100 26462 23102 26514
rect 23154 26462 23156 26514
rect 23100 26450 23156 26462
rect 24220 26402 24276 27132
rect 25004 27188 25060 28364
rect 25004 27094 25060 27132
rect 25452 27748 25508 27758
rect 25900 27748 25956 27758
rect 25508 27746 25956 27748
rect 25508 27694 25902 27746
rect 25954 27694 25956 27746
rect 25508 27692 25956 27694
rect 25452 27074 25508 27692
rect 25900 27682 25956 27692
rect 25452 27022 25454 27074
rect 25506 27022 25508 27074
rect 24220 26350 24222 26402
rect 24274 26350 24276 26402
rect 24220 26338 24276 26350
rect 24780 26964 24836 26974
rect 22988 26292 23044 26302
rect 22988 26198 23044 26236
rect 23212 26290 23268 26302
rect 23212 26238 23214 26290
rect 23266 26238 23268 26290
rect 22092 23214 22094 23266
rect 22146 23214 22148 23266
rect 22092 23202 22148 23214
rect 22204 23324 22484 23380
rect 23100 25844 23156 25854
rect 23100 25396 23156 25788
rect 21644 22764 21924 22820
rect 20300 22204 20468 22260
rect 20076 22092 20244 22148
rect 19404 22036 19460 22092
rect 19628 22036 19684 22046
rect 19404 21980 19572 22036
rect 19516 21700 19572 21980
rect 19628 21812 19684 21980
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19964 21812 20020 21822
rect 20188 21812 20244 22092
rect 19628 21810 20020 21812
rect 19628 21758 19966 21810
rect 20018 21758 20020 21810
rect 19628 21756 20020 21758
rect 19964 21746 20020 21756
rect 20076 21756 20244 21812
rect 19516 21698 19684 21700
rect 19516 21646 19518 21698
rect 19570 21646 19684 21698
rect 19516 21644 19684 21646
rect 19516 21634 19572 21644
rect 19404 21586 19460 21598
rect 19404 21534 19406 21586
rect 19458 21534 19460 21586
rect 18732 20526 18734 20578
rect 18786 20526 18788 20578
rect 18508 20020 18564 20030
rect 18508 19926 18564 19964
rect 18172 19842 18228 19852
rect 18732 19796 18788 20526
rect 18508 19740 18788 19796
rect 18844 20748 19012 20804
rect 19068 21140 19124 21150
rect 18172 19348 18228 19358
rect 18172 19236 18228 19292
rect 18396 19236 18452 19246
rect 18172 19234 18452 19236
rect 18172 19182 18398 19234
rect 18450 19182 18452 19234
rect 18172 19180 18452 19182
rect 18396 19170 18452 19180
rect 18508 19124 18564 19740
rect 18620 19460 18676 19470
rect 18620 19346 18676 19404
rect 18620 19294 18622 19346
rect 18674 19294 18676 19346
rect 18620 19282 18676 19294
rect 18732 19236 18788 19246
rect 18732 19142 18788 19180
rect 18060 19068 18340 19124
rect 18508 19068 18676 19124
rect 17948 18956 18116 19012
rect 17612 18732 17892 18788
rect 17724 18564 17780 18574
rect 17164 17556 17220 17566
rect 17164 17462 17220 17500
rect 16828 17108 16884 17118
rect 16772 17106 16884 17108
rect 16772 17054 16830 17106
rect 16882 17054 16884 17106
rect 16772 17052 16884 17054
rect 16716 17014 16772 17052
rect 16828 17042 16884 17052
rect 16268 16996 16324 17006
rect 17276 16996 17332 18060
rect 17388 18562 17780 18564
rect 17388 18510 17726 18562
rect 17778 18510 17780 18562
rect 17388 18508 17780 18510
rect 17388 17666 17444 18508
rect 17724 18498 17780 18508
rect 17836 18564 17892 18732
rect 18060 18564 18116 18956
rect 17836 18562 18004 18564
rect 17836 18510 17838 18562
rect 17890 18510 18004 18562
rect 17836 18508 18004 18510
rect 17836 18498 17892 18508
rect 17724 18228 17780 18238
rect 17948 18228 18004 18508
rect 18060 18498 18116 18508
rect 18172 18562 18228 18574
rect 18172 18510 18174 18562
rect 18226 18510 18228 18562
rect 18060 18228 18116 18238
rect 17724 18226 17892 18228
rect 17724 18174 17726 18226
rect 17778 18174 17892 18226
rect 17724 18172 17892 18174
rect 17948 18172 18060 18228
rect 17724 18162 17780 18172
rect 17388 17614 17390 17666
rect 17442 17614 17444 17666
rect 17388 17602 17444 17614
rect 17724 17666 17780 17678
rect 17724 17614 17726 17666
rect 17778 17614 17780 17666
rect 17500 17554 17556 17566
rect 17500 17502 17502 17554
rect 17554 17502 17556 17554
rect 17500 17444 17556 17502
rect 17724 17556 17780 17614
rect 17724 17490 17780 17500
rect 17500 17378 17556 17388
rect 17388 16996 17444 17006
rect 17276 16994 17444 16996
rect 17276 16942 17390 16994
rect 17442 16942 17444 16994
rect 17276 16940 17444 16942
rect 16268 16902 16324 16940
rect 17388 16930 17444 16940
rect 17724 16996 17780 17006
rect 17836 16996 17892 18172
rect 18060 18162 18116 18172
rect 18172 17780 18228 18510
rect 18172 17714 18228 17724
rect 17948 17666 18004 17678
rect 17948 17614 17950 17666
rect 18002 17614 18004 17666
rect 17948 17556 18004 17614
rect 18284 17556 18340 19068
rect 17948 17500 18340 17556
rect 18396 19012 18452 19022
rect 18396 17780 18452 18956
rect 18508 18452 18564 18462
rect 18620 18452 18676 19068
rect 18844 19012 18900 20748
rect 18564 18396 18676 18452
rect 18732 18956 18900 19012
rect 18956 20580 19012 20590
rect 18508 18358 18564 18396
rect 18732 18004 18788 18956
rect 18844 18228 18900 18238
rect 18844 18134 18900 18172
rect 18956 18116 19012 20524
rect 19068 19234 19124 21084
rect 19180 21028 19236 21038
rect 19180 20934 19236 20972
rect 19292 20804 19348 20814
rect 19292 20710 19348 20748
rect 19292 20356 19348 20366
rect 19068 19182 19070 19234
rect 19122 19182 19124 19234
rect 19068 19170 19124 19182
rect 19180 20244 19236 20254
rect 19180 18452 19236 20188
rect 19068 18450 19236 18452
rect 19068 18398 19182 18450
rect 19234 18398 19236 18450
rect 19068 18396 19236 18398
rect 19068 18340 19124 18396
rect 19180 18386 19236 18396
rect 19292 19346 19348 20300
rect 19292 19294 19294 19346
rect 19346 19294 19348 19346
rect 19292 18340 19348 19294
rect 19404 19236 19460 21534
rect 19516 21364 19572 21374
rect 19516 21270 19572 21308
rect 19404 19142 19460 19180
rect 19628 18676 19684 21644
rect 20076 21140 20132 21756
rect 20076 21074 20132 21084
rect 20188 20916 20244 20926
rect 19852 20804 19908 20814
rect 19852 20710 19908 20748
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19740 20020 19796 20030
rect 19740 19926 19796 19964
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 18620 19908 18676
rect 19516 18562 19572 18574
rect 19516 18510 19518 18562
rect 19570 18510 19572 18562
rect 19516 18340 19572 18510
rect 19292 18284 19460 18340
rect 19068 18274 19124 18284
rect 19180 18228 19236 18238
rect 19180 18226 19348 18228
rect 19180 18174 19182 18226
rect 19234 18174 19348 18226
rect 19180 18172 19348 18174
rect 19180 18162 19236 18172
rect 18956 18060 19124 18116
rect 18732 17948 18900 18004
rect 18396 17666 18452 17724
rect 18508 17780 18564 17790
rect 18508 17778 18788 17780
rect 18508 17726 18510 17778
rect 18562 17726 18788 17778
rect 18508 17724 18788 17726
rect 18508 17714 18564 17724
rect 18396 17614 18398 17666
rect 18450 17614 18452 17666
rect 17948 16996 18004 17006
rect 18396 16996 18452 17614
rect 18620 17556 18676 17566
rect 18620 17462 18676 17500
rect 17836 16994 18340 16996
rect 17836 16942 17950 16994
rect 18002 16942 18340 16994
rect 17836 16940 18340 16942
rect 15708 16830 15710 16882
rect 15762 16830 15764 16882
rect 15708 16818 15764 16830
rect 16156 16882 16212 16894
rect 16156 16830 16158 16882
rect 16210 16830 16212 16882
rect 14924 16098 15092 16100
rect 14924 16046 14926 16098
rect 14978 16046 15092 16098
rect 14924 16044 15092 16046
rect 15148 16772 15204 16782
rect 14924 16034 14980 16044
rect 15148 15986 15204 16716
rect 15148 15934 15150 15986
rect 15202 15934 15204 15986
rect 15148 15922 15204 15934
rect 15260 15988 15316 15998
rect 15260 15894 15316 15932
rect 15596 15988 15652 15998
rect 14588 15876 14644 15886
rect 14588 15782 14644 15820
rect 13356 15374 13358 15426
rect 13410 15374 13412 15426
rect 13356 15362 13412 15374
rect 14140 15596 14644 15652
rect 14140 15314 14196 15596
rect 14140 15262 14142 15314
rect 14194 15262 14196 15314
rect 14140 15250 14196 15262
rect 14588 15538 14644 15596
rect 14588 15486 14590 15538
rect 14642 15486 14644 15538
rect 11228 15150 11230 15202
rect 11282 15150 11284 15202
rect 11228 15138 11284 15150
rect 13580 15092 13636 15102
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 13580 13746 13636 15036
rect 14588 15092 14644 15486
rect 14588 15026 14644 15036
rect 15596 14530 15652 15932
rect 16156 15988 16212 16830
rect 17724 16882 17780 16940
rect 17948 16930 18004 16940
rect 17724 16830 17726 16882
rect 17778 16830 17780 16882
rect 17724 16818 17780 16830
rect 17836 16772 17892 16782
rect 17836 16678 17892 16716
rect 17164 16100 17220 16110
rect 17164 16006 17220 16044
rect 16156 15922 16212 15932
rect 16828 15988 16884 15998
rect 16828 15894 16884 15932
rect 18172 15876 18228 15886
rect 18172 15426 18228 15820
rect 18172 15374 18174 15426
rect 18226 15374 18228 15426
rect 18172 15362 18228 15374
rect 15596 14478 15598 14530
rect 15650 14478 15652 14530
rect 15596 14466 15652 14478
rect 16156 15092 16212 15102
rect 18060 15092 18116 15102
rect 16156 14532 16212 15036
rect 16940 15090 18116 15092
rect 16940 15038 18062 15090
rect 18114 15038 18116 15090
rect 16940 15036 18116 15038
rect 16940 14642 16996 15036
rect 18060 15026 18116 15036
rect 16940 14590 16942 14642
rect 16994 14590 16996 14642
rect 16940 14578 16996 14590
rect 16156 14530 16772 14532
rect 16156 14478 16158 14530
rect 16210 14478 16772 14530
rect 16156 14476 16772 14478
rect 16156 14466 16212 14476
rect 13580 13694 13582 13746
rect 13634 13694 13636 13746
rect 13580 13682 13636 13694
rect 15708 14306 15764 14318
rect 15708 14254 15710 14306
rect 15762 14254 15764 14306
rect 14364 13634 14420 13646
rect 14364 13582 14366 13634
rect 14418 13582 14420 13634
rect 14364 13524 14420 13582
rect 15708 13636 15764 14254
rect 15932 14308 15988 14318
rect 15932 14214 15988 14252
rect 15708 13570 15764 13580
rect 16492 13636 16548 13646
rect 16492 13542 16548 13580
rect 14364 13458 14420 13468
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 16716 13076 16772 14476
rect 17388 14308 17444 14318
rect 17388 13858 17444 14252
rect 17388 13806 17390 13858
rect 17442 13806 17444 13858
rect 17388 13794 17444 13806
rect 17948 13860 18004 13870
rect 17612 13748 17668 13758
rect 17612 13654 17668 13692
rect 17948 13746 18004 13804
rect 17948 13694 17950 13746
rect 18002 13694 18004 13746
rect 17948 13682 18004 13694
rect 18172 13748 18228 13758
rect 18284 13748 18340 16940
rect 18396 16930 18452 16940
rect 18508 17108 18564 17118
rect 18508 16994 18564 17052
rect 18508 16942 18510 16994
rect 18562 16942 18564 16994
rect 18508 16930 18564 16942
rect 18732 16660 18788 17724
rect 18732 16594 18788 16604
rect 18620 15986 18676 15998
rect 18620 15934 18622 15986
rect 18674 15934 18676 15986
rect 18620 14644 18676 15934
rect 18844 15148 18900 17948
rect 18956 17892 19012 17902
rect 18956 17666 19012 17836
rect 18956 17614 18958 17666
rect 19010 17614 19012 17666
rect 18956 17602 19012 17614
rect 19068 17556 19124 18060
rect 19068 17490 19124 17500
rect 19068 16772 19124 16782
rect 19068 16322 19124 16716
rect 19068 16270 19070 16322
rect 19122 16270 19124 16322
rect 19068 16258 19124 16270
rect 19292 16212 19348 18172
rect 18956 16100 19012 16138
rect 19292 16118 19348 16156
rect 19012 16044 19124 16100
rect 18956 16034 19012 16044
rect 19068 15988 19124 16044
rect 19404 15988 19460 18284
rect 19516 18116 19572 18284
rect 19516 18050 19572 18060
rect 19740 18452 19796 18462
rect 19516 17780 19572 17790
rect 19516 17666 19572 17724
rect 19516 17614 19518 17666
rect 19570 17614 19572 17666
rect 19516 17602 19572 17614
rect 19740 17666 19796 18396
rect 19852 18450 19908 18620
rect 19852 18398 19854 18450
rect 19906 18398 19908 18450
rect 19852 18386 19908 18398
rect 19740 17614 19742 17666
rect 19794 17614 19796 17666
rect 19740 17602 19796 17614
rect 19628 17442 19684 17454
rect 19628 17390 19630 17442
rect 19682 17390 19684 17442
rect 19516 17332 19572 17342
rect 19516 16660 19572 17276
rect 19516 16098 19572 16604
rect 19516 16046 19518 16098
rect 19570 16046 19572 16098
rect 19516 16034 19572 16046
rect 19068 15932 19460 15988
rect 18956 15876 19012 15886
rect 18956 15782 19012 15820
rect 19628 15876 19684 17390
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 15810 19684 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20188 15316 20244 20860
rect 20300 19346 20356 19358
rect 20300 19294 20302 19346
rect 20354 19294 20356 19346
rect 20300 19236 20356 19294
rect 20300 19170 20356 19180
rect 20412 18564 20468 22204
rect 20524 22194 20580 22204
rect 21308 22260 21364 22270
rect 21308 22166 21364 22204
rect 21420 21924 21476 22764
rect 21756 22596 21812 22606
rect 21644 22484 21700 22494
rect 21420 21858 21476 21868
rect 21532 22146 21588 22158
rect 21532 22094 21534 22146
rect 21586 22094 21588 22146
rect 20972 21698 21028 21710
rect 20972 21646 20974 21698
rect 21026 21646 21028 21698
rect 20860 21586 20916 21598
rect 20860 21534 20862 21586
rect 20914 21534 20916 21586
rect 20524 21474 20580 21486
rect 20524 21422 20526 21474
rect 20578 21422 20580 21474
rect 20524 19348 20580 21422
rect 20860 19460 20916 21534
rect 20972 20916 21028 21646
rect 20972 20850 21028 20860
rect 21532 20804 21588 22094
rect 21644 21810 21700 22428
rect 21756 22482 21812 22540
rect 21756 22430 21758 22482
rect 21810 22430 21812 22482
rect 21756 22418 21812 22430
rect 21868 22372 21924 22764
rect 22092 22372 22148 22382
rect 21868 22370 22148 22372
rect 21868 22318 22094 22370
rect 22146 22318 22148 22370
rect 21868 22316 22148 22318
rect 21756 22146 21812 22158
rect 21756 22094 21758 22146
rect 21810 22094 21812 22146
rect 21756 21924 21812 22094
rect 21756 21858 21812 21868
rect 21644 21758 21646 21810
rect 21698 21758 21700 21810
rect 21644 21746 21700 21758
rect 21532 20738 21588 20748
rect 21756 21698 21812 21710
rect 21756 21646 21758 21698
rect 21810 21646 21812 21698
rect 21756 20802 21812 21646
rect 21868 21028 21924 22316
rect 22092 22306 22148 22316
rect 22204 22148 22260 23324
rect 21868 20962 21924 20972
rect 21980 22146 22260 22148
rect 21980 22094 22206 22146
rect 22258 22094 22260 22146
rect 21980 22092 22260 22094
rect 21756 20750 21758 20802
rect 21810 20750 21812 20802
rect 21756 20244 21812 20750
rect 21756 20178 21812 20188
rect 20860 19394 20916 19404
rect 20524 19282 20580 19292
rect 21868 19236 21924 19246
rect 20748 19012 20804 19022
rect 20412 18498 20468 18508
rect 20524 19010 21140 19012
rect 20524 18958 20750 19010
rect 20802 18958 21140 19010
rect 20524 18956 21140 18958
rect 20300 18450 20356 18462
rect 20300 18398 20302 18450
rect 20354 18398 20356 18450
rect 20300 18340 20356 18398
rect 20524 18340 20580 18956
rect 20748 18946 20804 18956
rect 21084 18674 21140 18956
rect 21084 18622 21086 18674
rect 21138 18622 21140 18674
rect 21084 18610 21140 18622
rect 21196 18564 21252 18574
rect 21196 18450 21252 18508
rect 21196 18398 21198 18450
rect 21250 18398 21252 18450
rect 21196 18386 21252 18398
rect 21756 18452 21812 18462
rect 21756 18358 21812 18396
rect 20300 18284 20580 18340
rect 20748 18338 20804 18350
rect 20748 18286 20750 18338
rect 20802 18286 20804 18338
rect 20748 18004 20804 18286
rect 20748 17938 20804 17948
rect 20412 17892 20468 17902
rect 20300 15316 20356 15326
rect 20188 15260 20300 15316
rect 20300 15250 20356 15260
rect 18844 15092 19236 15148
rect 19068 14644 19124 14654
rect 18620 14642 19124 14644
rect 18620 14590 19070 14642
rect 19122 14590 19124 14642
rect 18620 14588 19124 14590
rect 18172 13746 18340 13748
rect 18172 13694 18174 13746
rect 18226 13694 18340 13746
rect 18172 13692 18340 13694
rect 18172 13682 18228 13692
rect 16716 12982 16772 13020
rect 16940 13636 16996 13646
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 16940 3554 16996 13580
rect 17500 13524 17556 13534
rect 17500 13430 17556 13468
rect 17724 13076 17780 13086
rect 17724 12962 17780 13020
rect 17724 12910 17726 12962
rect 17778 12910 17780 12962
rect 17724 12898 17780 12910
rect 18508 12852 18564 12862
rect 18508 12758 18564 12796
rect 19068 4338 19124 14588
rect 19180 13860 19236 15092
rect 19516 14644 19572 14654
rect 19516 14550 19572 14588
rect 20300 14532 20356 14542
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19404 13860 19460 13870
rect 19236 13858 19460 13860
rect 19236 13806 19406 13858
rect 19458 13806 19460 13858
rect 19236 13804 19460 13806
rect 19180 13766 19236 13804
rect 19404 13794 19460 13804
rect 19516 13860 19572 13870
rect 19516 13766 19572 13804
rect 19740 13858 19796 13870
rect 19740 13806 19742 13858
rect 19794 13806 19796 13858
rect 19740 13748 19796 13806
rect 20300 13858 20356 14476
rect 20300 13806 20302 13858
rect 20354 13806 20356 13858
rect 20300 13794 20356 13806
rect 19852 13748 19908 13758
rect 19740 13746 19908 13748
rect 19740 13694 19854 13746
rect 19906 13694 19908 13746
rect 19740 13692 19908 13694
rect 19852 13682 19908 13692
rect 20412 13748 20468 17836
rect 21868 17554 21924 19180
rect 21868 17502 21870 17554
rect 21922 17502 21924 17554
rect 21868 17490 21924 17502
rect 21980 18452 22036 22092
rect 22204 22082 22260 22092
rect 22428 23156 22484 23166
rect 22204 20802 22260 20814
rect 22204 20750 22206 20802
rect 22258 20750 22260 20802
rect 22204 18676 22260 20750
rect 22204 18610 22260 18620
rect 22316 19908 22372 19918
rect 22428 19908 22484 23100
rect 22988 22708 23044 22718
rect 22988 21698 23044 22652
rect 22988 21646 22990 21698
rect 23042 21646 23044 21698
rect 22876 21588 22932 21598
rect 22876 21494 22932 21532
rect 22316 19906 22484 19908
rect 22316 19854 22318 19906
rect 22370 19854 22484 19906
rect 22316 19852 22484 19854
rect 22540 21028 22596 21038
rect 21980 17444 22036 18396
rect 20524 16212 20580 16222
rect 20524 16098 20580 16156
rect 20524 16046 20526 16098
rect 20578 16046 20580 16098
rect 20524 16034 20580 16046
rect 21196 16212 21252 16222
rect 21196 16098 21252 16156
rect 21196 16046 21198 16098
rect 21250 16046 21252 16098
rect 21196 16034 21252 16046
rect 21868 16100 21924 16110
rect 21980 16100 22036 17388
rect 22316 16882 22372 19852
rect 22428 18564 22484 18574
rect 22540 18564 22596 20972
rect 22764 20690 22820 20702
rect 22764 20638 22766 20690
rect 22818 20638 22820 20690
rect 22764 20244 22820 20638
rect 22764 20178 22820 20188
rect 22988 20132 23044 21646
rect 23100 22258 23156 25340
rect 23212 24052 23268 26238
rect 23548 26292 23604 26302
rect 23548 26290 23828 26292
rect 23548 26238 23550 26290
rect 23602 26238 23828 26290
rect 23548 26236 23828 26238
rect 23548 26226 23604 26236
rect 23212 23986 23268 23996
rect 23772 25620 23828 26236
rect 23884 26290 23940 26302
rect 23884 26238 23886 26290
rect 23938 26238 23940 26290
rect 23884 26180 23940 26238
rect 23996 26292 24052 26302
rect 23996 26198 24052 26236
rect 24444 26292 24500 26302
rect 24668 26292 24724 26302
rect 24444 26290 24668 26292
rect 24444 26238 24446 26290
rect 24498 26238 24668 26290
rect 24444 26236 24668 26238
rect 24444 26226 24500 26236
rect 23884 25844 23940 26124
rect 23884 25778 23940 25788
rect 23772 25564 24612 25620
rect 23100 22206 23102 22258
rect 23154 22206 23156 22258
rect 23100 21700 23156 22206
rect 23100 21634 23156 21644
rect 23436 23828 23492 23838
rect 23324 20916 23380 20926
rect 23324 20822 23380 20860
rect 22988 20066 23044 20076
rect 23100 20802 23156 20814
rect 23100 20750 23102 20802
rect 23154 20750 23156 20802
rect 23100 19122 23156 20750
rect 23436 20188 23492 23772
rect 23772 21812 23828 25564
rect 24556 25506 24612 25564
rect 24556 25454 24558 25506
rect 24610 25454 24612 25506
rect 24556 25442 24612 25454
rect 24668 25396 24724 26236
rect 24780 25618 24836 26908
rect 25116 26290 25172 26302
rect 25116 26238 25118 26290
rect 25170 26238 25172 26290
rect 25116 26180 25172 26238
rect 25116 26114 25172 26124
rect 25340 26178 25396 26190
rect 25340 26126 25342 26178
rect 25394 26126 25396 26178
rect 25340 25844 25396 26126
rect 24892 25788 25396 25844
rect 24892 25730 24948 25788
rect 24892 25678 24894 25730
rect 24946 25678 24948 25730
rect 24892 25666 24948 25678
rect 24780 25566 24782 25618
rect 24834 25566 24836 25618
rect 24780 25554 24836 25566
rect 24668 25340 24836 25396
rect 23884 22370 23940 22382
rect 23884 22318 23886 22370
rect 23938 22318 23940 22370
rect 23884 21924 23940 22318
rect 23884 21858 23940 21868
rect 23772 21718 23828 21756
rect 23548 21698 23604 21710
rect 24668 21700 24724 21710
rect 23548 21646 23550 21698
rect 23602 21646 23604 21698
rect 23548 21364 23604 21646
rect 24444 21698 24724 21700
rect 24444 21646 24670 21698
rect 24722 21646 24724 21698
rect 24444 21644 24724 21646
rect 23548 20356 23604 21308
rect 24332 21586 24388 21598
rect 24332 21534 24334 21586
rect 24386 21534 24388 21586
rect 24332 21028 24388 21534
rect 24332 20962 24388 20972
rect 23660 20804 23716 20814
rect 23660 20710 23716 20748
rect 24220 20802 24276 20814
rect 24220 20750 24222 20802
rect 24274 20750 24276 20802
rect 23548 20290 23604 20300
rect 23436 20132 23716 20188
rect 23660 20020 23716 20132
rect 23100 19070 23102 19122
rect 23154 19070 23156 19122
rect 22428 18562 22596 18564
rect 22428 18510 22430 18562
rect 22482 18510 22596 18562
rect 22428 18508 22596 18510
rect 22988 18564 23044 18574
rect 22428 18498 22484 18508
rect 22988 18470 23044 18508
rect 23100 18450 23156 19070
rect 23100 18398 23102 18450
rect 23154 18398 23156 18450
rect 23100 18004 23156 18398
rect 23436 19348 23492 19358
rect 23436 19236 23492 19292
rect 23548 19236 23604 19246
rect 23436 19234 23604 19236
rect 23436 19182 23550 19234
rect 23602 19182 23604 19234
rect 23436 19180 23604 19182
rect 23324 18340 23380 18350
rect 23100 17938 23156 17948
rect 23212 18338 23380 18340
rect 23212 18286 23326 18338
rect 23378 18286 23380 18338
rect 23212 18284 23380 18286
rect 22316 16830 22318 16882
rect 22370 16830 22372 16882
rect 22316 16818 22372 16830
rect 23100 16324 23156 16334
rect 22764 16322 23156 16324
rect 22764 16270 23102 16322
rect 23154 16270 23156 16322
rect 22764 16268 23156 16270
rect 21868 16098 22036 16100
rect 21868 16046 21870 16098
rect 21922 16046 22036 16098
rect 21868 16044 22036 16046
rect 22652 16100 22708 16110
rect 22764 16100 22820 16268
rect 23100 16258 23156 16268
rect 22652 16098 22820 16100
rect 22652 16046 22654 16098
rect 22706 16046 22820 16098
rect 22652 16044 22820 16046
rect 22876 16100 22932 16110
rect 21868 16034 21924 16044
rect 22652 16034 22708 16044
rect 21644 15986 21700 15998
rect 21644 15934 21646 15986
rect 21698 15934 21700 15986
rect 20636 15876 20692 15886
rect 20860 15876 20916 15886
rect 20692 15820 20804 15876
rect 20636 15782 20692 15820
rect 20748 15428 20804 15820
rect 20860 15874 21252 15876
rect 20860 15822 20862 15874
rect 20914 15822 21252 15874
rect 20860 15820 21252 15822
rect 20860 15810 20916 15820
rect 21196 15540 21252 15820
rect 21532 15874 21588 15886
rect 21532 15822 21534 15874
rect 21586 15822 21588 15874
rect 21532 15652 21588 15822
rect 21644 15876 21700 15934
rect 22876 15986 22932 16044
rect 22876 15934 22878 15986
rect 22930 15934 22932 15986
rect 21644 15810 21700 15820
rect 22428 15876 22484 15886
rect 21532 15596 22036 15652
rect 21420 15540 21476 15550
rect 21196 15538 21476 15540
rect 21196 15486 21422 15538
rect 21474 15486 21476 15538
rect 21196 15484 21476 15486
rect 21420 15474 21476 15484
rect 20748 15372 21028 15428
rect 20972 15314 21028 15372
rect 21980 15426 22036 15596
rect 22428 15540 22484 15820
rect 22540 15540 22596 15550
rect 22428 15538 22596 15540
rect 22428 15486 22542 15538
rect 22594 15486 22596 15538
rect 22428 15484 22596 15486
rect 22540 15474 22596 15484
rect 21980 15374 21982 15426
rect 22034 15374 22036 15426
rect 21980 15362 22036 15374
rect 20972 15262 20974 15314
rect 21026 15262 21028 15314
rect 20972 15250 21028 15262
rect 21196 15316 21252 15326
rect 21196 15222 21252 15260
rect 21644 15314 21700 15326
rect 21644 15262 21646 15314
rect 21698 15262 21700 15314
rect 21308 15202 21364 15214
rect 21308 15150 21310 15202
rect 21362 15150 21364 15202
rect 21308 14196 21364 15150
rect 21644 14756 21700 15262
rect 22204 15314 22260 15326
rect 22204 15262 22206 15314
rect 22258 15262 22260 15314
rect 22204 14868 22260 15262
rect 22428 15316 22484 15326
rect 22428 15222 22484 15260
rect 22204 14802 22260 14812
rect 22316 15202 22372 15214
rect 22316 15150 22318 15202
rect 22370 15150 22372 15202
rect 21644 14690 21700 14700
rect 21308 14130 21364 14140
rect 21868 14644 21924 14654
rect 20972 13972 21028 13982
rect 21420 13972 21476 13982
rect 21868 13972 21924 14588
rect 20972 13970 21924 13972
rect 20972 13918 20974 13970
rect 21026 13918 21422 13970
rect 21474 13918 21924 13970
rect 20972 13916 21924 13918
rect 20972 13906 21028 13916
rect 20412 13654 20468 13692
rect 20636 13860 20692 13870
rect 20076 13634 20132 13646
rect 20076 13582 20078 13634
rect 20130 13582 20132 13634
rect 20076 12852 20132 13582
rect 20636 13076 20692 13804
rect 20636 13074 20804 13076
rect 20636 13022 20638 13074
rect 20690 13022 20804 13074
rect 20636 13020 20804 13022
rect 20636 13010 20692 13020
rect 20076 12786 20132 12796
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19068 4286 19070 4338
rect 19122 4286 19124 4338
rect 19068 4274 19124 4286
rect 16940 3502 16942 3554
rect 16994 3502 16996 3554
rect 16940 3490 16996 3502
rect 18844 4116 18900 4126
rect 16156 3444 16212 3454
rect 16156 800 16212 3388
rect 18508 3444 18564 3454
rect 18508 3350 18564 3388
rect 18844 800 18900 4060
rect 20076 4116 20132 4126
rect 20076 4022 20132 4060
rect 20748 3554 20804 13020
rect 21084 12402 21140 13916
rect 21420 12962 21476 13916
rect 21868 13746 21924 13916
rect 21868 13694 21870 13746
rect 21922 13694 21924 13746
rect 21868 13682 21924 13694
rect 22092 14196 22148 14206
rect 22092 13074 22148 14140
rect 22316 13860 22372 15150
rect 22876 15148 22932 15934
rect 22764 15092 22932 15148
rect 22652 14756 22708 14766
rect 22652 14662 22708 14700
rect 22540 14532 22596 14542
rect 22540 14438 22596 14476
rect 22764 14530 22820 15092
rect 22764 14478 22766 14530
rect 22818 14478 22820 14530
rect 22764 14466 22820 14478
rect 23212 14532 23268 18284
rect 23324 18274 23380 18284
rect 23324 17668 23380 17678
rect 23436 17668 23492 19180
rect 23548 19170 23604 19180
rect 23660 19124 23716 19964
rect 23996 19236 24052 19246
rect 23660 19058 23716 19068
rect 23772 19234 24052 19236
rect 23772 19182 23998 19234
rect 24050 19182 24052 19234
rect 23772 19180 24052 19182
rect 23324 17666 23492 17668
rect 23324 17614 23326 17666
rect 23378 17614 23492 17666
rect 23324 17612 23492 17614
rect 23548 18452 23604 18462
rect 23324 16322 23380 17612
rect 23548 16884 23604 18396
rect 23772 18228 23828 19180
rect 23996 19170 24052 19180
rect 24108 18452 24164 18462
rect 24108 18358 24164 18396
rect 24220 18340 24276 20750
rect 24444 20580 24500 21644
rect 24668 21634 24724 21644
rect 24780 21476 24836 25340
rect 25340 23716 25396 23726
rect 25452 23716 25508 27022
rect 28252 27186 28308 37214
rect 28252 27134 28254 27186
rect 28306 27134 28308 27186
rect 26124 26964 26180 26974
rect 26124 26870 26180 26908
rect 26236 26852 26292 26862
rect 25564 26404 25620 26414
rect 25564 26310 25620 26348
rect 26236 26404 26292 26796
rect 28252 26852 28308 27134
rect 28252 26786 28308 26796
rect 26460 26516 26516 26526
rect 26460 26422 26516 26460
rect 28588 26516 28644 37998
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 28588 26450 28644 26460
rect 25676 26292 25732 26302
rect 25676 26198 25732 26236
rect 26236 26290 26292 26348
rect 26236 26238 26238 26290
rect 26290 26238 26292 26290
rect 26236 26226 26292 26238
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 27020 24052 27076 24062
rect 25676 23938 25732 23950
rect 25676 23886 25678 23938
rect 25730 23886 25732 23938
rect 25676 23716 25732 23886
rect 25340 23714 25732 23716
rect 25340 23662 25342 23714
rect 25394 23662 25732 23714
rect 25340 23660 25732 23662
rect 26460 23826 26516 23838
rect 26460 23774 26462 23826
rect 26514 23774 26516 23826
rect 25340 23492 25396 23660
rect 25228 23436 25340 23492
rect 25228 22372 25284 23436
rect 25340 23426 25396 23436
rect 26460 23378 26516 23774
rect 26460 23326 26462 23378
rect 26514 23326 26516 23378
rect 26460 23314 26516 23326
rect 27020 23378 27076 23996
rect 28588 24052 28644 24062
rect 28588 23958 28644 23996
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 37660 23940 37716 23950
rect 37660 23846 37716 23884
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 27020 23326 27022 23378
rect 27074 23326 27076 23378
rect 27020 23314 27076 23326
rect 25452 23266 25508 23278
rect 25452 23214 25454 23266
rect 25506 23214 25508 23266
rect 25340 23154 25396 23166
rect 25340 23102 25342 23154
rect 25394 23102 25396 23154
rect 25340 22596 25396 23102
rect 25340 22530 25396 22540
rect 25340 22372 25396 22382
rect 25228 22370 25396 22372
rect 25228 22318 25342 22370
rect 25394 22318 25396 22370
rect 25228 22316 25396 22318
rect 25116 21924 25172 21934
rect 24668 21420 24836 21476
rect 24892 21588 24948 21598
rect 24556 21140 24612 21150
rect 24556 20802 24612 21084
rect 24556 20750 24558 20802
rect 24610 20750 24612 20802
rect 24556 20738 24612 20750
rect 24556 20580 24612 20590
rect 24444 20524 24556 20580
rect 24556 20514 24612 20524
rect 24556 20356 24612 20366
rect 24556 20242 24612 20300
rect 24556 20190 24558 20242
rect 24610 20190 24612 20242
rect 24556 20178 24612 20190
rect 24444 20132 24500 20142
rect 24444 20038 24500 20076
rect 24668 19346 24724 21420
rect 24892 20692 24948 21532
rect 25116 20804 25172 21868
rect 25228 20916 25284 22316
rect 25340 22306 25396 22316
rect 25452 21812 25508 23214
rect 25676 23156 25732 23166
rect 25676 23062 25732 23100
rect 26012 23154 26068 23166
rect 26012 23102 26014 23154
rect 26066 23102 26068 23154
rect 25340 21756 25508 21812
rect 25340 21588 25396 21756
rect 25676 21700 25732 21710
rect 25676 21606 25732 21644
rect 25900 21700 25956 21710
rect 25900 21606 25956 21644
rect 25340 21494 25396 21532
rect 25452 21586 25508 21598
rect 25452 21534 25454 21586
rect 25506 21534 25508 21586
rect 25340 20916 25396 20926
rect 25228 20914 25396 20916
rect 25228 20862 25342 20914
rect 25394 20862 25396 20914
rect 25228 20860 25396 20862
rect 25116 20748 25284 20804
rect 24892 20598 24948 20636
rect 25116 20356 25172 20366
rect 24780 20244 24836 20254
rect 24780 20150 24836 20188
rect 24668 19294 24670 19346
rect 24722 19294 24724 19346
rect 24668 19282 24724 19294
rect 24556 19124 24612 19134
rect 24556 19030 24612 19068
rect 23772 17666 23828 18172
rect 23884 18228 23940 18238
rect 23884 18226 24052 18228
rect 23884 18174 23886 18226
rect 23938 18174 24052 18226
rect 23884 18172 24052 18174
rect 23884 18162 23940 18172
rect 23772 17614 23774 17666
rect 23826 17614 23828 17666
rect 23772 17602 23828 17614
rect 23884 18004 23940 18014
rect 23884 17106 23940 17948
rect 23884 17054 23886 17106
rect 23938 17054 23940 17106
rect 23884 17042 23940 17054
rect 23324 16270 23326 16322
rect 23378 16270 23380 16322
rect 23324 16258 23380 16270
rect 23436 16828 23604 16884
rect 23324 16100 23380 16110
rect 23436 16100 23492 16828
rect 23996 16772 24052 18172
rect 24220 17220 24276 18284
rect 24332 18564 24388 18574
rect 24332 17554 24388 18508
rect 24332 17502 24334 17554
rect 24386 17502 24388 17554
rect 24332 17490 24388 17502
rect 24444 18450 24500 18462
rect 24444 18398 24446 18450
rect 24498 18398 24500 18450
rect 23996 16706 24052 16716
rect 24108 17164 24276 17220
rect 24332 17332 24388 17342
rect 24108 16548 24164 17164
rect 24220 16994 24276 17006
rect 24220 16942 24222 16994
rect 24274 16942 24276 16994
rect 24220 16660 24276 16942
rect 24220 16594 24276 16604
rect 23884 16492 24164 16548
rect 23324 16098 23492 16100
rect 23324 16046 23326 16098
rect 23378 16046 23492 16098
rect 23324 16044 23492 16046
rect 23548 16100 23604 16110
rect 23324 16034 23380 16044
rect 23548 15204 23604 16044
rect 23884 16098 23940 16492
rect 23884 16046 23886 16098
rect 23938 16046 23940 16098
rect 23884 16034 23940 16046
rect 24220 16100 24276 16110
rect 24332 16100 24388 17276
rect 24220 16098 24388 16100
rect 24220 16046 24222 16098
rect 24274 16046 24388 16098
rect 24220 16044 24388 16046
rect 24444 16100 24500 18398
rect 25116 18452 25172 20300
rect 25228 20130 25284 20748
rect 25340 20356 25396 20860
rect 25452 20580 25508 21534
rect 25564 21476 25620 21486
rect 25564 21382 25620 21420
rect 26012 21028 26068 23102
rect 26236 23154 26292 23166
rect 26236 23102 26238 23154
rect 26290 23102 26292 23154
rect 26236 22484 26292 23102
rect 26684 23154 26740 23166
rect 26684 23102 26686 23154
rect 26738 23102 26740 23154
rect 26684 22932 26740 23102
rect 26908 23156 26964 23166
rect 26908 23062 26964 23100
rect 27020 22932 27076 22942
rect 26684 22930 27076 22932
rect 26684 22878 27022 22930
rect 27074 22878 27076 22930
rect 26684 22876 27076 22878
rect 27020 22866 27076 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 26236 22418 26292 22428
rect 28252 22484 28308 22494
rect 26124 22260 26180 22270
rect 26124 22258 26292 22260
rect 26124 22206 26126 22258
rect 26178 22206 26292 22258
rect 26124 22204 26292 22206
rect 26124 22194 26180 22204
rect 26236 21698 26292 22204
rect 26236 21646 26238 21698
rect 26290 21646 26292 21698
rect 26236 21634 26292 21646
rect 26348 21812 26404 21822
rect 26348 21586 26404 21756
rect 28252 21700 28308 22428
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 37660 22372 37716 22382
rect 37660 22278 37716 22316
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 28252 21634 28308 21644
rect 26348 21534 26350 21586
rect 26402 21534 26404 21586
rect 26348 21522 26404 21534
rect 27692 21588 27748 21598
rect 28140 21588 28196 21598
rect 27692 21586 28196 21588
rect 27692 21534 27694 21586
rect 27746 21534 28142 21586
rect 28194 21534 28196 21586
rect 27692 21532 28196 21534
rect 27692 21522 27748 21532
rect 28140 21522 28196 21532
rect 28364 21588 28420 21598
rect 37660 21588 37716 21598
rect 28420 21532 28644 21588
rect 28364 21494 28420 21532
rect 26684 21476 26740 21486
rect 26684 21382 26740 21420
rect 26460 21364 26516 21374
rect 26012 20972 26180 21028
rect 25452 20514 25508 20524
rect 25676 20802 25732 20814
rect 25676 20750 25678 20802
rect 25730 20750 25732 20802
rect 25676 20356 25732 20750
rect 25340 20300 26068 20356
rect 26012 20242 26068 20300
rect 26012 20190 26014 20242
rect 26066 20190 26068 20242
rect 26012 20178 26068 20190
rect 26124 20244 26180 20972
rect 26460 20914 26516 21308
rect 26460 20862 26462 20914
rect 26514 20862 26516 20914
rect 26460 20850 26516 20862
rect 26572 21362 26628 21374
rect 26572 21310 26574 21362
rect 26626 21310 26628 21362
rect 26572 20916 26628 21310
rect 27132 21364 27188 21374
rect 27132 21270 27188 21308
rect 27244 21362 27300 21374
rect 27244 21310 27246 21362
rect 27298 21310 27300 21362
rect 26572 20850 26628 20860
rect 26124 20178 26180 20188
rect 26348 20580 26404 20590
rect 25228 20078 25230 20130
rect 25282 20078 25284 20130
rect 25228 20066 25284 20078
rect 25452 19908 25508 19918
rect 25340 19906 25508 19908
rect 25340 19854 25454 19906
rect 25506 19854 25508 19906
rect 25340 19852 25508 19854
rect 25340 18564 25396 19852
rect 25452 19842 25508 19852
rect 26348 19234 26404 20524
rect 27244 20244 27300 21310
rect 27468 21362 27524 21374
rect 27468 21310 27470 21362
rect 27522 21310 27524 21362
rect 27468 20916 27524 21310
rect 27468 20850 27524 20860
rect 28028 21362 28084 21374
rect 28028 21310 28030 21362
rect 28082 21310 28084 21362
rect 27468 20692 27524 20702
rect 27468 20188 27524 20636
rect 28028 20692 28084 21310
rect 28588 20914 28644 21532
rect 37660 21494 37716 21532
rect 40012 21362 40068 21374
rect 40012 21310 40014 21362
rect 40066 21310 40068 21362
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 28588 20862 28590 20914
rect 28642 20862 28644 20914
rect 28588 20850 28644 20862
rect 40012 20916 40068 21310
rect 40012 20850 40068 20860
rect 28028 20626 28084 20636
rect 27244 20178 27300 20188
rect 27356 20132 27524 20188
rect 27244 19460 27300 19470
rect 27356 19460 27412 20132
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 27244 19458 27412 19460
rect 27244 19406 27246 19458
rect 27298 19406 27412 19458
rect 27244 19404 27412 19406
rect 27244 19394 27300 19404
rect 26348 19182 26350 19234
rect 26402 19182 26404 19234
rect 26348 19170 26404 19182
rect 26572 19234 26628 19246
rect 26572 19182 26574 19234
rect 26626 19182 26628 19234
rect 25340 18498 25396 18508
rect 26124 19122 26180 19134
rect 26124 19070 26126 19122
rect 26178 19070 26180 19122
rect 25116 18396 25284 18452
rect 24556 18226 24612 18238
rect 24556 18174 24558 18226
rect 24610 18174 24612 18226
rect 24556 16324 24612 18174
rect 24668 18226 24724 18238
rect 24668 18174 24670 18226
rect 24722 18174 24724 18226
rect 24668 17332 24724 18174
rect 24668 17266 24724 17276
rect 25004 17442 25060 17454
rect 25004 17390 25006 17442
rect 25058 17390 25060 17442
rect 24556 16258 24612 16268
rect 24668 17108 24724 17118
rect 24220 16034 24276 16044
rect 24444 16034 24500 16044
rect 23996 15988 24052 15998
rect 23996 15894 24052 15932
rect 23436 14868 23492 14878
rect 23436 14754 23492 14812
rect 23436 14702 23438 14754
rect 23490 14702 23492 14754
rect 23436 14690 23492 14702
rect 23212 14438 23268 14476
rect 23548 14530 23604 15148
rect 24332 14644 24388 14654
rect 24668 14644 24724 17052
rect 25004 16772 25060 17390
rect 25004 15428 25060 16716
rect 25228 16210 25284 18396
rect 25564 18450 25620 18462
rect 25564 18398 25566 18450
rect 25618 18398 25620 18450
rect 25340 17108 25396 17118
rect 25564 17108 25620 18398
rect 26124 17892 26180 19070
rect 26236 19010 26292 19022
rect 26236 18958 26238 19010
rect 26290 18958 26292 19010
rect 26236 18564 26292 18958
rect 26348 18564 26404 18574
rect 26236 18562 26404 18564
rect 26236 18510 26350 18562
rect 26402 18510 26404 18562
rect 26236 18508 26404 18510
rect 26348 18498 26404 18508
rect 26124 17826 26180 17836
rect 25900 17556 25956 17566
rect 25396 17052 25620 17108
rect 25340 17014 25396 17052
rect 25564 16884 25620 17052
rect 25788 17554 25956 17556
rect 25788 17502 25902 17554
rect 25954 17502 25956 17554
rect 25788 17500 25956 17502
rect 25676 16884 25732 16894
rect 25564 16882 25732 16884
rect 25564 16830 25678 16882
rect 25730 16830 25732 16882
rect 25564 16828 25732 16830
rect 25676 16818 25732 16828
rect 25452 16324 25508 16334
rect 25452 16230 25508 16268
rect 25788 16322 25844 17500
rect 25900 17490 25956 17500
rect 26236 17444 26292 17454
rect 26236 17442 26516 17444
rect 26236 17390 26238 17442
rect 26290 17390 26516 17442
rect 26236 17388 26516 17390
rect 26236 17378 26292 17388
rect 26460 16994 26516 17388
rect 26460 16942 26462 16994
rect 26514 16942 26516 16994
rect 26460 16930 26516 16942
rect 25788 16270 25790 16322
rect 25842 16270 25844 16322
rect 25788 16258 25844 16270
rect 26572 16660 26628 19182
rect 26908 19236 26964 19246
rect 27356 19236 27412 19246
rect 26908 19234 27412 19236
rect 26908 19182 26910 19234
rect 26962 19182 27358 19234
rect 27410 19182 27412 19234
rect 26908 19180 27412 19182
rect 26908 19170 26964 19180
rect 27356 19170 27412 19180
rect 27580 19234 27636 19246
rect 27580 19182 27582 19234
rect 27634 19182 27636 19234
rect 27580 18452 27636 19182
rect 27580 18386 27636 18396
rect 28476 18452 28532 18462
rect 28476 18338 28532 18396
rect 37660 18452 37716 18462
rect 37660 18358 37716 18396
rect 28476 18286 28478 18338
rect 28530 18286 28532 18338
rect 28476 18274 28532 18286
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 37660 17666 37716 17678
rect 37660 17614 37662 17666
rect 37714 17614 37716 17666
rect 25228 16158 25230 16210
rect 25282 16158 25284 16210
rect 25228 16146 25284 16158
rect 25676 15540 25732 15550
rect 25676 15538 26180 15540
rect 25676 15486 25678 15538
rect 25730 15486 26180 15538
rect 25676 15484 26180 15486
rect 25676 15474 25732 15484
rect 25228 15428 25284 15438
rect 25004 15426 25284 15428
rect 25004 15374 25230 15426
rect 25282 15374 25284 15426
rect 25004 15372 25284 15374
rect 25228 15362 25284 15372
rect 26124 15426 26180 15484
rect 26124 15374 26126 15426
rect 26178 15374 26180 15426
rect 26124 15362 26180 15374
rect 25564 15316 25620 15326
rect 25564 15222 25620 15260
rect 25788 15314 25844 15326
rect 25788 15262 25790 15314
rect 25842 15262 25844 15314
rect 25788 15204 25844 15262
rect 26460 15316 26516 15326
rect 26572 15316 26628 16604
rect 28588 16772 28644 16782
rect 28588 15988 28644 16716
rect 37660 16772 37716 17614
rect 40012 17556 40068 17726
rect 40012 17490 40068 17500
rect 37660 16706 37716 16716
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 28588 15922 28644 15932
rect 26460 15314 26628 15316
rect 26460 15262 26462 15314
rect 26514 15262 26628 15314
rect 26460 15260 26628 15262
rect 27580 15316 27636 15326
rect 26460 15250 26516 15260
rect 26236 15202 26292 15214
rect 26236 15150 26238 15202
rect 26290 15150 26292 15202
rect 26236 15148 26292 15150
rect 25788 15138 25844 15148
rect 25900 15092 26292 15148
rect 25900 14756 25956 15092
rect 24388 14588 24724 14644
rect 24332 14550 24388 14588
rect 23548 14478 23550 14530
rect 23602 14478 23604 14530
rect 23548 14466 23604 14478
rect 24668 14530 24724 14588
rect 25452 14700 25956 14756
rect 25452 14642 25508 14700
rect 25452 14590 25454 14642
rect 25506 14590 25508 14642
rect 25452 14578 25508 14590
rect 27580 14644 27636 15260
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 27580 14550 27636 14588
rect 28588 14644 28644 14654
rect 24668 14478 24670 14530
rect 24722 14478 24724 14530
rect 24668 14466 24724 14478
rect 22988 14308 23044 14318
rect 22988 14214 23044 14252
rect 23772 14306 23828 14318
rect 23772 14254 23774 14306
rect 23826 14254 23828 14306
rect 22540 13860 22596 13870
rect 22316 13858 22596 13860
rect 22316 13806 22542 13858
rect 22594 13806 22596 13858
rect 22316 13804 22596 13806
rect 22540 13794 22596 13804
rect 23772 13524 23828 14254
rect 23772 13458 23828 13468
rect 24220 14308 24276 14318
rect 22092 13022 22094 13074
rect 22146 13022 22148 13074
rect 22092 13010 22148 13022
rect 24220 13074 24276 14252
rect 25228 13860 25284 13870
rect 25228 13858 25396 13860
rect 25228 13806 25230 13858
rect 25282 13806 25396 13858
rect 25228 13804 25396 13806
rect 25228 13794 25284 13804
rect 24668 13634 24724 13646
rect 24668 13582 24670 13634
rect 24722 13582 24724 13634
rect 24668 13524 24724 13582
rect 24668 13458 24724 13468
rect 25228 13524 25284 13534
rect 24220 13022 24222 13074
rect 24274 13022 24276 13074
rect 21420 12910 21422 12962
rect 21474 12910 21476 12962
rect 21420 12898 21476 12910
rect 21084 12350 21086 12402
rect 21138 12350 21140 12402
rect 21084 12338 21140 12350
rect 24220 8428 24276 13022
rect 24220 8372 24612 8428
rect 20748 3502 20750 3554
rect 20802 3502 20804 3554
rect 20748 3490 20804 3502
rect 24220 4116 24276 4126
rect 20188 3444 20244 3454
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 800 20244 3388
rect 21756 3444 21812 3454
rect 21756 3330 21812 3388
rect 21756 3278 21758 3330
rect 21810 3278 21812 3330
rect 21756 3266 21812 3278
rect 23548 3444 23604 3454
rect 23548 800 23604 3388
rect 24220 800 24276 4060
rect 24556 3554 24612 8372
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 24892 5236 24948 5246
rect 24892 800 24948 5180
rect 25228 4338 25284 13468
rect 25340 5122 25396 13804
rect 25564 13746 25620 13758
rect 25564 13694 25566 13746
rect 25618 13694 25620 13746
rect 25564 13524 25620 13694
rect 25564 13458 25620 13468
rect 26124 5236 26180 5246
rect 26124 5142 26180 5180
rect 25340 5070 25342 5122
rect 25394 5070 25396 5122
rect 25340 5058 25396 5070
rect 25228 4286 25230 4338
rect 25282 4286 25284 4338
rect 25228 4274 25284 4286
rect 26236 4116 26292 4126
rect 26236 4022 26292 4060
rect 25564 3666 25620 3678
rect 25564 3614 25566 3666
rect 25618 3614 25620 3666
rect 25564 3444 25620 3614
rect 25564 3378 25620 3388
rect 25676 3668 25732 3678
rect 25676 1652 25732 3612
rect 28588 3554 28644 14588
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 29372 3668 29428 3678
rect 29372 3574 29428 3612
rect 28588 3502 28590 3554
rect 28642 3502 28644 3554
rect 28588 3490 28644 3502
rect 25564 1596 25732 1652
rect 25564 800 25620 1596
rect 16128 0 16240 800
rect 18816 0 18928 800
rect 20160 0 20272 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 24864 0 24976 800
rect 25536 0 25648 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 16828 38220 16884 38276
rect 18060 38274 18116 38276
rect 18060 38222 18062 38274
rect 18062 38222 18114 38274
rect 18114 38222 18116 38274
rect 18060 38220 18116 38222
rect 16156 37436 16212 37492
rect 15820 37212 15876 37268
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 1708 36370 1764 36372
rect 1708 36318 1710 36370
rect 1710 36318 1762 36370
rect 1762 36318 1764 36370
rect 1708 36316 1764 36318
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 15708 28700 15764 28756
rect 14588 28588 14644 28644
rect 4172 28252 4228 28308
rect 1932 24498 1988 24500
rect 1932 24446 1934 24498
rect 1934 24446 1986 24498
rect 1986 24446 1988 24498
rect 1932 24444 1988 24446
rect 1932 23548 1988 23604
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 18396 37490 18452 37492
rect 18396 37438 18398 37490
rect 18398 37438 18450 37490
rect 18450 37438 18452 37490
rect 18396 37436 18452 37438
rect 24892 38556 24948 38612
rect 20188 37436 20244 37492
rect 17388 37266 17444 37268
rect 17388 37214 17390 37266
rect 17390 37214 17442 37266
rect 17442 37214 17444 37266
rect 17388 37212 17444 37214
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 14924 28364 14980 28420
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4284 24722 4340 24724
rect 4284 24670 4286 24722
rect 4286 24670 4338 24722
rect 4338 24670 4340 24722
rect 4284 24668 4340 24670
rect 15932 28418 15988 28420
rect 15932 28366 15934 28418
rect 15934 28366 15986 28418
rect 15986 28366 15988 28418
rect 15932 28364 15988 28366
rect 16380 28642 16436 28644
rect 16380 28590 16382 28642
rect 16382 28590 16434 28642
rect 16434 28590 16436 28642
rect 16380 28588 16436 28590
rect 16156 28476 16212 28532
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 17276 28642 17332 28644
rect 17276 28590 17278 28642
rect 17278 28590 17330 28642
rect 17330 28590 17332 28642
rect 17276 28588 17332 28590
rect 19516 28530 19572 28532
rect 19516 28478 19518 28530
rect 19518 28478 19570 28530
rect 19570 28478 19572 28530
rect 19516 28476 19572 28478
rect 16940 28364 16996 28420
rect 16940 27074 16996 27076
rect 16940 27022 16942 27074
rect 16942 27022 16994 27074
rect 16994 27022 16996 27074
rect 16940 27020 16996 27022
rect 15148 25228 15204 25284
rect 10780 24668 10836 24724
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4284 23938 4340 23940
rect 4284 23886 4286 23938
rect 4286 23886 4338 23938
rect 4338 23886 4340 23938
rect 4284 23884 4340 23886
rect 12796 23996 12852 24052
rect 11004 23884 11060 23940
rect 10892 23772 10948 23828
rect 12796 23826 12852 23828
rect 12796 23774 12798 23826
rect 12798 23774 12850 23826
rect 12850 23774 12852 23826
rect 12796 23772 12852 23774
rect 13020 23772 13076 23828
rect 13132 23660 13188 23716
rect 13580 23884 13636 23940
rect 13468 23826 13524 23828
rect 13468 23774 13470 23826
rect 13470 23774 13522 23826
rect 13522 23774 13524 23826
rect 13468 23772 13524 23774
rect 13244 23324 13300 23380
rect 14028 23996 14084 24052
rect 15932 24556 15988 24612
rect 16604 26796 16660 26852
rect 17500 26796 17556 26852
rect 17612 27020 17668 27076
rect 18620 26796 18676 26852
rect 16156 23996 16212 24052
rect 13692 23548 13748 23604
rect 14140 23714 14196 23716
rect 14140 23662 14142 23714
rect 14142 23662 14194 23714
rect 14194 23662 14196 23714
rect 14140 23660 14196 23662
rect 14364 23660 14420 23716
rect 14588 23378 14644 23380
rect 14588 23326 14590 23378
rect 14590 23326 14642 23378
rect 14642 23326 14644 23378
rect 14588 23324 14644 23326
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 15148 23548 15204 23604
rect 14812 23378 14868 23380
rect 14812 23326 14814 23378
rect 14814 23326 14866 23378
rect 14866 23326 14868 23378
rect 14812 23324 14868 23326
rect 15820 23378 15876 23380
rect 15820 23326 15822 23378
rect 15822 23326 15874 23378
rect 15874 23326 15876 23378
rect 15820 23324 15876 23326
rect 17052 23660 17108 23716
rect 16380 23154 16436 23156
rect 16380 23102 16382 23154
rect 16382 23102 16434 23154
rect 16434 23102 16436 23154
rect 16380 23100 16436 23102
rect 14700 22428 14756 22484
rect 17052 22764 17108 22820
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 14476 20748 14532 20804
rect 4172 19964 4228 20020
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 12908 19906 12964 19908
rect 12908 19854 12910 19906
rect 12910 19854 12962 19906
rect 12962 19854 12964 19906
rect 12908 19852 12964 19854
rect 11788 18396 11844 18452
rect 12796 18396 12852 18452
rect 12348 18338 12404 18340
rect 12348 18286 12350 18338
rect 12350 18286 12402 18338
rect 12402 18286 12404 18338
rect 12348 18284 12404 18286
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 1932 17778 1988 17780
rect 1932 17726 1934 17778
rect 1934 17726 1986 17778
rect 1986 17726 1988 17778
rect 1932 17724 1988 17726
rect 4284 17666 4340 17668
rect 4284 17614 4286 17666
rect 4286 17614 4338 17666
rect 4338 17614 4340 17666
rect 4284 17612 4340 17614
rect 9996 17612 10052 17668
rect 1932 16828 1988 16884
rect 4284 16882 4340 16884
rect 4284 16830 4286 16882
rect 4286 16830 4338 16882
rect 4338 16830 4340 16882
rect 4284 16828 4340 16830
rect 15036 20802 15092 20804
rect 15036 20750 15038 20802
rect 15038 20750 15090 20802
rect 15090 20750 15092 20802
rect 15036 20748 15092 20750
rect 16492 20802 16548 20804
rect 16492 20750 16494 20802
rect 16494 20750 16546 20802
rect 16546 20750 16548 20802
rect 16492 20748 16548 20750
rect 15036 20076 15092 20132
rect 15260 19852 15316 19908
rect 15708 19852 15764 19908
rect 15484 19404 15540 19460
rect 14812 18732 14868 18788
rect 12796 17666 12852 17668
rect 12796 17614 12798 17666
rect 12798 17614 12850 17666
rect 12850 17614 12852 17666
rect 12796 17612 12852 17614
rect 13580 17666 13636 17668
rect 13580 17614 13582 17666
rect 13582 17614 13634 17666
rect 13634 17614 13636 17666
rect 13580 17612 13636 17614
rect 14252 17500 14308 17556
rect 14364 17612 14420 17668
rect 12124 17388 12180 17444
rect 14140 17442 14196 17444
rect 14140 17390 14142 17442
rect 14142 17390 14194 17442
rect 14194 17390 14196 17442
rect 14140 17388 14196 17390
rect 9996 16716 10052 16772
rect 12796 16828 12852 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4284 16098 4340 16100
rect 4284 16046 4286 16098
rect 4286 16046 4338 16098
rect 4338 16046 4340 16098
rect 4284 16044 4340 16046
rect 11228 16044 11284 16100
rect 1932 15484 1988 15540
rect 13692 16044 13748 16100
rect 13804 15986 13860 15988
rect 13804 15934 13806 15986
rect 13806 15934 13858 15986
rect 13858 15934 13860 15986
rect 13804 15932 13860 15934
rect 13356 15820 13412 15876
rect 14924 18338 14980 18340
rect 14924 18286 14926 18338
rect 14926 18286 14978 18338
rect 14978 18286 14980 18338
rect 14924 18284 14980 18286
rect 14924 17612 14980 17668
rect 17500 24610 17556 24612
rect 17500 24558 17502 24610
rect 17502 24558 17554 24610
rect 17554 24558 17556 24610
rect 17500 24556 17556 24558
rect 17612 23660 17668 23716
rect 17836 23100 17892 23156
rect 17388 22930 17444 22932
rect 17388 22878 17390 22930
rect 17390 22878 17442 22930
rect 17442 22878 17444 22930
rect 17388 22876 17444 22878
rect 17948 22764 18004 22820
rect 19628 28364 19684 28420
rect 20300 28476 20356 28532
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19292 27746 19348 27748
rect 19292 27694 19294 27746
rect 19294 27694 19346 27746
rect 19346 27694 19348 27746
rect 19292 27692 19348 27694
rect 20524 28530 20580 28532
rect 20524 28478 20526 28530
rect 20526 28478 20578 28530
rect 20578 28478 20580 28530
rect 20524 28476 20580 28478
rect 21420 37490 21476 37492
rect 21420 37438 21422 37490
rect 21422 37438 21474 37490
rect 21474 37438 21476 37490
rect 21420 37436 21476 37438
rect 22204 28588 22260 28644
rect 20636 27692 20692 27748
rect 22204 27692 22260 27748
rect 20748 26962 20804 26964
rect 20748 26910 20750 26962
rect 20750 26910 20802 26962
rect 20802 26910 20804 26962
rect 20748 26908 20804 26910
rect 21868 26908 21924 26964
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 18844 24892 18900 24948
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19740 24946 19796 24948
rect 19740 24894 19742 24946
rect 19742 24894 19794 24946
rect 19794 24894 19796 24946
rect 19740 24892 19796 24894
rect 19292 24722 19348 24724
rect 19292 24670 19294 24722
rect 19294 24670 19346 24722
rect 19346 24670 19348 24722
rect 19292 24668 19348 24670
rect 20300 24668 20356 24724
rect 19516 24108 19572 24164
rect 19852 24220 19908 24276
rect 18844 23714 18900 23716
rect 18844 23662 18846 23714
rect 18846 23662 18898 23714
rect 18898 23662 18900 23714
rect 18844 23660 18900 23662
rect 18284 23154 18340 23156
rect 18284 23102 18286 23154
rect 18286 23102 18338 23154
rect 18338 23102 18340 23154
rect 18284 23100 18340 23102
rect 18060 21980 18116 22036
rect 17388 20802 17444 20804
rect 17388 20750 17390 20802
rect 17390 20750 17442 20802
rect 17442 20750 17444 20802
rect 17388 20748 17444 20750
rect 18060 21308 18116 21364
rect 17724 20748 17780 20804
rect 17724 20524 17780 20580
rect 17388 20130 17444 20132
rect 17388 20078 17390 20130
rect 17390 20078 17442 20130
rect 17442 20078 17444 20130
rect 17388 20076 17444 20078
rect 17612 20076 17668 20132
rect 17052 18732 17108 18788
rect 16716 18284 16772 18340
rect 14700 17388 14756 17444
rect 14700 16604 14756 16660
rect 15484 17500 15540 17556
rect 15484 17276 15540 17332
rect 16492 17500 16548 17556
rect 15708 17052 15764 17108
rect 17612 19516 17668 19572
rect 17948 20076 18004 20132
rect 17948 19516 18004 19572
rect 17724 19122 17780 19124
rect 17724 19070 17726 19122
rect 17726 19070 17778 19122
rect 17778 19070 17780 19122
rect 17724 19068 17780 19070
rect 18396 21084 18452 21140
rect 18620 22540 18676 22596
rect 18620 21980 18676 22036
rect 18844 22146 18900 22148
rect 18844 22094 18846 22146
rect 18846 22094 18898 22146
rect 18898 22094 18900 22146
rect 18844 22092 18900 22094
rect 18508 20578 18564 20580
rect 18508 20526 18510 20578
rect 18510 20526 18562 20578
rect 18562 20526 18564 20578
rect 18508 20524 18564 20526
rect 18620 20300 18676 20356
rect 18844 21532 18900 21588
rect 19852 23884 19908 23940
rect 19516 23660 19572 23716
rect 19068 22876 19124 22932
rect 20412 23884 20468 23940
rect 20300 23772 20356 23828
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20076 23154 20132 23156
rect 20076 23102 20078 23154
rect 20078 23102 20130 23154
rect 20130 23102 20132 23154
rect 20076 23100 20132 23102
rect 20076 22876 20132 22932
rect 19516 22258 19572 22260
rect 19516 22206 19518 22258
rect 19518 22206 19570 22258
rect 19570 22206 19572 22258
rect 19516 22204 19572 22206
rect 19404 22092 19460 22148
rect 20524 23714 20580 23716
rect 20524 23662 20526 23714
rect 20526 23662 20578 23714
rect 20578 23662 20580 23714
rect 20524 23660 20580 23662
rect 20412 22652 20468 22708
rect 26124 38556 26180 38612
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 26236 38220 26292 38276
rect 29372 38274 29428 38276
rect 29372 38222 29374 38274
rect 29374 38222 29426 38274
rect 29426 38222 29428 38274
rect 29372 38220 29428 38222
rect 22764 27746 22820 27748
rect 22764 27694 22766 27746
rect 22766 27694 22818 27746
rect 22818 27694 22820 27746
rect 22764 27692 22820 27694
rect 24220 27132 24276 27188
rect 21420 24220 21476 24276
rect 21980 25340 22036 25396
rect 22092 25228 22148 25284
rect 21308 23938 21364 23940
rect 21308 23886 21310 23938
rect 21310 23886 21362 23938
rect 21362 23886 21364 23938
rect 21308 23884 21364 23886
rect 21868 23996 21924 24052
rect 21420 23772 21476 23828
rect 21196 22652 21252 22708
rect 21420 22764 21476 22820
rect 22204 23826 22260 23828
rect 22204 23774 22206 23826
rect 22206 23774 22258 23826
rect 22258 23774 22260 23826
rect 22204 23772 22260 23774
rect 22092 23436 22148 23492
rect 25004 27186 25060 27188
rect 25004 27134 25006 27186
rect 25006 27134 25058 27186
rect 25058 27134 25060 27186
rect 25004 27132 25060 27134
rect 25452 27746 25508 27748
rect 25452 27694 25454 27746
rect 25454 27694 25506 27746
rect 25506 27694 25508 27746
rect 25452 27692 25508 27694
rect 24780 26908 24836 26964
rect 22988 26290 23044 26292
rect 22988 26238 22990 26290
rect 22990 26238 23042 26290
rect 23042 26238 23044 26290
rect 22988 26236 23044 26238
rect 23100 25788 23156 25844
rect 23100 25340 23156 25396
rect 19628 21980 19684 22036
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 18508 20018 18564 20020
rect 18508 19966 18510 20018
rect 18510 19966 18562 20018
rect 18562 19966 18564 20018
rect 18508 19964 18564 19966
rect 18172 19852 18228 19908
rect 19068 21084 19124 21140
rect 18172 19292 18228 19348
rect 18620 19404 18676 19460
rect 18732 19234 18788 19236
rect 18732 19182 18734 19234
rect 18734 19182 18786 19234
rect 18786 19182 18788 19234
rect 18732 19180 18788 19182
rect 17276 18060 17332 18116
rect 17164 17554 17220 17556
rect 17164 17502 17166 17554
rect 17166 17502 17218 17554
rect 17218 17502 17220 17554
rect 17164 17500 17220 17502
rect 16716 17052 16772 17108
rect 16268 16994 16324 16996
rect 16268 16942 16270 16994
rect 16270 16942 16322 16994
rect 16322 16942 16324 16994
rect 16268 16940 16324 16942
rect 18060 18508 18116 18564
rect 18060 18172 18116 18228
rect 17724 17500 17780 17556
rect 17500 17388 17556 17444
rect 17724 16940 17780 16996
rect 18172 17724 18228 17780
rect 18396 18956 18452 19012
rect 18508 18450 18564 18452
rect 18508 18398 18510 18450
rect 18510 18398 18562 18450
rect 18562 18398 18564 18450
rect 18508 18396 18564 18398
rect 18956 20524 19012 20580
rect 18844 18226 18900 18228
rect 18844 18174 18846 18226
rect 18846 18174 18898 18226
rect 18898 18174 18900 18226
rect 18844 18172 18900 18174
rect 19180 21026 19236 21028
rect 19180 20974 19182 21026
rect 19182 20974 19234 21026
rect 19234 20974 19236 21026
rect 19180 20972 19236 20974
rect 19292 20802 19348 20804
rect 19292 20750 19294 20802
rect 19294 20750 19346 20802
rect 19346 20750 19348 20802
rect 19292 20748 19348 20750
rect 19292 20300 19348 20356
rect 19180 20188 19236 20244
rect 19068 18284 19124 18340
rect 19516 21362 19572 21364
rect 19516 21310 19518 21362
rect 19518 21310 19570 21362
rect 19570 21310 19572 21362
rect 19516 21308 19572 21310
rect 19404 19234 19460 19236
rect 19404 19182 19406 19234
rect 19406 19182 19458 19234
rect 19458 19182 19460 19234
rect 19404 19180 19460 19182
rect 20076 21084 20132 21140
rect 20188 20914 20244 20916
rect 20188 20862 20190 20914
rect 20190 20862 20242 20914
rect 20242 20862 20244 20914
rect 20188 20860 20244 20862
rect 19852 20802 19908 20804
rect 19852 20750 19854 20802
rect 19854 20750 19906 20802
rect 19906 20750 19908 20802
rect 19852 20748 19908 20750
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19740 20018 19796 20020
rect 19740 19966 19742 20018
rect 19742 19966 19794 20018
rect 19794 19966 19796 20018
rect 19740 19964 19796 19966
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 18396 17724 18452 17780
rect 18620 17554 18676 17556
rect 18620 17502 18622 17554
rect 18622 17502 18674 17554
rect 18674 17502 18676 17554
rect 18620 17500 18676 17502
rect 15148 16716 15204 16772
rect 15260 15986 15316 15988
rect 15260 15934 15262 15986
rect 15262 15934 15314 15986
rect 15314 15934 15316 15986
rect 15260 15932 15316 15934
rect 15596 15932 15652 15988
rect 14588 15874 14644 15876
rect 14588 15822 14590 15874
rect 14590 15822 14642 15874
rect 14642 15822 14644 15874
rect 14588 15820 14644 15822
rect 13580 15036 13636 15092
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 14588 15036 14644 15092
rect 17836 16770 17892 16772
rect 17836 16718 17838 16770
rect 17838 16718 17890 16770
rect 17890 16718 17892 16770
rect 17836 16716 17892 16718
rect 17164 16098 17220 16100
rect 17164 16046 17166 16098
rect 17166 16046 17218 16098
rect 17218 16046 17220 16098
rect 17164 16044 17220 16046
rect 16156 15932 16212 15988
rect 16828 15986 16884 15988
rect 16828 15934 16830 15986
rect 16830 15934 16882 15986
rect 16882 15934 16884 15986
rect 16828 15932 16884 15934
rect 18172 15820 18228 15876
rect 16156 15036 16212 15092
rect 15932 14306 15988 14308
rect 15932 14254 15934 14306
rect 15934 14254 15986 14306
rect 15986 14254 15988 14306
rect 15932 14252 15988 14254
rect 15708 13580 15764 13636
rect 16492 13634 16548 13636
rect 16492 13582 16494 13634
rect 16494 13582 16546 13634
rect 16546 13582 16548 13634
rect 16492 13580 16548 13582
rect 14364 13468 14420 13524
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 17388 14252 17444 14308
rect 17948 13804 18004 13860
rect 17612 13746 17668 13748
rect 17612 13694 17614 13746
rect 17614 13694 17666 13746
rect 17666 13694 17668 13746
rect 17612 13692 17668 13694
rect 18396 16940 18452 16996
rect 18508 17052 18564 17108
rect 18732 16604 18788 16660
rect 18956 17836 19012 17892
rect 19068 17500 19124 17556
rect 19068 16716 19124 16772
rect 19292 16210 19348 16212
rect 19292 16158 19294 16210
rect 19294 16158 19346 16210
rect 19346 16158 19348 16210
rect 19292 16156 19348 16158
rect 18956 16098 19012 16100
rect 18956 16046 18958 16098
rect 18958 16046 19010 16098
rect 19010 16046 19012 16098
rect 18956 16044 19012 16046
rect 19516 18284 19572 18340
rect 19516 18060 19572 18116
rect 19740 18396 19796 18452
rect 19516 17724 19572 17780
rect 19516 17276 19572 17332
rect 19516 16604 19572 16660
rect 18956 15874 19012 15876
rect 18956 15822 18958 15874
rect 18958 15822 19010 15874
rect 19010 15822 19012 15874
rect 18956 15820 19012 15822
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19628 15820 19684 15876
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20300 19180 20356 19236
rect 20524 22204 20580 22260
rect 21308 22258 21364 22260
rect 21308 22206 21310 22258
rect 21310 22206 21362 22258
rect 21362 22206 21364 22258
rect 21308 22204 21364 22206
rect 21756 22540 21812 22596
rect 21644 22428 21700 22484
rect 21420 21868 21476 21924
rect 20972 20860 21028 20916
rect 21756 21868 21812 21924
rect 21532 20748 21588 20804
rect 21868 20972 21924 21028
rect 21756 20188 21812 20244
rect 20860 19404 20916 19460
rect 20524 19292 20580 19348
rect 21868 19180 21924 19236
rect 20412 18508 20468 18564
rect 21196 18508 21252 18564
rect 21756 18450 21812 18452
rect 21756 18398 21758 18450
rect 21758 18398 21810 18450
rect 21810 18398 21812 18450
rect 21756 18396 21812 18398
rect 20748 17948 20804 18004
rect 20412 17836 20468 17892
rect 20300 15260 20356 15316
rect 16716 13074 16772 13076
rect 16716 13022 16718 13074
rect 16718 13022 16770 13074
rect 16770 13022 16772 13074
rect 16716 13020 16772 13022
rect 16940 13580 16996 13636
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 17500 13522 17556 13524
rect 17500 13470 17502 13522
rect 17502 13470 17554 13522
rect 17554 13470 17556 13522
rect 17500 13468 17556 13470
rect 17724 13020 17780 13076
rect 18508 12850 18564 12852
rect 18508 12798 18510 12850
rect 18510 12798 18562 12850
rect 18562 12798 18564 12850
rect 18508 12796 18564 12798
rect 19516 14642 19572 14644
rect 19516 14590 19518 14642
rect 19518 14590 19570 14642
rect 19570 14590 19572 14642
rect 19516 14588 19572 14590
rect 20300 14476 20356 14532
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19180 13804 19236 13860
rect 19516 13858 19572 13860
rect 19516 13806 19518 13858
rect 19518 13806 19570 13858
rect 19570 13806 19572 13858
rect 19516 13804 19572 13806
rect 22428 23100 22484 23156
rect 22204 18620 22260 18676
rect 22988 22652 23044 22708
rect 22876 21586 22932 21588
rect 22876 21534 22878 21586
rect 22878 21534 22930 21586
rect 22930 21534 22932 21586
rect 22876 21532 22932 21534
rect 22540 20972 22596 21028
rect 21980 18396 22036 18452
rect 21980 17388 22036 17444
rect 20524 16156 20580 16212
rect 21196 16156 21252 16212
rect 22764 20188 22820 20244
rect 23212 23996 23268 24052
rect 23996 26290 24052 26292
rect 23996 26238 23998 26290
rect 23998 26238 24050 26290
rect 24050 26238 24052 26290
rect 23996 26236 24052 26238
rect 24668 26236 24724 26292
rect 23884 26124 23940 26180
rect 23884 25788 23940 25844
rect 23100 21644 23156 21700
rect 23436 23772 23492 23828
rect 23324 20914 23380 20916
rect 23324 20862 23326 20914
rect 23326 20862 23378 20914
rect 23378 20862 23380 20914
rect 23324 20860 23380 20862
rect 22988 20076 23044 20132
rect 25116 26124 25172 26180
rect 23884 21868 23940 21924
rect 23772 21810 23828 21812
rect 23772 21758 23774 21810
rect 23774 21758 23826 21810
rect 23826 21758 23828 21810
rect 23772 21756 23828 21758
rect 23548 21308 23604 21364
rect 24332 20972 24388 21028
rect 23660 20802 23716 20804
rect 23660 20750 23662 20802
rect 23662 20750 23714 20802
rect 23714 20750 23716 20802
rect 23660 20748 23716 20750
rect 23548 20300 23604 20356
rect 23660 19964 23716 20020
rect 22988 18562 23044 18564
rect 22988 18510 22990 18562
rect 22990 18510 23042 18562
rect 23042 18510 23044 18562
rect 22988 18508 23044 18510
rect 23436 19292 23492 19348
rect 23100 17948 23156 18004
rect 22876 16044 22932 16100
rect 20636 15874 20692 15876
rect 20636 15822 20638 15874
rect 20638 15822 20690 15874
rect 20690 15822 20692 15874
rect 20636 15820 20692 15822
rect 21644 15820 21700 15876
rect 22428 15820 22484 15876
rect 21196 15314 21252 15316
rect 21196 15262 21198 15314
rect 21198 15262 21250 15314
rect 21250 15262 21252 15314
rect 21196 15260 21252 15262
rect 22428 15314 22484 15316
rect 22428 15262 22430 15314
rect 22430 15262 22482 15314
rect 22482 15262 22484 15314
rect 22428 15260 22484 15262
rect 22204 14812 22260 14868
rect 21644 14700 21700 14756
rect 21308 14140 21364 14196
rect 21868 14588 21924 14644
rect 20412 13746 20468 13748
rect 20412 13694 20414 13746
rect 20414 13694 20466 13746
rect 20466 13694 20468 13746
rect 20412 13692 20468 13694
rect 20636 13804 20692 13860
rect 20076 12796 20132 12852
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 18844 4060 18900 4116
rect 16156 3388 16212 3444
rect 18508 3442 18564 3444
rect 18508 3390 18510 3442
rect 18510 3390 18562 3442
rect 18562 3390 18564 3442
rect 18508 3388 18564 3390
rect 20076 4114 20132 4116
rect 20076 4062 20078 4114
rect 20078 4062 20130 4114
rect 20130 4062 20132 4114
rect 20076 4060 20132 4062
rect 22092 14140 22148 14196
rect 22652 14754 22708 14756
rect 22652 14702 22654 14754
rect 22654 14702 22706 14754
rect 22706 14702 22708 14754
rect 22652 14700 22708 14702
rect 22540 14530 22596 14532
rect 22540 14478 22542 14530
rect 22542 14478 22594 14530
rect 22594 14478 22596 14530
rect 22540 14476 22596 14478
rect 23660 19068 23716 19124
rect 23548 18396 23604 18452
rect 24108 18450 24164 18452
rect 24108 18398 24110 18450
rect 24110 18398 24162 18450
rect 24162 18398 24164 18450
rect 24108 18396 24164 18398
rect 26124 26962 26180 26964
rect 26124 26910 26126 26962
rect 26126 26910 26178 26962
rect 26178 26910 26180 26962
rect 26124 26908 26180 26910
rect 26236 26796 26292 26852
rect 25564 26402 25620 26404
rect 25564 26350 25566 26402
rect 25566 26350 25618 26402
rect 25618 26350 25620 26402
rect 25564 26348 25620 26350
rect 28252 26796 28308 26852
rect 26460 26514 26516 26516
rect 26460 26462 26462 26514
rect 26462 26462 26514 26514
rect 26514 26462 26516 26514
rect 26460 26460 26516 26462
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 28588 26460 28644 26516
rect 26236 26348 26292 26404
rect 25676 26290 25732 26292
rect 25676 26238 25678 26290
rect 25678 26238 25730 26290
rect 25730 26238 25732 26290
rect 25676 26236 25732 26238
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 27020 23996 27076 24052
rect 25340 23436 25396 23492
rect 28588 24050 28644 24052
rect 28588 23998 28590 24050
rect 28590 23998 28642 24050
rect 28642 23998 28644 24050
rect 28588 23996 28644 23998
rect 37660 23938 37716 23940
rect 37660 23886 37662 23938
rect 37662 23886 37714 23938
rect 37714 23886 37716 23938
rect 37660 23884 37716 23886
rect 40012 23548 40068 23604
rect 25340 22540 25396 22596
rect 25116 21868 25172 21924
rect 24892 21532 24948 21588
rect 24556 21084 24612 21140
rect 24556 20524 24612 20580
rect 24556 20300 24612 20356
rect 24444 20130 24500 20132
rect 24444 20078 24446 20130
rect 24446 20078 24498 20130
rect 24498 20078 24500 20130
rect 24444 20076 24500 20078
rect 25676 23154 25732 23156
rect 25676 23102 25678 23154
rect 25678 23102 25730 23154
rect 25730 23102 25732 23154
rect 25676 23100 25732 23102
rect 25676 21698 25732 21700
rect 25676 21646 25678 21698
rect 25678 21646 25730 21698
rect 25730 21646 25732 21698
rect 25676 21644 25732 21646
rect 25900 21698 25956 21700
rect 25900 21646 25902 21698
rect 25902 21646 25954 21698
rect 25954 21646 25956 21698
rect 25900 21644 25956 21646
rect 25340 21586 25396 21588
rect 25340 21534 25342 21586
rect 25342 21534 25394 21586
rect 25394 21534 25396 21586
rect 25340 21532 25396 21534
rect 24892 20690 24948 20692
rect 24892 20638 24894 20690
rect 24894 20638 24946 20690
rect 24946 20638 24948 20690
rect 24892 20636 24948 20638
rect 25116 20300 25172 20356
rect 24780 20242 24836 20244
rect 24780 20190 24782 20242
rect 24782 20190 24834 20242
rect 24834 20190 24836 20242
rect 24780 20188 24836 20190
rect 24556 19122 24612 19124
rect 24556 19070 24558 19122
rect 24558 19070 24610 19122
rect 24610 19070 24612 19122
rect 24556 19068 24612 19070
rect 24220 18284 24276 18340
rect 23772 18172 23828 18228
rect 23884 17948 23940 18004
rect 24332 18508 24388 18564
rect 23996 16716 24052 16772
rect 24332 17276 24388 17332
rect 24220 16604 24276 16660
rect 23548 16044 23604 16100
rect 25564 21474 25620 21476
rect 25564 21422 25566 21474
rect 25566 21422 25618 21474
rect 25618 21422 25620 21474
rect 25564 21420 25620 21422
rect 26908 23154 26964 23156
rect 26908 23102 26910 23154
rect 26910 23102 26962 23154
rect 26962 23102 26964 23154
rect 26908 23100 26964 23102
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 26236 22428 26292 22484
rect 28252 22482 28308 22484
rect 28252 22430 28254 22482
rect 28254 22430 28306 22482
rect 28306 22430 28308 22482
rect 28252 22428 28308 22430
rect 26348 21756 26404 21812
rect 37660 22370 37716 22372
rect 37660 22318 37662 22370
rect 37662 22318 37714 22370
rect 37714 22318 37716 22370
rect 37660 22316 37716 22318
rect 40012 22204 40068 22260
rect 28252 21644 28308 21700
rect 28364 21586 28420 21588
rect 28364 21534 28366 21586
rect 28366 21534 28418 21586
rect 28418 21534 28420 21586
rect 28364 21532 28420 21534
rect 26684 21474 26740 21476
rect 26684 21422 26686 21474
rect 26686 21422 26738 21474
rect 26738 21422 26740 21474
rect 26684 21420 26740 21422
rect 26460 21308 26516 21364
rect 25452 20524 25508 20580
rect 27132 21362 27188 21364
rect 27132 21310 27134 21362
rect 27134 21310 27186 21362
rect 27186 21310 27188 21362
rect 27132 21308 27188 21310
rect 26572 20860 26628 20916
rect 26124 20188 26180 20244
rect 26348 20524 26404 20580
rect 27468 20860 27524 20916
rect 27244 20188 27300 20244
rect 27468 20636 27524 20692
rect 37660 21586 37716 21588
rect 37660 21534 37662 21586
rect 37662 21534 37714 21586
rect 37714 21534 37716 21586
rect 37660 21532 37716 21534
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 40012 20860 40068 20916
rect 28028 20636 28084 20692
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 25340 18508 25396 18564
rect 24668 17276 24724 17332
rect 24556 16268 24612 16324
rect 24668 17106 24724 17108
rect 24668 17054 24670 17106
rect 24670 17054 24722 17106
rect 24722 17054 24724 17106
rect 24668 17052 24724 17054
rect 24444 16044 24500 16100
rect 23996 15986 24052 15988
rect 23996 15934 23998 15986
rect 23998 15934 24050 15986
rect 24050 15934 24052 15986
rect 23996 15932 24052 15934
rect 23548 15148 23604 15204
rect 23436 14812 23492 14868
rect 23212 14530 23268 14532
rect 23212 14478 23214 14530
rect 23214 14478 23266 14530
rect 23266 14478 23268 14530
rect 23212 14476 23268 14478
rect 25004 16716 25060 16772
rect 26124 17836 26180 17892
rect 25340 17106 25396 17108
rect 25340 17054 25342 17106
rect 25342 17054 25394 17106
rect 25394 17054 25396 17106
rect 25340 17052 25396 17054
rect 25452 16322 25508 16324
rect 25452 16270 25454 16322
rect 25454 16270 25506 16322
rect 25506 16270 25508 16322
rect 25452 16268 25508 16270
rect 27580 18396 27636 18452
rect 28476 18396 28532 18452
rect 37660 18450 37716 18452
rect 37660 18398 37662 18450
rect 37662 18398 37714 18450
rect 37714 18398 37716 18450
rect 37660 18396 37716 18398
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 26572 16604 26628 16660
rect 25564 15314 25620 15316
rect 25564 15262 25566 15314
rect 25566 15262 25618 15314
rect 25618 15262 25620 15314
rect 25564 15260 25620 15262
rect 28588 16770 28644 16772
rect 28588 16718 28590 16770
rect 28590 16718 28642 16770
rect 28642 16718 28644 16770
rect 28588 16716 28644 16718
rect 40012 17500 40068 17556
rect 37660 16716 37716 16772
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 28588 15932 28644 15988
rect 27580 15260 27636 15316
rect 25788 15148 25844 15204
rect 24332 14642 24388 14644
rect 24332 14590 24334 14642
rect 24334 14590 24386 14642
rect 24386 14590 24388 14642
rect 24332 14588 24388 14590
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 27580 14642 27636 14644
rect 27580 14590 27582 14642
rect 27582 14590 27634 14642
rect 27634 14590 27636 14642
rect 27580 14588 27636 14590
rect 28588 14588 28644 14644
rect 22988 14306 23044 14308
rect 22988 14254 22990 14306
rect 22990 14254 23042 14306
rect 23042 14254 23044 14306
rect 22988 14252 23044 14254
rect 23772 13468 23828 13524
rect 24220 14252 24276 14308
rect 24668 13468 24724 13524
rect 25228 13468 25284 13524
rect 24220 4060 24276 4116
rect 20188 3388 20244 3444
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 21756 3388 21812 3444
rect 23548 3388 23604 3444
rect 24892 5180 24948 5236
rect 25564 13468 25620 13524
rect 26124 5234 26180 5236
rect 26124 5182 26126 5234
rect 26126 5182 26178 5234
rect 26178 5182 26180 5234
rect 26124 5180 26180 5182
rect 26236 4114 26292 4116
rect 26236 4062 26238 4114
rect 26238 4062 26290 4114
rect 26290 4062 26292 4114
rect 26236 4060 26292 4062
rect 25564 3388 25620 3444
rect 25676 3612 25732 3668
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 29372 3666 29428 3668
rect 29372 3614 29374 3666
rect 29374 3614 29426 3666
rect 29426 3614 29428 3666
rect 29372 3612 29428 3614
<< metal3 >>
rect 24882 38556 24892 38612
rect 24948 38556 26124 38612
rect 26180 38556 26190 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 16818 38220 16828 38276
rect 16884 38220 18060 38276
rect 18116 38220 18126 38276
rect 26226 38220 26236 38276
rect 26292 38220 29372 38276
rect 29428 38220 29438 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 16146 37436 16156 37492
rect 16212 37436 18396 37492
rect 18452 37436 18462 37492
rect 20178 37436 20188 37492
rect 20244 37436 21420 37492
rect 21476 37436 21486 37492
rect 15810 37212 15820 37268
rect 15876 37212 17388 37268
rect 17444 37212 17454 37268
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 0 36372 800 36400
rect 0 36316 1708 36372
rect 1764 36316 1774 36372
rect 0 36288 800 36316
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 15698 28700 15708 28756
rect 15764 28700 17332 28756
rect 17276 28644 17332 28700
rect 14578 28588 14588 28644
rect 14644 28588 16380 28644
rect 16436 28588 16446 28644
rect 17266 28588 17276 28644
rect 17332 28588 22204 28644
rect 22260 28588 22270 28644
rect 16146 28476 16156 28532
rect 16212 28476 16324 28532
rect 19506 28476 19516 28532
rect 19572 28476 20300 28532
rect 20356 28476 20366 28532
rect 20514 28476 20524 28532
rect 20580 28476 20590 28532
rect 16268 28420 16324 28476
rect 20524 28420 20580 28476
rect 14914 28364 14924 28420
rect 14980 28364 15932 28420
rect 15988 28364 15998 28420
rect 16268 28364 16940 28420
rect 16996 28364 19628 28420
rect 19684 28364 20580 28420
rect 0 28308 800 28336
rect 0 28252 4172 28308
rect 4228 28252 4238 28308
rect 0 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 19282 27692 19292 27748
rect 19348 27692 20636 27748
rect 20692 27692 20702 27748
rect 22194 27692 22204 27748
rect 22260 27692 22764 27748
rect 22820 27692 25452 27748
rect 25508 27692 25518 27748
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 24210 27132 24220 27188
rect 24276 27132 25004 27188
rect 25060 27132 25070 27188
rect 16930 27020 16940 27076
rect 16996 27020 17612 27076
rect 17668 27020 17678 27076
rect 20132 26908 20748 26964
rect 20804 26908 21868 26964
rect 21924 26908 21934 26964
rect 24770 26908 24780 26964
rect 24836 26908 26124 26964
rect 26180 26908 26190 26964
rect 20132 26852 20188 26908
rect 16594 26796 16604 26852
rect 16660 26796 17500 26852
rect 17556 26796 18620 26852
rect 18676 26796 20188 26852
rect 26226 26796 26236 26852
rect 26292 26796 28252 26852
rect 28308 26796 28318 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 26450 26460 26460 26516
rect 26516 26460 28588 26516
rect 28644 26460 28654 26516
rect 25554 26348 25564 26404
rect 25620 26348 26236 26404
rect 26292 26348 26302 26404
rect 22978 26236 22988 26292
rect 23044 26236 23996 26292
rect 24052 26236 24062 26292
rect 24658 26236 24668 26292
rect 24724 26236 25676 26292
rect 25732 26236 25742 26292
rect 23874 26124 23884 26180
rect 23940 26124 25116 26180
rect 25172 26124 25182 26180
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 23090 25788 23100 25844
rect 23156 25788 23884 25844
rect 23940 25788 23950 25844
rect 21970 25340 21980 25396
rect 22036 25340 23100 25396
rect 23156 25340 23166 25396
rect 15138 25228 15148 25284
rect 15204 25228 22092 25284
rect 22148 25228 22158 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 18834 24892 18844 24948
rect 18900 24892 19740 24948
rect 19796 24892 19806 24948
rect 4274 24668 4284 24724
rect 4340 24668 10780 24724
rect 10836 24668 10846 24724
rect 19282 24668 19292 24724
rect 19348 24668 20300 24724
rect 20356 24668 20366 24724
rect 15922 24556 15932 24612
rect 15988 24556 17500 24612
rect 17556 24556 17566 24612
rect 1922 24444 1932 24500
rect 1988 24444 1998 24500
rect 0 24276 800 24304
rect 1932 24276 1988 24444
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 0 24220 1988 24276
rect 19842 24220 19852 24276
rect 19908 24220 21420 24276
rect 21476 24220 21486 24276
rect 0 24192 800 24220
rect 19478 24108 19516 24164
rect 19572 24108 19582 24164
rect 12786 23996 12796 24052
rect 12852 23996 14028 24052
rect 14084 23996 14094 24052
rect 16146 23996 16156 24052
rect 16212 23996 21868 24052
rect 21924 23996 23212 24052
rect 23268 23996 23278 24052
rect 27010 23996 27020 24052
rect 27076 23996 28588 24052
rect 28644 23996 31948 24052
rect 31892 23940 31948 23996
rect 4274 23884 4284 23940
rect 4340 23884 11004 23940
rect 11060 23884 13580 23940
rect 13636 23884 13646 23940
rect 19842 23884 19852 23940
rect 19908 23884 20412 23940
rect 20468 23884 21308 23940
rect 21364 23884 21374 23940
rect 31892 23884 37660 23940
rect 37716 23884 37726 23940
rect 10882 23772 10892 23828
rect 10948 23772 12796 23828
rect 12852 23772 12862 23828
rect 13010 23772 13020 23828
rect 13076 23772 13468 23828
rect 13524 23772 18900 23828
rect 20290 23772 20300 23828
rect 20356 23772 21420 23828
rect 21476 23772 21486 23828
rect 22194 23772 22204 23828
rect 22260 23772 23436 23828
rect 23492 23772 23502 23828
rect 18844 23716 18900 23772
rect 13122 23660 13132 23716
rect 13188 23660 14140 23716
rect 14196 23660 14206 23716
rect 14354 23660 14364 23716
rect 14420 23660 17052 23716
rect 17108 23660 17612 23716
rect 17668 23660 17678 23716
rect 18834 23660 18844 23716
rect 18900 23660 18910 23716
rect 19506 23660 19516 23716
rect 19572 23660 20524 23716
rect 20580 23660 20590 23716
rect 0 23604 800 23632
rect 41200 23604 42000 23632
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 13682 23548 13692 23604
rect 13748 23548 15148 23604
rect 15204 23548 15214 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 41200 23520 42000 23548
rect 22082 23436 22092 23492
rect 22148 23436 25340 23492
rect 25396 23436 25406 23492
rect 13234 23324 13244 23380
rect 13300 23324 14588 23380
rect 14644 23324 14654 23380
rect 14802 23324 14812 23380
rect 14868 23324 15820 23380
rect 15876 23324 15886 23380
rect 16370 23100 16380 23156
rect 16436 23100 17836 23156
rect 17892 23100 18284 23156
rect 18340 23100 18350 23156
rect 20066 23100 20076 23156
rect 20132 23100 22428 23156
rect 22484 23100 22494 23156
rect 25666 23100 25676 23156
rect 25732 23100 26908 23156
rect 26964 23100 26974 23156
rect 17378 22876 17388 22932
rect 17444 22876 19068 22932
rect 19124 22876 20076 22932
rect 20132 22876 20142 22932
rect 17042 22764 17052 22820
rect 17108 22764 17948 22820
rect 18004 22764 21420 22820
rect 21476 22764 21486 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 20402 22652 20412 22708
rect 20468 22652 21196 22708
rect 21252 22652 22988 22708
rect 23044 22652 23054 22708
rect 18610 22540 18620 22596
rect 18676 22540 21756 22596
rect 21812 22540 25340 22596
rect 25396 22540 25406 22596
rect 14690 22428 14700 22484
rect 14756 22428 21644 22484
rect 21700 22428 26236 22484
rect 26292 22428 26302 22484
rect 28242 22428 28252 22484
rect 28308 22428 31948 22484
rect 31892 22372 31948 22428
rect 31892 22316 37660 22372
rect 37716 22316 37726 22372
rect 41200 22260 42000 22288
rect 19506 22204 19516 22260
rect 19572 22204 20524 22260
rect 20580 22204 21308 22260
rect 21364 22204 21374 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 41200 22176 42000 22204
rect 18834 22092 18844 22148
rect 18900 22092 19404 22148
rect 19460 22092 19470 22148
rect 18050 21980 18060 22036
rect 18116 21980 18620 22036
rect 18676 21980 19628 22036
rect 19684 21980 19694 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 21410 21868 21420 21924
rect 21476 21868 21756 21924
rect 21812 21868 23884 21924
rect 23940 21868 25116 21924
rect 25172 21868 25182 21924
rect 23762 21756 23772 21812
rect 23828 21756 26348 21812
rect 26404 21756 26414 21812
rect 23090 21644 23100 21700
rect 23156 21644 25676 21700
rect 25732 21644 25742 21700
rect 25890 21644 25900 21700
rect 25956 21644 28252 21700
rect 28308 21644 28318 21700
rect 18834 21532 18844 21588
rect 18900 21532 22876 21588
rect 22932 21532 22942 21588
rect 24882 21532 24892 21588
rect 24948 21532 25340 21588
rect 25396 21532 25406 21588
rect 28354 21532 28364 21588
rect 28420 21532 37660 21588
rect 37716 21532 37726 21588
rect 25554 21420 25564 21476
rect 25620 21420 26684 21476
rect 26740 21420 26750 21476
rect 18050 21308 18060 21364
rect 18116 21308 19516 21364
rect 19572 21308 23548 21364
rect 23604 21308 23614 21364
rect 26450 21308 26460 21364
rect 26516 21308 27132 21364
rect 27188 21308 27198 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 18386 21084 18396 21140
rect 18452 21084 19068 21140
rect 19124 21084 20076 21140
rect 20132 21084 24556 21140
rect 24612 21084 24622 21140
rect 19170 20972 19180 21028
rect 19236 20972 21868 21028
rect 21924 20972 22540 21028
rect 22596 20972 24332 21028
rect 24388 20972 24398 21028
rect 41200 20916 42000 20944
rect 20178 20860 20188 20916
rect 20244 20860 20972 20916
rect 21028 20860 22932 20916
rect 23314 20860 23324 20916
rect 23380 20860 26572 20916
rect 26628 20860 27468 20916
rect 27524 20860 27534 20916
rect 40002 20860 40012 20916
rect 40068 20860 42000 20916
rect 22876 20804 22932 20860
rect 41200 20832 42000 20860
rect 14466 20748 14476 20804
rect 14532 20748 15036 20804
rect 15092 20748 16492 20804
rect 16548 20748 17388 20804
rect 17444 20748 17454 20804
rect 17714 20748 17724 20804
rect 17780 20748 19292 20804
rect 19348 20748 19852 20804
rect 19908 20748 21532 20804
rect 21588 20748 21598 20804
rect 22876 20748 23660 20804
rect 23716 20748 23726 20804
rect 24882 20636 24892 20692
rect 24948 20636 27468 20692
rect 27524 20636 28028 20692
rect 28084 20636 28094 20692
rect 17714 20524 17724 20580
rect 17780 20524 18508 20580
rect 18564 20524 18574 20580
rect 18946 20524 18956 20580
rect 19012 20524 24556 20580
rect 24612 20524 25452 20580
rect 25508 20524 26348 20580
rect 26404 20524 26414 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 18610 20300 18620 20356
rect 18676 20300 19292 20356
rect 19348 20300 19358 20356
rect 23538 20300 23548 20356
rect 23604 20300 24556 20356
rect 24612 20300 25116 20356
rect 25172 20300 25182 20356
rect 19170 20188 19180 20244
rect 19236 20188 21756 20244
rect 21812 20188 22764 20244
rect 22820 20188 22830 20244
rect 24770 20188 24780 20244
rect 24836 20188 26124 20244
rect 26180 20188 27244 20244
rect 27300 20188 27310 20244
rect 15026 20076 15036 20132
rect 15092 20076 17388 20132
rect 17444 20076 17454 20132
rect 17602 20076 17612 20132
rect 17668 20076 17948 20132
rect 18004 20076 20020 20132
rect 22978 20076 22988 20132
rect 23044 20076 24444 20132
rect 24500 20076 24510 20132
rect 19964 20020 20020 20076
rect 4162 19964 4172 20020
rect 4228 19964 18508 20020
rect 18564 19964 19740 20020
rect 19796 19964 19806 20020
rect 19964 19964 23660 20020
rect 23716 19964 23726 20020
rect 12898 19852 12908 19908
rect 12964 19852 15260 19908
rect 15316 19852 15708 19908
rect 15764 19852 18172 19908
rect 18228 19852 18238 19908
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 17602 19516 17612 19572
rect 17668 19516 17948 19572
rect 18004 19516 18014 19572
rect 15474 19404 15484 19460
rect 15540 19404 18620 19460
rect 18676 19404 20860 19460
rect 20916 19404 20926 19460
rect 18162 19292 18172 19348
rect 18228 19292 20524 19348
rect 20580 19292 23436 19348
rect 23492 19292 23502 19348
rect 18722 19180 18732 19236
rect 18788 19180 19404 19236
rect 19460 19180 20300 19236
rect 20356 19180 21868 19236
rect 21924 19180 21934 19236
rect 17714 19068 17724 19124
rect 17780 19068 18452 19124
rect 23650 19068 23660 19124
rect 23716 19068 24556 19124
rect 24612 19068 24622 19124
rect 18396 19012 18452 19068
rect 18386 18956 18396 19012
rect 18452 18956 18462 19012
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 14802 18732 14812 18788
rect 14868 18732 17052 18788
rect 17108 18732 17118 18788
rect 22194 18620 22204 18676
rect 22260 18620 22270 18676
rect 22204 18564 22260 18620
rect 18050 18508 18060 18564
rect 18116 18508 20412 18564
rect 20468 18508 21196 18564
rect 21252 18508 21262 18564
rect 22204 18508 22988 18564
rect 23044 18508 24332 18564
rect 24388 18508 25340 18564
rect 25396 18508 25406 18564
rect 11778 18396 11788 18452
rect 11844 18396 12796 18452
rect 12852 18396 12862 18452
rect 14700 18396 18340 18452
rect 18498 18396 18508 18452
rect 18564 18396 19740 18452
rect 19796 18396 19806 18452
rect 21746 18396 21756 18452
rect 21812 18396 21980 18452
rect 22036 18396 23548 18452
rect 23604 18396 24108 18452
rect 24164 18396 24174 18452
rect 27570 18396 27580 18452
rect 27636 18396 28476 18452
rect 28532 18396 37660 18452
rect 37716 18396 37726 18452
rect 14700 18340 14756 18396
rect 18284 18340 18340 18396
rect 12338 18284 12348 18340
rect 12404 18284 14756 18340
rect 14914 18284 14924 18340
rect 14980 18284 16716 18340
rect 16772 18284 16782 18340
rect 18284 18284 19068 18340
rect 19124 18284 19134 18340
rect 19506 18284 19516 18340
rect 19572 18284 24220 18340
rect 24276 18284 24286 18340
rect 41200 18228 42000 18256
rect 18050 18172 18060 18228
rect 18116 18172 18844 18228
rect 18900 18172 23772 18228
rect 23828 18172 23838 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 41200 18144 42000 18172
rect 17266 18060 17276 18116
rect 17332 18060 19516 18116
rect 19572 18060 19582 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 20738 17948 20748 18004
rect 20804 17948 23100 18004
rect 23156 17948 23884 18004
rect 23940 17948 23950 18004
rect 18172 17836 18956 17892
rect 19012 17836 20412 17892
rect 20468 17836 26124 17892
rect 26180 17836 26190 17892
rect 18172 17780 18228 17836
rect 1922 17724 1932 17780
rect 1988 17724 1998 17780
rect 18162 17724 18172 17780
rect 18228 17724 18238 17780
rect 18386 17724 18396 17780
rect 18452 17724 19516 17780
rect 19572 17724 19582 17780
rect 0 17556 800 17584
rect 1932 17556 1988 17724
rect 4274 17612 4284 17668
rect 4340 17612 9996 17668
rect 10052 17612 10062 17668
rect 12786 17612 12796 17668
rect 12852 17612 13580 17668
rect 13636 17612 14364 17668
rect 14420 17612 14924 17668
rect 14980 17612 14990 17668
rect 41200 17556 42000 17584
rect 0 17500 1988 17556
rect 14242 17500 14252 17556
rect 14308 17500 15484 17556
rect 15540 17500 15550 17556
rect 16482 17500 16492 17556
rect 16548 17500 17164 17556
rect 17220 17500 17230 17556
rect 17714 17500 17724 17556
rect 17780 17500 18620 17556
rect 18676 17500 19068 17556
rect 19124 17500 19134 17556
rect 40002 17500 40012 17556
rect 40068 17500 42000 17556
rect 0 17472 800 17500
rect 41200 17472 42000 17500
rect 12114 17388 12124 17444
rect 12180 17388 14140 17444
rect 14196 17388 14206 17444
rect 14690 17388 14700 17444
rect 14756 17388 17500 17444
rect 17556 17388 17566 17444
rect 17724 17388 21980 17444
rect 22036 17388 22046 17444
rect 17724 17332 17780 17388
rect 15474 17276 15484 17332
rect 15540 17276 17780 17332
rect 19478 17276 19516 17332
rect 19572 17276 19582 17332
rect 24322 17276 24332 17332
rect 24388 17276 24668 17332
rect 24724 17276 24734 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 15698 17052 15708 17108
rect 15764 17052 16716 17108
rect 16772 17052 18508 17108
rect 18564 17052 24668 17108
rect 24724 17052 25340 17108
rect 25396 17052 25406 17108
rect 12796 16940 16268 16996
rect 16324 16940 16334 16996
rect 17714 16940 17724 16996
rect 17780 16940 18396 16996
rect 18452 16940 18462 16996
rect 0 16884 800 16912
rect 12796 16884 12852 16940
rect 0 16828 1932 16884
rect 1988 16828 1998 16884
rect 4274 16828 4284 16884
rect 4340 16828 12796 16884
rect 12852 16828 12862 16884
rect 0 16800 800 16828
rect 9986 16716 9996 16772
rect 10052 16716 15148 16772
rect 15204 16716 15214 16772
rect 17826 16716 17836 16772
rect 17892 16716 19068 16772
rect 19124 16716 19134 16772
rect 23986 16716 23996 16772
rect 24052 16716 25004 16772
rect 25060 16716 25070 16772
rect 28578 16716 28588 16772
rect 28644 16716 37660 16772
rect 37716 16716 37726 16772
rect 14690 16604 14700 16660
rect 14756 16604 18732 16660
rect 18788 16604 18798 16660
rect 19506 16604 19516 16660
rect 19572 16604 24220 16660
rect 24276 16604 26572 16660
rect 26628 16604 26638 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 24546 16268 24556 16324
rect 24612 16268 25452 16324
rect 25508 16268 25518 16324
rect 19282 16156 19292 16212
rect 19348 16156 20524 16212
rect 20580 16156 21196 16212
rect 21252 16156 21262 16212
rect 4274 16044 4284 16100
rect 4340 16044 11228 16100
rect 11284 16044 13692 16100
rect 13748 16044 13758 16100
rect 17154 16044 17164 16100
rect 17220 16044 18956 16100
rect 19012 16044 19022 16100
rect 22866 16044 22876 16100
rect 22932 16044 23548 16100
rect 23604 16044 24444 16100
rect 24500 16044 24510 16100
rect 13794 15932 13804 15988
rect 13860 15932 15260 15988
rect 15316 15932 15596 15988
rect 15652 15932 16156 15988
rect 16212 15932 16828 15988
rect 16884 15932 16894 15988
rect 23986 15932 23996 15988
rect 24052 15932 28588 15988
rect 28644 15932 28654 15988
rect 13346 15820 13356 15876
rect 13412 15820 14588 15876
rect 14644 15820 14654 15876
rect 18162 15820 18172 15876
rect 18228 15820 18956 15876
rect 19012 15820 19022 15876
rect 19618 15820 19628 15876
rect 19684 15820 20636 15876
rect 20692 15820 21644 15876
rect 21700 15820 22428 15876
rect 22484 15820 22494 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 0 15540 800 15568
rect 0 15484 1932 15540
rect 1988 15484 1998 15540
rect 0 15456 800 15484
rect 20290 15260 20300 15316
rect 20356 15260 21196 15316
rect 21252 15260 22428 15316
rect 22484 15260 22494 15316
rect 25554 15260 25564 15316
rect 25620 15260 27580 15316
rect 27636 15260 27646 15316
rect 23538 15148 23548 15204
rect 23604 15148 25788 15204
rect 25844 15148 25854 15204
rect 13570 15036 13580 15092
rect 13636 15036 14588 15092
rect 14644 15036 16156 15092
rect 16212 15036 16222 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 22194 14812 22204 14868
rect 22260 14812 23436 14868
rect 23492 14812 23502 14868
rect 21634 14700 21644 14756
rect 21700 14700 22652 14756
rect 22708 14700 22718 14756
rect 19506 14588 19516 14644
rect 19572 14588 21868 14644
rect 21924 14588 24332 14644
rect 24388 14588 24398 14644
rect 27570 14588 27580 14644
rect 27636 14588 28588 14644
rect 28644 14588 28654 14644
rect 20290 14476 20300 14532
rect 20356 14476 22540 14532
rect 22596 14476 23212 14532
rect 23268 14476 23278 14532
rect 15922 14252 15932 14308
rect 15988 14252 17388 14308
rect 17444 14252 17454 14308
rect 22978 14252 22988 14308
rect 23044 14252 24220 14308
rect 24276 14252 24286 14308
rect 21298 14140 21308 14196
rect 21364 14140 22092 14196
rect 22148 14140 22158 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 17938 13804 17948 13860
rect 18004 13804 19180 13860
rect 19236 13804 19246 13860
rect 19506 13804 19516 13860
rect 19572 13804 20636 13860
rect 20692 13804 20702 13860
rect 17602 13692 17612 13748
rect 17668 13692 20412 13748
rect 20468 13692 20478 13748
rect 15698 13580 15708 13636
rect 15764 13580 16492 13636
rect 16548 13580 16940 13636
rect 16996 13580 17006 13636
rect 14354 13468 14364 13524
rect 14420 13468 17500 13524
rect 17556 13468 17566 13524
rect 23762 13468 23772 13524
rect 23828 13468 24668 13524
rect 24724 13468 25228 13524
rect 25284 13468 25564 13524
rect 25620 13468 25630 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 16706 13020 16716 13076
rect 16772 13020 17724 13076
rect 17780 13020 17790 13076
rect 18498 12796 18508 12852
rect 18564 12796 20076 12852
rect 20132 12796 20142 12852
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 24882 5180 24892 5236
rect 24948 5180 26124 5236
rect 26180 5180 26190 5236
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 18834 4060 18844 4116
rect 18900 4060 20076 4116
rect 20132 4060 20142 4116
rect 24210 4060 24220 4116
rect 24276 4060 26236 4116
rect 26292 4060 26302 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 25666 3612 25676 3668
rect 25732 3612 29372 3668
rect 29428 3612 29438 3668
rect 16146 3388 16156 3444
rect 16212 3388 18508 3444
rect 18564 3388 18574 3444
rect 20178 3388 20188 3444
rect 20244 3388 21756 3444
rect 21812 3388 21822 3444
rect 23538 3388 23548 3444
rect 23604 3388 25564 3444
rect 25620 3388 25630 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19516 24108 19572 24164
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19516 17276 19572 17332
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 19516 24164 19572 24174
rect 19516 17332 19572 24108
rect 19516 17266 19572 17276
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16352 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18928 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21392 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _112_
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23408 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1698175906
transform 1 0 20048 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform -1 0 19376 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17920 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698175906
transform 1 0 18144 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform -1 0 18704 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19824 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _121_
timestamp 1698175906
transform -1 0 22512 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _122_
timestamp 1698175906
transform 1 0 19600 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19824 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _124_
timestamp 1698175906
transform -1 0 20944 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18928 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _126_
timestamp 1698175906
transform -1 0 22176 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _127_
timestamp 1698175906
transform 1 0 24416 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _128_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _129_
timestamp 1698175906
transform 1 0 25200 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _130_
timestamp 1698175906
transform 1 0 26768 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform 1 0 18368 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _132_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19824 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18144 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _134_
timestamp 1698175906
transform -1 0 20496 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _135_
timestamp 1698175906
transform 1 0 24304 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _136_
timestamp 1698175906
transform -1 0 26768 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14560 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15232 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _139_
timestamp 1698175906
transform 1 0 23744 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _140_
timestamp 1698175906
transform 1 0 19376 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _141_
timestamp 1698175906
transform -1 0 20608 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _142_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19152 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _143_
timestamp 1698175906
transform -1 0 20048 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _144_
timestamp 1698175906
transform -1 0 17584 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _145_
timestamp 1698175906
transform -1 0 19040 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _146_
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _147_
timestamp 1698175906
transform -1 0 18256 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _148_
timestamp 1698175906
transform 1 0 18144 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _149_
timestamp 1698175906
transform -1 0 24192 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _150_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21280 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _151_
timestamp 1698175906
transform 1 0 17248 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _152_
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _153_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21840 0 1 18816
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _154_
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _155_
timestamp 1698175906
transform -1 0 25088 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _156_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19376 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _157_
timestamp 1698175906
transform 1 0 18704 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698175906
transform 1 0 20384 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _159_
timestamp 1698175906
transform 1 0 22400 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _160_
timestamp 1698175906
transform 1 0 22400 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _161_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21840 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _162_
timestamp 1698175906
transform -1 0 19600 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _163_
timestamp 1698175906
transform -1 0 18144 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _164_
timestamp 1698175906
transform -1 0 19824 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _165_
timestamp 1698175906
transform -1 0 19152 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _166_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21952 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _167_
timestamp 1698175906
transform -1 0 16352 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _168_
timestamp 1698175906
transform -1 0 15120 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _169_
timestamp 1698175906
transform -1 0 22624 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _170_
timestamp 1698175906
transform -1 0 17136 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _171_
timestamp 1698175906
transform -1 0 16912 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _172_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22512 0 1 20384
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _173_
timestamp 1698175906
transform 1 0 24192 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _174_
timestamp 1698175906
transform -1 0 26096 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _175_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 26992 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _176_
timestamp 1698175906
transform -1 0 13104 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _177_
timestamp 1698175906
transform -1 0 16576 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _178_
timestamp 1698175906
transform 1 0 13888 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _179_
timestamp 1698175906
transform -1 0 15680 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _180_
timestamp 1698175906
transform 1 0 18256 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _181_
timestamp 1698175906
transform -1 0 17360 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _182_
timestamp 1698175906
transform -1 0 14000 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _183_
timestamp 1698175906
transform -1 0 14896 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _184_
timestamp 1698175906
transform -1 0 15456 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _185_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15232 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _186_
timestamp 1698175906
transform 1 0 21616 0 1 17248
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _187_
timestamp 1698175906
transform 1 0 23744 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _188_
timestamp 1698175906
transform -1 0 24864 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _189_
timestamp 1698175906
transform 1 0 25088 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _190_
timestamp 1698175906
transform 1 0 25760 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _191_
timestamp 1698175906
transform 1 0 27104 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _192_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25984 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _193_
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _194_
timestamp 1698175906
transform 1 0 14112 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _195_
timestamp 1698175906
transform 1 0 27888 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _196_
timestamp 1698175906
transform -1 0 27888 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _197_
timestamp 1698175906
transform 1 0 23744 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _198_
timestamp 1698175906
transform 1 0 22848 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _199_
timestamp 1698175906
transform -1 0 25984 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _200_
timestamp 1698175906
transform 1 0 25984 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _201_
timestamp 1698175906
transform 1 0 16016 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _202_
timestamp 1698175906
transform 1 0 17024 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _203_
timestamp 1698175906
transform -1 0 18032 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _204_
timestamp 1698175906
transform 1 0 15456 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _205_
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _206_
timestamp 1698175906
transform 1 0 23184 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _207_
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _208_
timestamp 1698175906
transform 1 0 21840 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _209_
timestamp 1698175906
transform -1 0 18144 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _210_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18480 0 1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _211_
timestamp 1698175906
transform -1 0 18368 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _212_
timestamp 1698175906
transform 1 0 20384 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _213_
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17584 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 25536 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 11424 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 11984 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 18368 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 15008 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 25200 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 17248 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 13664 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 25200 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform -1 0 14112 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform -1 0 14336 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform -1 0 13104 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 25536 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 25424 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform -1 0 14112 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 25536 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform 1 0 21952 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 24528 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform -1 0 15904 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform 1 0 13440 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 21616 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698175906
transform 1 0 16016 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform -1 0 22400 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _242_
timestamp 1698175906
transform -1 0 25760 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _243_
timestamp 1698175906
transform 1 0 25984 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__B dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17360 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__A3
timestamp 1698175906
transform 1 0 15456 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__A2
timestamp 1698175906
transform 1 0 21728 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__B
timestamp 1698175906
transform 1 0 23296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 20944 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 25312 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 14896 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform -1 0 16352 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 21840 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 18480 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform -1 0 25536 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform -1 0 21168 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 16576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform -1 0 17696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 25312 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 14112 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 14560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 13552 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 14336 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 25984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform -1 0 25984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 24304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform 1 0 16688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 21392 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform 1 0 19488 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform -1 0 22848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 18480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18704 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 23744 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 19264 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_164 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19712 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_168 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_198
timestamp 1698175906
transform 1 0 23520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_202
timestamp 1698175906
transform 1 0 23968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_266
timestamp 1698175906
transform 1 0 31136 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_270
timestamp 1698175906
transform 1 0 31584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698175906
transform 1 0 18144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_154
timestamp 1698175906
transform 1 0 18592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_156
timestamp 1698175906
transform 1 0 18816 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_183 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21840 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_199
timestamp 1698175906
transform 1 0 23632 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 28000 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 31584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_209
timestamp 1698175906
transform 1 0 24752 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_237
timestamp 1698175906
transform 1 0 27888 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_174
timestamp 1698175906
transform 1 0 20832 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_177
timestamp 1698175906
transform 1 0 21168 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698175906
transform 1 0 24752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_123
timestamp 1698175906
transform 1 0 15120 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_131
timestamp 1698175906
transform 1 0 16016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_135
timestamp 1698175906
transform 1 0 16464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_139
timestamp 1698175906
transform 1 0 16912 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_143
timestamp 1698175906
transform 1 0 17360 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_206
timestamp 1698175906
transform 1 0 24416 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_238
timestamp 1698175906
transform 1 0 28000 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_242
timestamp 1698175906
transform 1 0 28448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698175906
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_104
timestamp 1698175906
transform 1 0 12992 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_137
timestamp 1698175906
transform 1 0 16688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698175906
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_153
timestamp 1698175906
transform 1 0 18480 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_157
timestamp 1698175906
transform 1 0 18928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_159
timestamp 1698175906
transform 1 0 19152 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_173
timestamp 1698175906
transform 1 0 20720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_177
timestamp 1698175906
transform 1 0 21168 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_218
timestamp 1698175906
transform 1 0 25760 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_250
timestamp 1698175906
transform 1 0 29344 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_266
timestamp 1698175906
transform 1 0 31136 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_274
timestamp 1698175906
transform 1 0 32032 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_278
timestamp 1698175906
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_125
timestamp 1698175906
transform 1 0 15344 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_160
timestamp 1698175906
transform 1 0 19264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_164
timestamp 1698175906
transform 1 0 19712 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698175906
transform 1 0 20608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_185
timestamp 1698175906
transform 1 0 22064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_187
timestamp 1698175906
transform 1 0 22288 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_202
timestamp 1698175906
transform 1 0 23968 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_204
timestamp 1698175906
transform 1 0 24192 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_236
timestamp 1698175906
transform 1 0 27776 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_80
timestamp 1698175906
transform 1 0 10304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_84
timestamp 1698175906
transform 1 0 10752 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_86
timestamp 1698175906
transform 1 0 10976 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_116
timestamp 1698175906
transform 1 0 14336 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_120
timestamp 1698175906
transform 1 0 14784 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_146
timestamp 1698175906
transform 1 0 17696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_152
timestamp 1698175906
transform 1 0 18368 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_168
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_172
timestamp 1698175906
transform 1 0 20608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_192
timestamp 1698175906
transform 1 0 22848 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698175906
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_226
timestamp 1698175906
transform 1 0 26656 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_258
timestamp 1698175906
transform 1 0 30240 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_274
timestamp 1698175906
transform 1 0 32032 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698175906
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_28
timestamp 1698175906
transform 1 0 4480 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698175906
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_126
timestamp 1698175906
transform 1 0 15456 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_134
timestamp 1698175906
transform 1 0 16352 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_136
timestamp 1698175906
transform 1 0 16576 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_143
timestamp 1698175906
transform 1 0 17360 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_151
timestamp 1698175906
transform 1 0 18256 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_164
timestamp 1698175906
transform 1 0 19712 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_168
timestamp 1698175906
transform 1 0 20160 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_185
timestamp 1698175906
transform 1 0 22064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_187
timestamp 1698175906
transform 1 0 22288 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_194
timestamp 1698175906
transform 1 0 23072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_198
timestamp 1698175906
transform 1 0 23520 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_205
timestamp 1698175906
transform 1 0 24304 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_209
timestamp 1698175906
transform 1 0 24752 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_211
timestamp 1698175906
transform 1 0 24976 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_220
timestamp 1698175906
transform 1 0 25984 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_236
timestamp 1698175906
transform 1 0 27776 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 4480 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_88
timestamp 1698175906
transform 1 0 11200 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_96
timestamp 1698175906
transform 1 0 12096 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_100
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_130
timestamp 1698175906
transform 1 0 15904 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_136
timestamp 1698175906
transform 1 0 16576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_206
timestamp 1698175906
transform 1 0 24416 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_245
timestamp 1698175906
transform 1 0 28784 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698175906
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_69
timestamp 1698175906
transform 1 0 9072 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_73
timestamp 1698175906
transform 1 0 9520 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_75
timestamp 1698175906
transform 1 0 9744 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_111
timestamp 1698175906
transform 1 0 13776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_124
timestamp 1698175906
transform 1 0 15232 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_128
timestamp 1698175906
transform 1 0 15680 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_136
timestamp 1698175906
transform 1 0 16576 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_159
timestamp 1698175906
transform 1 0 19152 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698175906
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_224
timestamp 1698175906
transform 1 0 26432 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_240
timestamp 1698175906
transform 1 0 28224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_88
timestamp 1698175906
transform 1 0 11200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_119
timestamp 1698175906
transform 1 0 14672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_123
timestamp 1698175906
transform 1 0 15120 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_179
timestamp 1698175906
transform 1 0 21392 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_181
timestamp 1698175906
transform 1 0 21616 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_197
timestamp 1698175906
transform 1 0 23408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_214
timestamp 1698175906
transform 1 0 25312 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_244
timestamp 1698175906
transform 1 0 28672 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698175906
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_115
timestamp 1698175906
transform 1 0 14224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_119
timestamp 1698175906
transform 1 0 14672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_128
timestamp 1698175906
transform 1 0 15680 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_136
timestamp 1698175906
transform 1 0 16576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_138
timestamp 1698175906
transform 1 0 16800 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_163
timestamp 1698175906
transform 1 0 19600 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_181
timestamp 1698175906
transform 1 0 21616 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_236
timestamp 1698175906
transform 1 0 27776 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_88
timestamp 1698175906
transform 1 0 11200 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_92
timestamp 1698175906
transform 1 0 11648 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_94
timestamp 1698175906
transform 1 0 11872 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_130
timestamp 1698175906
transform 1 0 15904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_134
timestamp 1698175906
transform 1 0 16352 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_138
timestamp 1698175906
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_150
timestamp 1698175906
transform 1 0 18144 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_152
timestamp 1698175906
transform 1 0 18368 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_218
timestamp 1698175906
transform 1 0 25760 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_222
timestamp 1698175906
transform 1 0 26208 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_254
timestamp 1698175906
transform 1 0 29792 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_270
timestamp 1698175906
transform 1 0 31584 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 40320 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_115
timestamp 1698175906
transform 1 0 14224 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_117
timestamp 1698175906
transform 1 0 14448 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_130
timestamp 1698175906
transform 1 0 15904 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698175906
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_212
timestamp 1698175906
transform 1 0 25088 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698175906
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_148
timestamp 1698175906
transform 1 0 17920 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_186
timestamp 1698175906
transform 1 0 22176 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_190
timestamp 1698175906
transform 1 0 22624 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_243
timestamp 1698175906
transform 1 0 28560 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_275
timestamp 1698175906
transform 1 0 32144 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_111
timestamp 1698175906
transform 1 0 13776 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_113
timestamp 1698175906
transform 1 0 14000 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_116
timestamp 1698175906
transform 1 0 14336 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698175906
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_210
timestamp 1698175906
transform 1 0 24864 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_212
timestamp 1698175906
transform 1 0 25088 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_242
timestamp 1698175906
transform 1 0 28448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_80
timestamp 1698175906
transform 1 0 10304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_84
timestamp 1698175906
transform 1 0 10752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_123
timestamp 1698175906
transform 1 0 15120 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_127
timestamp 1698175906
transform 1 0 15568 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698175906
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_158
timestamp 1698175906
transform 1 0 19040 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_218
timestamp 1698175906
transform 1 0 25760 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_232
timestamp 1698175906
transform 1 0 27328 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_264
timestamp 1698175906
transform 1 0 30912 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 40320 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_69
timestamp 1698175906
transform 1 0 9072 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_85
timestamp 1698175906
transform 1 0 10864 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_93
timestamp 1698175906
transform 1 0 11760 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_97
timestamp 1698175906
transform 1 0 12208 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_99
timestamp 1698175906
transform 1 0 12432 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_120
timestamp 1698175906
transform 1 0 14784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_151
timestamp 1698175906
transform 1 0 18256 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_173
timestamp 1698175906
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_190
timestamp 1698175906
transform 1 0 22624 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_206
timestamp 1698175906
transform 1 0 24416 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 4480 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 8064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698175906
transform 1 0 10304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_84
timestamp 1698175906
transform 1 0 10752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_114
timestamp 1698175906
transform 1 0 14112 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_118
timestamp 1698175906
transform 1 0 14560 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_134
timestamp 1698175906
transform 1 0 16352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_150
timestamp 1698175906
transform 1 0 18144 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_158
timestamp 1698175906
transform 1 0 19040 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_172
timestamp 1698175906
transform 1 0 20608 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_176
timestamp 1698175906
transform 1 0 21056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_188
timestamp 1698175906
transform 1 0 22400 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_204
timestamp 1698175906
transform 1 0 24192 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698175906
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698175906
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_193
timestamp 1698175906
transform 1 0 22960 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_201
timestamp 1698175906
transform 1 0 23856 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_205
timestamp 1698175906
transform 1 0 24304 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_212
timestamp 1698175906
transform 1 0 25088 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_104
timestamp 1698175906
transform 1 0 12992 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_112
timestamp 1698175906
transform 1 0 13888 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_116
timestamp 1698175906
transform 1 0 14336 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_118
timestamp 1698175906
transform 1 0 14560 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_123
timestamp 1698175906
transform 1 0 15120 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_131
timestamp 1698175906
transform 1 0 16016 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_135
timestamp 1698175906
transform 1 0 16464 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698175906
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_150
timestamp 1698175906
transform 1 0 18144 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_181
timestamp 1698175906
transform 1 0 21616 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_185
timestamp 1698175906
transform 1 0 22064 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_189
timestamp 1698175906
transform 1 0 22512 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_191
timestamp 1698175906
transform 1 0 22736 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698175906
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_226
timestamp 1698175906
transform 1 0 26656 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_258
timestamp 1698175906
transform 1 0 30240 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_274
timestamp 1698175906
transform 1 0 32032 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698175906
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_141
timestamp 1698175906
transform 1 0 17136 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_171
timestamp 1698175906
transform 1 0 20496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_182
timestamp 1698175906
transform 1 0 21728 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_104
timestamp 1698175906
transform 1 0 12992 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_108
timestamp 1698175906
transform 1 0 13440 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698175906
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_146
timestamp 1698175906
transform 1 0 17696 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_188
timestamp 1698175906
transform 1 0 22400 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_192
timestamp 1698175906
transform 1 0 22848 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698175906
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_216
timestamp 1698175906
transform 1 0 25536 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_220
timestamp 1698175906
transform 1 0 25984 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_252
timestamp 1698175906
transform 1 0 29568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_268
timestamp 1698175906
transform 1 0 31360 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_123
timestamp 1698175906
transform 1 0 15120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_125
timestamp 1698175906
transform 1 0 15344 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_139
timestamp 1698175906
transform 1 0 16912 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_143
timestamp 1698175906
transform 1 0 17360 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_159
timestamp 1698175906
transform 1 0 19152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_165
timestamp 1698175906
transform 1 0 19824 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_169
timestamp 1698175906
transform 1 0 20272 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_6
timestamp 1698175906
transform 1 0 2016 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_22
timestamp 1698175906
transform 1 0 3808 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_30
timestamp 1698175906
transform 1 0 4704 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_168
timestamp 1698175906
transform 1 0 20160 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_195
timestamp 1698175906
transform 1 0 23184 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698175906
transform 1 0 24080 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 25536 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_243
timestamp 1698175906
transform 1 0 28560 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698175906
transform 1 0 32144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_169
timestamp 1698175906
transform 1 0 20272 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_206
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_210
timestamp 1698175906
transform 1 0 24864 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_237
timestamp 1698175906
transform 1 0 27888 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_266
timestamp 1698175906
transform 1 0 31136 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_270
timestamp 1698175906
transform 1 0 31584 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita59_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 2016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita59_26
timestamp 1698175906
transform -1 0 20272 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 18928 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 24976 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 24976 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 28560 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform -1 0 4480 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform -1 0 4480 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform -1 0 4480 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 4480 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 16912 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 20272 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 21280 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 24864 41200 24976 42000 0 FreeSans 448 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 25536 41200 25648 42000 0 FreeSans 448 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 18816 41200 18928 42000 0 FreeSans 448 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 0 15456 800 15568 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 41200 17472 42000 17584 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 16800 41200 16912 42000 0 FreeSans 448 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 16128 41200 16240 42000 0 FreeSans 448 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 20160 41200 20272 42000 0 FreeSans 448 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 26208 41200 26320 42000 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 14616 28280 14616 28280 0 _000_
rlabel metal2 26264 21952 26264 21952 0 _001_
rlabel metal2 13160 23464 13160 23464 0 _002_
rlabel metal2 13384 15624 13384 15624 0 _003_
rlabel metal2 12152 17472 12152 17472 0 _004_
rlabel metal2 26488 17192 26488 17192 0 _005_
rlabel metal2 26320 18536 26320 18536 0 _006_
rlabel metal3 13944 23352 13944 23352 0 _007_
rlabel metal2 26488 21112 26488 21112 0 _008_
rlabel metal2 23016 26936 23016 26936 0 _009_
rlabel metal2 25480 14672 25480 14672 0 _010_
rlabel metal2 14728 17136 14728 17136 0 _011_
rlabel metal2 14392 13552 14392 13552 0 _012_
rlabel metal2 22456 13832 22456 13832 0 _013_
rlabel metal2 16968 14840 16968 14840 0 _014_
rlabel metal2 21448 27496 21448 27496 0 _015_
rlabel metal3 19320 12824 19320 12824 0 _016_
rlabel metal2 26488 23576 26488 23576 0 _017_
rlabel metal3 14728 18368 14728 18368 0 _018_
rlabel metal2 15736 19992 15736 19992 0 _019_
rlabel metal2 19432 25536 19432 25536 0 _020_
rlabel metal2 15960 24304 15960 24304 0 _021_
rlabel metal3 25480 26936 25480 26936 0 _022_
rlabel metal2 22120 13608 22120 13608 0 _023_
rlabel metal2 18200 27496 18200 27496 0 _024_
rlabel metal2 14840 26712 14840 26712 0 _025_
rlabel metal2 24920 25760 24920 25760 0 _026_
rlabel metal3 20160 15848 20160 15848 0 _027_
rlabel metal2 19320 17192 19320 17192 0 _028_
rlabel metal2 21336 15512 21336 15512 0 _029_
rlabel metal2 22792 14812 22792 14812 0 _030_
rlabel metal3 22176 14728 22176 14728 0 _031_
rlabel metal2 19320 19824 19320 19824 0 _032_
rlabel metal3 20552 28448 20552 28448 0 _033_
rlabel metal2 18984 28168 18984 28168 0 _034_
rlabel metal2 22288 28616 22288 28616 0 _035_
rlabel metal2 14952 27384 14952 27384 0 _036_
rlabel metal2 16576 28392 16576 28392 0 _037_
rlabel metal2 16632 27496 16632 27496 0 _038_
rlabel metal2 27496 21112 27496 21112 0 _039_
rlabel metal3 18200 17528 18200 17528 0 _040_
rlabel metal3 26152 21448 26152 21448 0 _041_
rlabel metal2 12824 24080 12824 24080 0 _042_
rlabel metal2 14840 23576 14840 23576 0 _043_
rlabel metal2 14560 17864 14560 17864 0 _044_
rlabel metal2 14728 16352 14728 16352 0 _045_
rlabel metal3 16520 15960 16520 15960 0 _046_
rlabel metal2 14056 16184 14056 16184 0 _047_
rlabel metal2 15008 16072 15008 16072 0 _048_
rlabel metal2 25032 16408 25032 16408 0 _049_
rlabel metal2 24304 16072 24304 16072 0 _050_
rlabel metal3 25032 16296 25032 16296 0 _051_
rlabel metal2 25816 16912 25816 16912 0 _052_
rlabel metal2 27160 19208 27160 19208 0 _053_
rlabel metal2 14504 23016 14504 23016 0 _054_
rlabel metal2 27944 21560 27944 21560 0 _055_
rlabel metal3 23520 26264 23520 26264 0 _056_
rlabel metal2 26152 15456 26152 15456 0 _057_
rlabel metal2 16520 17304 16520 17304 0 _058_
rlabel metal2 18256 13720 18256 13720 0 _059_
rlabel metal2 17416 14056 17416 14056 0 _060_
rlabel metal2 23464 14784 23464 14784 0 _061_
rlabel metal2 22008 15512 22008 15512 0 _062_
rlabel metal2 19096 16520 19096 16520 0 _063_
rlabel metal2 18200 15624 18200 15624 0 _064_
rlabel metal2 21336 27720 21336 27720 0 _065_
rlabel metal2 23912 22120 23912 22120 0 _066_
rlabel metal3 23688 18536 23688 18536 0 _067_
rlabel metal3 20720 20776 20720 20776 0 _068_
rlabel metal2 22008 22344 22008 22344 0 _069_
rlabel metal2 21112 18816 21112 18816 0 _070_
rlabel metal2 23128 18200 23128 18200 0 _071_
rlabel metal3 22904 14504 22904 14504 0 _072_
rlabel metal3 20440 22232 20440 22232 0 _073_
rlabel metal2 12992 23912 12992 23912 0 _074_
rlabel metal2 19768 13776 19768 13776 0 _075_
rlabel metal2 20104 22176 20104 22176 0 _076_
rlabel metal3 19152 18424 19152 18424 0 _077_
rlabel metal3 19040 13720 19040 13720 0 _078_
rlabel metal3 21840 15288 21840 15288 0 _079_
rlabel metal2 23352 16968 23352 16968 0 _080_
rlabel metal2 20328 19264 20328 19264 0 _081_
rlabel metal2 18648 19376 18648 19376 0 _082_
rlabel metal2 14728 22792 14728 22792 0 _083_
rlabel metal2 28056 21000 28056 21000 0 _084_
rlabel metal2 21784 22512 21784 22512 0 _085_
rlabel metal3 26320 23128 26320 23128 0 _086_
rlabel metal2 26712 23016 26712 23016 0 _087_
rlabel metal2 19768 24024 19768 24024 0 _088_
rlabel metal2 24584 20272 24584 20272 0 _089_
rlabel metal3 18760 22904 18760 22904 0 _090_
rlabel metal2 20440 22568 20440 22568 0 _091_
rlabel metal2 27272 20776 27272 20776 0 _092_
rlabel metal2 15512 20328 15512 20328 0 _093_
rlabel metal2 19544 16688 19544 16688 0 _094_
rlabel metal2 19880 23968 19880 23968 0 _095_
rlabel metal3 19320 24920 19320 24920 0 _096_
rlabel metal2 23912 16296 23912 16296 0 _097_
rlabel metal2 14392 23744 14392 23744 0 _098_
rlabel metal3 17360 23128 17360 23128 0 _099_
rlabel metal2 17752 19824 17752 19824 0 _100_
rlabel metal2 18872 21280 18872 21280 0 _101_
rlabel metal2 24584 25536 24584 25536 0 _102_
rlabel metal2 23128 21952 23128 21952 0 _103_
rlabel metal3 22848 23800 22848 23800 0 _104_
rlabel metal2 23912 19208 23912 19208 0 _105_
rlabel metal2 24584 26264 24584 26264 0 _106_
rlabel metal3 2478 28280 2478 28280 0 clk
rlabel metal2 22344 18368 22344 18368 0 clknet_0_clk
rlabel metal2 24528 14616 24528 14616 0 clknet_1_0__leaf_clk
rlabel metal2 25480 27384 25480 27384 0 clknet_1_1__leaf_clk
rlabel metal3 14784 20776 14784 20776 0 dut59.count\[0\]
rlabel metal2 14840 20468 14840 20468 0 dut59.count\[1\]
rlabel metal2 21224 18480 21224 18480 0 dut59.count\[2\]
rlabel metal2 18648 22176 18648 22176 0 dut59.count\[3\]
rlabel metal2 28616 21224 28616 21224 0 net1
rlabel metal2 11256 15624 11256 15624 0 net10
rlabel metal2 10024 17248 10024 17248 0 net11
rlabel metal2 28616 16352 28616 16352 0 net12
rlabel metal2 28280 22064 28280 22064 0 net13
rlabel metal2 12824 16800 12824 16800 0 net14
rlabel metal3 16744 13608 16744 13608 0 net15
rlabel metal2 16800 27720 16800 27720 0 net16
rlabel metal2 16408 27720 16408 27720 0 net17
rlabel metal2 20328 27832 20328 27832 0 net18
rlabel metal2 28616 32256 28616 32256 0 net19
rlabel metal2 28504 18368 28504 18368 0 net2
rlabel metal3 28112 14616 28112 14616 0 net20
rlabel metal2 27048 23688 27048 23688 0 net21
rlabel metal2 20664 28112 20664 28112 0 net22
rlabel metal2 20720 13048 20720 13048 0 net23
rlabel metal2 24584 5964 24584 5964 0 net24
rlabel metal3 1246 36344 1246 36344 0 net25
rlabel metal2 19992 38248 19992 38248 0 net26
rlabel metal2 11032 24248 11032 24248 0 net3
rlabel metal2 18872 14616 18872 14616 0 net4
rlabel metal2 25312 13832 25312 13832 0 net5
rlabel metal2 25032 27776 25032 27776 0 net6
rlabel metal2 28280 26992 28280 26992 0 net7
rlabel metal2 25592 13608 25592 13608 0 net8
rlabel metal2 10976 23016 10976 23016 0 net9
rlabel metal2 40040 21112 40040 21112 0 segm[10]
rlabel metal3 40642 18200 40642 18200 0 segm[11]
rlabel metal3 1358 23576 1358 23576 0 segm[12]
rlabel metal2 18872 2422 18872 2422 0 segm[13]
rlabel metal2 24920 2982 24920 2982 0 segm[1]
rlabel metal2 24920 39914 24920 39914 0 segm[2]
rlabel metal2 25592 39186 25592 39186 0 segm[3]
rlabel metal2 24248 2422 24248 2422 0 segm[4]
rlabel metal3 1358 24248 1358 24248 0 segm[6]
rlabel metal3 1358 15512 1358 15512 0 segm[7]
rlabel metal3 1358 17528 1358 17528 0 segm[8]
rlabel metal2 40040 17640 40040 17640 0 segm[9]
rlabel metal2 40040 22344 40040 22344 0 sel[0]
rlabel metal3 1358 16856 1358 16856 0 sel[10]
rlabel metal2 16184 2086 16184 2086 0 sel[11]
rlabel metal2 16856 39746 16856 39746 0 sel[1]
rlabel metal2 16184 39354 16184 39354 0 sel[2]
rlabel metal2 20216 39354 20216 39354 0 sel[3]
rlabel metal2 26264 39746 26264 39746 0 sel[4]
rlabel metal2 25592 1190 25592 1190 0 sel[5]
rlabel metal2 40040 23800 40040 23800 0 sel[6]
rlabel metal2 22232 39746 22232 39746 0 sel[7]
rlabel metal2 20216 2086 20216 2086 0 sel[8]
rlabel metal2 23576 2086 23576 2086 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
