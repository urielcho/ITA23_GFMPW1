magic
tech gf180mcuD
magscale 1 5
timestamp 1699643053
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 11215 19137 11241 19143
rect 11215 19105 11241 19111
rect 14687 19137 14713 19143
rect 14687 19105 14713 19111
rect 12833 19055 12839 19081
rect 12865 19055 12871 19081
rect 10873 18999 10879 19025
rect 10905 18999 10911 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 14289 18999 14295 19025
rect 14321 18999 14327 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 12223 18745 12249 18751
rect 12223 18713 12249 18719
rect 13119 18745 13145 18751
rect 13119 18713 13145 18719
rect 12833 18607 12839 18633
rect 12865 18607 12871 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 11999 18353 12025 18359
rect 11999 18321 12025 18327
rect 12945 18215 12951 18241
rect 12977 18215 12983 18241
rect 20119 18129 20145 18135
rect 20119 18097 20145 18103
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 967 13593 993 13599
rect 9417 13567 9423 13593
rect 9449 13567 9455 13593
rect 12721 13567 12727 13593
rect 12753 13567 12759 13593
rect 967 13561 993 13567
rect 2025 13511 2031 13537
rect 2057 13511 2063 13537
rect 8017 13511 8023 13537
rect 8049 13511 8055 13537
rect 11265 13511 11271 13537
rect 11297 13511 11303 13537
rect 13001 13511 13007 13537
rect 13033 13511 13039 13537
rect 6847 13481 6873 13487
rect 10711 13481 10737 13487
rect 13287 13481 13313 13487
rect 8353 13455 8359 13481
rect 8385 13455 8391 13481
rect 11657 13455 11663 13481
rect 11689 13455 11695 13481
rect 12889 13455 12895 13481
rect 12921 13455 12927 13481
rect 6847 13449 6873 13455
rect 10711 13449 10737 13455
rect 13287 13449 13313 13455
rect 6903 13425 6929 13431
rect 6903 13393 6929 13399
rect 9647 13425 9673 13431
rect 9647 13393 9673 13399
rect 10655 13425 10681 13431
rect 10655 13393 10681 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 8415 13257 8441 13263
rect 12777 13231 12783 13257
rect 12809 13231 12815 13257
rect 8415 13225 8441 13231
rect 7065 13175 7071 13201
rect 7097 13175 7103 13201
rect 10089 13175 10095 13201
rect 10121 13175 10127 13201
rect 7687 13145 7713 13151
rect 9535 13145 9561 13151
rect 2137 13119 2143 13145
rect 2169 13119 2175 13145
rect 7457 13119 7463 13145
rect 7489 13119 7495 13145
rect 8297 13119 8303 13145
rect 8329 13119 8335 13145
rect 9697 13119 9703 13145
rect 9729 13119 9735 13145
rect 12665 13119 12671 13145
rect 12697 13119 12703 13145
rect 7687 13113 7713 13119
rect 9535 13113 9561 13119
rect 6001 13063 6007 13089
rect 6033 13063 6039 13089
rect 11153 13063 11159 13089
rect 11185 13063 11191 13089
rect 967 13033 993 13039
rect 967 13001 993 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 8303 12865 8329 12871
rect 8303 12833 8329 12839
rect 10823 12809 10849 12815
rect 10823 12777 10849 12783
rect 11495 12809 11521 12815
rect 11495 12777 11521 12783
rect 11663 12809 11689 12815
rect 20007 12809 20033 12815
rect 12105 12783 12111 12809
rect 12137 12783 12143 12809
rect 11663 12777 11689 12783
rect 20007 12777 20033 12783
rect 6903 12753 6929 12759
rect 6903 12721 6929 12727
rect 7015 12753 7041 12759
rect 7407 12753 7433 12759
rect 8135 12753 8161 12759
rect 9815 12753 9841 12759
rect 7233 12727 7239 12753
rect 7265 12727 7271 12753
rect 7569 12727 7575 12753
rect 7601 12727 7607 12753
rect 9585 12727 9591 12753
rect 9617 12727 9623 12753
rect 7015 12721 7041 12727
rect 7407 12721 7433 12727
rect 8135 12721 8161 12727
rect 9815 12721 9841 12727
rect 10767 12753 10793 12759
rect 10767 12721 10793 12727
rect 10879 12753 10905 12759
rect 10879 12721 10905 12727
rect 11607 12753 11633 12759
rect 12223 12753 12249 12759
rect 11713 12727 11719 12753
rect 11745 12727 11751 12753
rect 12329 12727 12335 12753
rect 12361 12727 12367 12753
rect 18825 12727 18831 12753
rect 18857 12727 18863 12753
rect 11607 12721 11633 12727
rect 12223 12721 12249 12727
rect 6343 12697 6369 12703
rect 6343 12665 6369 12671
rect 6791 12697 6817 12703
rect 6791 12665 6817 12671
rect 6847 12697 6873 12703
rect 6847 12665 6873 12671
rect 8023 12697 8049 12703
rect 8023 12665 8049 12671
rect 10655 12697 10681 12703
rect 10655 12665 10681 12671
rect 11439 12697 11465 12703
rect 11439 12665 11465 12671
rect 13455 12697 13481 12703
rect 13455 12665 13481 12671
rect 6399 12641 6425 12647
rect 6399 12609 6425 12615
rect 7351 12641 7377 12647
rect 7351 12609 7377 12615
rect 7463 12641 7489 12647
rect 10935 12641 10961 12647
rect 9473 12615 9479 12641
rect 9505 12615 9511 12641
rect 9977 12615 9983 12641
rect 10009 12615 10015 12641
rect 7463 12609 7489 12615
rect 10935 12609 10961 12615
rect 12055 12641 12081 12647
rect 12055 12609 12081 12615
rect 12111 12641 12137 12647
rect 12111 12609 12137 12615
rect 13511 12641 13537 12647
rect 13511 12609 13537 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 7239 12473 7265 12479
rect 10593 12447 10599 12473
rect 10625 12447 10631 12473
rect 7239 12441 7265 12447
rect 9815 12417 9841 12423
rect 6617 12391 6623 12417
rect 6649 12391 6655 12417
rect 9305 12391 9311 12417
rect 9337 12391 9343 12417
rect 9815 12385 9841 12391
rect 9871 12417 9897 12423
rect 9871 12385 9897 12391
rect 9927 12417 9953 12423
rect 13505 12391 13511 12417
rect 13537 12391 13543 12417
rect 9927 12385 9953 12391
rect 9479 12361 9505 12367
rect 12671 12361 12697 12367
rect 7009 12335 7015 12361
rect 7041 12335 7047 12361
rect 10481 12335 10487 12361
rect 10513 12335 10519 12361
rect 10929 12335 10935 12361
rect 10961 12335 10967 12361
rect 13113 12335 13119 12361
rect 13145 12335 13151 12361
rect 9479 12329 9505 12335
rect 12671 12329 12697 12335
rect 14799 12305 14825 12311
rect 5553 12279 5559 12305
rect 5585 12279 5591 12305
rect 11265 12279 11271 12305
rect 11297 12279 11303 12305
rect 12329 12279 12335 12305
rect 12361 12279 12367 12305
rect 14569 12279 14575 12305
rect 14601 12279 14607 12305
rect 14799 12273 14825 12279
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 9983 12081 10009 12087
rect 9983 12049 10009 12055
rect 967 12025 993 12031
rect 10039 12025 10065 12031
rect 9473 11999 9479 12025
rect 9505 11999 9511 12025
rect 967 11993 993 11999
rect 10039 11993 10065 11999
rect 10263 12025 10289 12031
rect 10263 11993 10289 11999
rect 11551 12025 11577 12031
rect 11551 11993 11577 11999
rect 13343 12025 13369 12031
rect 13343 11993 13369 11999
rect 9815 11969 9841 11975
rect 2137 11943 2143 11969
rect 2169 11943 2175 11969
rect 8073 11943 8079 11969
rect 8105 11943 8111 11969
rect 9815 11937 9841 11943
rect 11439 11969 11465 11975
rect 11439 11937 11465 11943
rect 11663 11969 11689 11975
rect 11663 11937 11689 11943
rect 11943 11969 11969 11975
rect 11943 11937 11969 11943
rect 13231 11969 13257 11975
rect 13231 11937 13257 11943
rect 13399 11969 13425 11975
rect 13399 11937 13425 11943
rect 6847 11913 6873 11919
rect 13287 11913 13313 11919
rect 8409 11887 8415 11913
rect 8441 11887 8447 11913
rect 11769 11887 11775 11913
rect 11801 11887 11807 11913
rect 6847 11881 6873 11887
rect 13287 11881 13313 11887
rect 6679 11857 6705 11863
rect 6679 11825 6705 11831
rect 6791 11857 6817 11863
rect 11495 11857 11521 11863
rect 9641 11831 9647 11857
rect 9673 11831 9679 11857
rect 6791 11825 6817 11831
rect 11495 11825 11521 11831
rect 13455 11857 13481 11863
rect 13455 11825 13481 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 7127 11689 7153 11695
rect 7127 11657 7153 11663
rect 7687 11689 7713 11695
rect 7687 11657 7713 11663
rect 6791 11633 6817 11639
rect 6791 11601 6817 11607
rect 6847 11633 6873 11639
rect 6847 11601 6873 11607
rect 7575 11633 7601 11639
rect 7575 11601 7601 11607
rect 11327 11633 11353 11639
rect 11327 11601 11353 11607
rect 15023 11633 15049 11639
rect 15023 11601 15049 11607
rect 7743 11577 7769 11583
rect 11383 11577 11409 11583
rect 2137 11551 2143 11577
rect 2169 11551 2175 11577
rect 6617 11551 6623 11577
rect 6649 11551 6655 11577
rect 7457 11551 7463 11577
rect 7489 11551 7495 11577
rect 9473 11551 9479 11577
rect 9505 11551 9511 11577
rect 9697 11551 9703 11577
rect 9729 11551 9735 11577
rect 7743 11545 7769 11551
rect 11383 11545 11409 11551
rect 11495 11577 11521 11583
rect 11495 11545 11521 11551
rect 11551 11577 11577 11583
rect 11713 11551 11719 11577
rect 11745 11551 11751 11577
rect 13337 11551 13343 11577
rect 13369 11551 13375 11577
rect 18825 11551 18831 11577
rect 18857 11551 18863 11577
rect 11551 11545 11577 11551
rect 7631 11521 7657 11527
rect 5161 11495 5167 11521
rect 5193 11495 5199 11521
rect 6225 11495 6231 11521
rect 6257 11495 6263 11521
rect 13729 11495 13735 11521
rect 13761 11495 13767 11521
rect 14793 11495 14799 11521
rect 14825 11495 14831 11521
rect 7631 11489 7657 11495
rect 967 11465 993 11471
rect 967 11433 993 11439
rect 6847 11465 6873 11471
rect 20007 11465 20033 11471
rect 9697 11439 9703 11465
rect 9729 11439 9735 11465
rect 6847 11433 6873 11439
rect 20007 11433 20033 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 7407 11297 7433 11303
rect 7407 11265 7433 11271
rect 7519 11297 7545 11303
rect 10039 11297 10065 11303
rect 9753 11271 9759 11297
rect 9785 11271 9791 11297
rect 7519 11265 7545 11271
rect 10039 11265 10065 11271
rect 12111 11297 12137 11303
rect 12111 11265 12137 11271
rect 967 11241 993 11247
rect 967 11209 993 11215
rect 9927 11241 9953 11247
rect 13567 11241 13593 11247
rect 12273 11215 12279 11241
rect 12305 11215 12311 11241
rect 9927 11209 9953 11215
rect 13567 11209 13593 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 7575 11185 7601 11191
rect 2137 11159 2143 11185
rect 2169 11159 2175 11185
rect 7575 11153 7601 11159
rect 7799 11185 7825 11191
rect 7799 11153 7825 11159
rect 7967 11185 7993 11191
rect 9199 11185 9225 11191
rect 8913 11159 8919 11185
rect 8945 11159 8951 11185
rect 7967 11153 7993 11159
rect 9199 11153 9225 11159
rect 9479 11185 9505 11191
rect 9479 11153 9505 11159
rect 11215 11185 11241 11191
rect 11215 11153 11241 11159
rect 11383 11185 11409 11191
rect 11383 11153 11409 11159
rect 11439 11185 11465 11191
rect 13847 11185 13873 11191
rect 11489 11159 11495 11185
rect 11521 11159 11527 11185
rect 11439 11153 11465 11159
rect 13847 11153 13873 11159
rect 14015 11185 14041 11191
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 14015 11153 14041 11159
rect 7351 11129 7377 11135
rect 7351 11097 7377 11103
rect 8751 11129 8777 11135
rect 8751 11097 8777 11103
rect 9143 11129 9169 11135
rect 9143 11097 9169 11103
rect 9423 11129 9449 11135
rect 9423 11097 9449 11103
rect 9535 11129 9561 11135
rect 12223 11129 12249 11135
rect 11937 11103 11943 11129
rect 11969 11103 11975 11129
rect 9535 11097 9561 11103
rect 12223 11097 12249 11103
rect 14127 11129 14153 11135
rect 14127 11097 14153 11103
rect 14183 11129 14209 11135
rect 14183 11097 14209 11103
rect 7911 11073 7937 11079
rect 7911 11041 7937 11047
rect 8807 11073 8833 11079
rect 8807 11041 8833 11047
rect 9031 11073 9057 11079
rect 11607 11073 11633 11079
rect 10201 11047 10207 11073
rect 10233 11047 10239 11073
rect 9031 11041 9057 11047
rect 11607 11041 11633 11047
rect 11775 11073 11801 11079
rect 11775 11041 11801 11047
rect 13511 11073 13537 11079
rect 13511 11041 13537 11047
rect 13623 11073 13649 11079
rect 13623 11041 13649 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 7631 10905 7657 10911
rect 7631 10873 7657 10879
rect 8863 10905 8889 10911
rect 11047 10905 11073 10911
rect 10425 10879 10431 10905
rect 10457 10879 10463 10905
rect 11433 10879 11439 10905
rect 11465 10879 11471 10905
rect 8863 10873 8889 10879
rect 11047 10873 11073 10879
rect 9591 10849 9617 10855
rect 8689 10823 8695 10849
rect 8721 10823 8727 10849
rect 9081 10823 9087 10849
rect 9113 10823 9119 10849
rect 9591 10817 9617 10823
rect 10879 10849 10905 10855
rect 11881 10823 11887 10849
rect 11913 10823 11919 10849
rect 13169 10823 13175 10849
rect 13201 10823 13207 10849
rect 10879 10817 10905 10823
rect 10039 10793 10065 10799
rect 2137 10767 2143 10793
rect 2169 10767 2175 10793
rect 7009 10767 7015 10793
rect 7041 10767 7047 10793
rect 7401 10767 7407 10793
rect 7433 10767 7439 10793
rect 9193 10767 9199 10793
rect 9225 10767 9231 10793
rect 10039 10761 10065 10767
rect 10095 10793 10121 10799
rect 10095 10761 10121 10767
rect 10263 10793 10289 10799
rect 10263 10761 10289 10767
rect 10599 10793 10625 10799
rect 10599 10761 10625 10767
rect 10991 10793 11017 10799
rect 10991 10761 11017 10767
rect 11103 10793 11129 10799
rect 11103 10761 11129 10767
rect 11271 10793 11297 10799
rect 11769 10767 11775 10793
rect 11801 10767 11807 10793
rect 13057 10767 13063 10793
rect 13089 10767 13095 10793
rect 13393 10767 13399 10793
rect 13425 10767 13431 10793
rect 11271 10761 11297 10767
rect 10207 10737 10233 10743
rect 15079 10737 15105 10743
rect 5945 10711 5951 10737
rect 5977 10711 5983 10737
rect 13785 10711 13791 10737
rect 13817 10711 13823 10737
rect 14849 10711 14855 10737
rect 14881 10711 14887 10737
rect 10207 10705 10233 10711
rect 15079 10705 15105 10711
rect 967 10681 993 10687
rect 967 10649 993 10655
rect 9535 10681 9561 10687
rect 9535 10649 9561 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 6903 10513 6929 10519
rect 6903 10481 6929 10487
rect 7015 10513 7041 10519
rect 7015 10481 7041 10487
rect 10711 10457 10737 10463
rect 10711 10425 10737 10431
rect 11439 10457 11465 10463
rect 14631 10457 14657 10463
rect 13393 10431 13399 10457
rect 13425 10431 13431 10457
rect 11439 10425 11465 10431
rect 14631 10425 14657 10431
rect 7407 10401 7433 10407
rect 10767 10401 10793 10407
rect 14575 10401 14601 10407
rect 7121 10375 7127 10401
rect 7153 10375 7159 10401
rect 10033 10375 10039 10401
rect 10065 10375 10071 10401
rect 11657 10375 11663 10401
rect 11689 10375 11695 10401
rect 7407 10369 7433 10375
rect 10767 10369 10793 10375
rect 14575 10369 14601 10375
rect 14687 10401 14713 10407
rect 14687 10369 14713 10375
rect 6847 10345 6873 10351
rect 6847 10313 6873 10319
rect 7295 10345 7321 10351
rect 7295 10313 7321 10319
rect 7575 10345 7601 10351
rect 10655 10345 10681 10351
rect 7849 10319 7855 10345
rect 7881 10319 7887 10345
rect 7575 10313 7601 10319
rect 10655 10313 10681 10319
rect 10935 10345 10961 10351
rect 10935 10313 10961 10319
rect 11159 10345 11185 10351
rect 11159 10313 11185 10319
rect 11495 10345 11521 10351
rect 11495 10313 11521 10319
rect 7463 10289 7489 10295
rect 7463 10257 7489 10263
rect 11103 10289 11129 10295
rect 11103 10257 11129 10263
rect 11383 10289 11409 10295
rect 11383 10257 11409 10263
rect 14799 10289 14825 10295
rect 14799 10257 14825 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 7855 10121 7881 10127
rect 7855 10089 7881 10095
rect 8863 10121 8889 10127
rect 8863 10089 8889 10095
rect 14295 10121 14321 10127
rect 14295 10089 14321 10095
rect 14575 10121 14601 10127
rect 14575 10089 14601 10095
rect 7631 10065 7657 10071
rect 6897 10039 6903 10065
rect 6929 10039 6935 10065
rect 7457 10039 7463 10065
rect 7489 10039 7495 10065
rect 7631 10033 7657 10039
rect 9423 10065 9449 10071
rect 9423 10033 9449 10039
rect 9479 10065 9505 10071
rect 14239 10065 14265 10071
rect 11657 10039 11663 10065
rect 11689 10039 11695 10065
rect 9479 10033 9505 10039
rect 14239 10033 14265 10039
rect 8807 10009 8833 10015
rect 2137 9983 2143 10009
rect 2169 9983 2175 10009
rect 7289 9983 7295 10009
rect 7321 9983 7327 10009
rect 8807 9977 8833 9983
rect 8975 10009 9001 10015
rect 14407 10009 14433 10015
rect 9081 9983 9087 10009
rect 9113 9983 9119 10009
rect 9697 9983 9703 10009
rect 9729 9983 9735 10009
rect 12665 9983 12671 10009
rect 12697 9983 12703 10009
rect 18825 9983 18831 10009
rect 18857 9983 18863 10009
rect 8975 9977 9001 9983
rect 14407 9977 14433 9983
rect 8919 9953 8945 9959
rect 5833 9927 5839 9953
rect 5865 9927 5871 9953
rect 13001 9927 13007 9953
rect 13033 9927 13039 9953
rect 14065 9927 14071 9953
rect 14097 9927 14103 9953
rect 8919 9921 8945 9927
rect 967 9897 993 9903
rect 967 9865 993 9871
rect 9535 9897 9561 9903
rect 9535 9865 9561 9871
rect 20007 9897 20033 9903
rect 20007 9865 20033 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 9983 9673 10009 9679
rect 7737 9647 7743 9673
rect 7769 9647 7775 9673
rect 9983 9641 10009 9647
rect 12279 9673 12305 9679
rect 12279 9641 12305 9647
rect 7183 9617 7209 9623
rect 9703 9617 9729 9623
rect 10935 9617 10961 9623
rect 9137 9591 9143 9617
rect 9169 9591 9175 9617
rect 9865 9591 9871 9617
rect 9897 9591 9903 9617
rect 7183 9585 7209 9591
rect 9703 9585 9729 9591
rect 10935 9585 10961 9591
rect 11159 9617 11185 9623
rect 11159 9585 11185 9591
rect 11495 9617 11521 9623
rect 11495 9585 11521 9591
rect 12223 9617 12249 9623
rect 12223 9585 12249 9591
rect 12335 9617 12361 9623
rect 12335 9585 12361 9591
rect 13063 9617 13089 9623
rect 13337 9591 13343 9617
rect 13369 9591 13375 9617
rect 13063 9585 13089 9591
rect 6735 9561 6761 9567
rect 10039 9561 10065 9567
rect 8801 9535 8807 9561
rect 8833 9535 8839 9561
rect 9529 9535 9535 9561
rect 9561 9535 9567 9561
rect 6735 9529 6761 9535
rect 10039 9529 10065 9535
rect 11663 9561 11689 9567
rect 11663 9529 11689 9535
rect 12055 9561 12081 9567
rect 12055 9529 12081 9535
rect 13119 9561 13145 9567
rect 13119 9529 13145 9535
rect 6791 9505 6817 9511
rect 6791 9473 6817 9479
rect 6903 9505 6929 9511
rect 10375 9505 10401 9511
rect 7009 9479 7015 9505
rect 7041 9479 7047 9505
rect 10201 9479 10207 9505
rect 10233 9479 10239 9505
rect 6903 9473 6929 9479
rect 10375 9473 10401 9479
rect 10711 9505 10737 9511
rect 10711 9473 10737 9479
rect 10823 9505 10849 9511
rect 10823 9473 10849 9479
rect 10879 9505 10905 9511
rect 13175 9505 13201 9511
rect 11321 9479 11327 9505
rect 11353 9479 11359 9505
rect 10879 9473 10905 9479
rect 13175 9473 13201 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 8807 9337 8833 9343
rect 8807 9305 8833 9311
rect 9591 9337 9617 9343
rect 9591 9305 9617 9311
rect 13623 9337 13649 9343
rect 13623 9305 13649 9311
rect 7183 9281 7209 9287
rect 7183 9249 7209 9255
rect 7463 9281 7489 9287
rect 7463 9249 7489 9255
rect 7687 9281 7713 9287
rect 7687 9249 7713 9255
rect 8863 9281 8889 9287
rect 8863 9249 8889 9255
rect 11775 9281 11801 9287
rect 11775 9249 11801 9255
rect 13567 9281 13593 9287
rect 13567 9249 13593 9255
rect 7295 9225 7321 9231
rect 9311 9225 9337 9231
rect 12111 9225 12137 9231
rect 2137 9199 2143 9225
rect 2169 9199 2175 9225
rect 6449 9199 6455 9225
rect 6481 9199 6487 9225
rect 6785 9199 6791 9225
rect 6817 9199 6823 9225
rect 8689 9199 8695 9225
rect 8721 9199 8727 9225
rect 11153 9199 11159 9225
rect 11185 9199 11191 9225
rect 11545 9199 11551 9225
rect 11577 9199 11583 9225
rect 7295 9193 7321 9199
rect 9311 9193 9337 9199
rect 12111 9193 12137 9199
rect 13735 9225 13761 9231
rect 13735 9193 13761 9199
rect 7239 9169 7265 9175
rect 5385 9143 5391 9169
rect 5417 9143 5423 9169
rect 10089 9143 10095 9169
rect 10121 9143 10127 9169
rect 11713 9143 11719 9169
rect 11745 9143 11751 9169
rect 7239 9137 7265 9143
rect 967 9113 993 9119
rect 967 9081 993 9087
rect 11887 9113 11913 9119
rect 11887 9081 11913 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 6791 8945 6817 8951
rect 6791 8913 6817 8919
rect 7239 8945 7265 8951
rect 7239 8913 7265 8919
rect 9759 8945 9785 8951
rect 9759 8913 9785 8919
rect 13903 8945 13929 8951
rect 13903 8913 13929 8919
rect 967 8889 993 8895
rect 13287 8889 13313 8895
rect 7065 8863 7071 8889
rect 7097 8863 7103 8889
rect 967 8857 993 8863
rect 13287 8857 13313 8863
rect 20007 8889 20033 8895
rect 20007 8857 20033 8863
rect 6847 8833 6873 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 6847 8801 6873 8807
rect 8583 8833 8609 8839
rect 13231 8833 13257 8839
rect 9641 8807 9647 8833
rect 9673 8807 9679 8833
rect 10201 8807 10207 8833
rect 10233 8807 10239 8833
rect 10313 8807 10319 8833
rect 10345 8807 10351 8833
rect 11209 8807 11215 8833
rect 11241 8807 11247 8833
rect 8583 8801 8609 8807
rect 13231 8801 13257 8807
rect 13343 8833 13369 8839
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 13343 8801 13369 8807
rect 6791 8777 6817 8783
rect 13847 8777 13873 8783
rect 10929 8751 10935 8777
rect 10961 8751 10967 8777
rect 11097 8751 11103 8777
rect 11129 8751 11135 8777
rect 12889 8751 12895 8777
rect 12921 8751 12927 8777
rect 6791 8745 6817 8751
rect 13847 8745 13873 8751
rect 13903 8777 13929 8783
rect 13903 8745 13929 8751
rect 7127 8721 7153 8727
rect 7127 8689 7153 8695
rect 8639 8721 8665 8727
rect 8639 8689 8665 8695
rect 8751 8721 8777 8727
rect 12727 8721 12753 8727
rect 10761 8695 10767 8721
rect 10793 8695 10799 8721
rect 8751 8689 8777 8695
rect 12727 8689 12753 8695
rect 13119 8721 13145 8727
rect 13119 8689 13145 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 7575 8553 7601 8559
rect 7575 8521 7601 8527
rect 8303 8553 8329 8559
rect 8303 8521 8329 8527
rect 8919 8553 8945 8559
rect 8919 8521 8945 8527
rect 9087 8553 9113 8559
rect 9087 8521 9113 8527
rect 10655 8553 10681 8559
rect 10655 8521 10681 8527
rect 11215 8553 11241 8559
rect 15023 8553 15049 8559
rect 11377 8527 11383 8553
rect 11409 8527 11415 8553
rect 11215 8521 11241 8527
rect 15023 8521 15049 8527
rect 8807 8497 8833 8503
rect 6953 8471 6959 8497
rect 6985 8471 6991 8497
rect 8807 8465 8833 8471
rect 12839 8497 12865 8503
rect 13729 8471 13735 8497
rect 13761 8471 13767 8497
rect 12839 8465 12865 8471
rect 9031 8441 9057 8447
rect 12951 8441 12977 8447
rect 7345 8415 7351 8441
rect 7377 8415 7383 8441
rect 10145 8415 10151 8441
rect 10177 8415 10183 8441
rect 13393 8415 13399 8441
rect 13425 8415 13431 8441
rect 9031 8409 9057 8415
rect 12951 8409 12977 8415
rect 8975 8385 9001 8391
rect 5889 8359 5895 8385
rect 5921 8359 5927 8385
rect 8975 8353 9001 8359
rect 9983 8385 10009 8391
rect 10543 8385 10569 8391
rect 10089 8359 10095 8385
rect 10121 8359 10127 8385
rect 9983 8353 10009 8359
rect 10543 8353 10569 8359
rect 10599 8385 10625 8391
rect 14793 8359 14799 8385
rect 14825 8359 14831 8385
rect 10599 8353 10625 8359
rect 8247 8329 8273 8335
rect 8247 8297 8273 8303
rect 8415 8329 8441 8335
rect 8415 8297 8441 8303
rect 13119 8329 13145 8335
rect 13119 8297 13145 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 10767 8161 10793 8167
rect 10767 8129 10793 8135
rect 10879 8161 10905 8167
rect 10879 8129 10905 8135
rect 9255 8105 9281 8111
rect 7961 8079 7967 8105
rect 7993 8079 7999 8105
rect 9025 8079 9031 8105
rect 9057 8079 9063 8105
rect 9255 8073 9281 8079
rect 20007 8105 20033 8111
rect 20007 8073 20033 8079
rect 13679 8049 13705 8055
rect 7569 8023 7575 8049
rect 7601 8023 7607 8049
rect 10649 8023 10655 8049
rect 10681 8023 10687 8049
rect 12497 8023 12503 8049
rect 12529 8023 12535 8049
rect 12833 8023 12839 8049
rect 12865 8023 12871 8049
rect 18825 8023 18831 8049
rect 18857 8023 18863 8049
rect 13679 8017 13705 8023
rect 10935 7993 10961 7999
rect 13175 7993 13201 7999
rect 11153 7967 11159 7993
rect 11185 7967 11191 7993
rect 13225 7967 13231 7993
rect 13257 7967 13263 7993
rect 10935 7961 10961 7967
rect 13175 7961 13201 7967
rect 11327 7937 11353 7943
rect 11327 7905 11353 7911
rect 12615 7937 12641 7943
rect 12615 7905 12641 7911
rect 12671 7937 12697 7943
rect 12671 7905 12697 7911
rect 12727 7937 12753 7943
rect 12727 7905 12753 7911
rect 13007 7937 13033 7943
rect 13007 7905 13033 7911
rect 13063 7937 13089 7943
rect 13063 7905 13089 7911
rect 13119 7937 13145 7943
rect 13119 7905 13145 7911
rect 13511 7937 13537 7943
rect 13511 7905 13537 7911
rect 13623 7937 13649 7943
rect 13623 7905 13649 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 10207 7769 10233 7775
rect 11607 7769 11633 7775
rect 14407 7769 14433 7775
rect 11265 7743 11271 7769
rect 11297 7743 11303 7769
rect 11769 7743 11775 7769
rect 11801 7743 11807 7769
rect 10207 7737 10233 7743
rect 11607 7737 11633 7743
rect 14407 7737 14433 7743
rect 8695 7713 8721 7719
rect 8695 7681 8721 7687
rect 8807 7713 8833 7719
rect 8807 7681 8833 7687
rect 9087 7713 9113 7719
rect 9087 7681 9113 7687
rect 9199 7713 9225 7719
rect 9199 7681 9225 7687
rect 9255 7713 9281 7719
rect 9255 7681 9281 7687
rect 12279 7713 12305 7719
rect 12279 7681 12305 7687
rect 8919 7657 8945 7663
rect 8919 7625 8945 7631
rect 9031 7657 9057 7663
rect 10095 7657 10121 7663
rect 9921 7631 9927 7657
rect 9953 7631 9959 7657
rect 9031 7625 9057 7631
rect 10095 7625 10121 7631
rect 11047 7657 11073 7663
rect 11047 7625 11073 7631
rect 11439 7657 11465 7663
rect 12777 7631 12783 7657
rect 12809 7631 12815 7657
rect 13113 7631 13119 7657
rect 13145 7631 13151 7657
rect 18825 7631 18831 7657
rect 18857 7631 18863 7657
rect 11439 7625 11465 7631
rect 10151 7601 10177 7607
rect 10151 7569 10177 7575
rect 11103 7601 11129 7607
rect 20007 7601 20033 7607
rect 14177 7575 14183 7601
rect 14209 7575 14215 7601
rect 11103 7569 11129 7575
rect 20007 7569 20033 7575
rect 12335 7545 12361 7551
rect 12335 7513 12361 7519
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 9815 7377 9841 7383
rect 9815 7345 9841 7351
rect 8975 7321 9001 7327
rect 14015 7321 14041 7327
rect 7681 7295 7687 7321
rect 7713 7295 7719 7321
rect 8745 7295 8751 7321
rect 8777 7295 8783 7321
rect 9641 7295 9647 7321
rect 9673 7295 9679 7321
rect 11041 7295 11047 7321
rect 11073 7295 11079 7321
rect 12105 7295 12111 7321
rect 12137 7295 12143 7321
rect 12721 7295 12727 7321
rect 12753 7295 12759 7321
rect 13785 7295 13791 7321
rect 13817 7295 13823 7321
rect 8975 7289 9001 7295
rect 14015 7289 14041 7295
rect 7345 7239 7351 7265
rect 7377 7239 7383 7265
rect 10705 7239 10711 7265
rect 10737 7239 10743 7265
rect 12329 7239 12335 7265
rect 12361 7239 12367 7265
rect 9703 7209 9729 7215
rect 9703 7177 9729 7183
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 12279 6985 12305 6991
rect 12279 6953 12305 6959
rect 9305 6903 9311 6929
rect 9337 6903 9343 6929
rect 8751 6873 8777 6879
rect 8969 6847 8975 6873
rect 9001 6847 9007 6873
rect 8751 6841 8777 6847
rect 10369 6791 10375 6817
rect 10401 6791 10407 6817
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 8857 2143 8863 2169
rect 8889 2143 8895 2169
rect 9367 2057 9393 2063
rect 9367 2025 9393 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 9311 1833 9337 1839
rect 9311 1801 9337 1807
rect 8969 1751 8975 1777
rect 9001 1751 9007 1777
rect 10369 1751 10375 1777
rect 10401 1751 10407 1777
rect 10879 1665 10905 1671
rect 10879 1633 10905 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 11215 19111 11241 19137
rect 14687 19111 14713 19137
rect 12839 19055 12865 19081
rect 10879 18999 10905 19025
rect 12279 18999 12305 19025
rect 14295 18999 14321 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 12223 18719 12249 18745
rect 13119 18719 13145 18745
rect 12839 18607 12865 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 11999 18327 12025 18353
rect 12951 18215 12977 18241
rect 20119 18103 20145 18129
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 967 13567 993 13593
rect 9423 13567 9449 13593
rect 12727 13567 12753 13593
rect 2031 13511 2057 13537
rect 8023 13511 8049 13537
rect 11271 13511 11297 13537
rect 13007 13511 13033 13537
rect 6847 13455 6873 13481
rect 8359 13455 8385 13481
rect 10711 13455 10737 13481
rect 11663 13455 11689 13481
rect 12895 13455 12921 13481
rect 13287 13455 13313 13481
rect 6903 13399 6929 13425
rect 9647 13399 9673 13425
rect 10655 13399 10681 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 8415 13231 8441 13257
rect 12783 13231 12809 13257
rect 7071 13175 7097 13201
rect 10095 13175 10121 13201
rect 2143 13119 2169 13145
rect 7463 13119 7489 13145
rect 7687 13119 7713 13145
rect 8303 13119 8329 13145
rect 9535 13119 9561 13145
rect 9703 13119 9729 13145
rect 12671 13119 12697 13145
rect 6007 13063 6033 13089
rect 11159 13063 11185 13089
rect 967 13007 993 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 8303 12839 8329 12865
rect 10823 12783 10849 12809
rect 11495 12783 11521 12809
rect 11663 12783 11689 12809
rect 12111 12783 12137 12809
rect 20007 12783 20033 12809
rect 6903 12727 6929 12753
rect 7015 12727 7041 12753
rect 7239 12727 7265 12753
rect 7407 12727 7433 12753
rect 7575 12727 7601 12753
rect 8135 12727 8161 12753
rect 9591 12727 9617 12753
rect 9815 12727 9841 12753
rect 10767 12727 10793 12753
rect 10879 12727 10905 12753
rect 11607 12727 11633 12753
rect 11719 12727 11745 12753
rect 12223 12727 12249 12753
rect 12335 12727 12361 12753
rect 18831 12727 18857 12753
rect 6343 12671 6369 12697
rect 6791 12671 6817 12697
rect 6847 12671 6873 12697
rect 8023 12671 8049 12697
rect 10655 12671 10681 12697
rect 11439 12671 11465 12697
rect 13455 12671 13481 12697
rect 6399 12615 6425 12641
rect 7351 12615 7377 12641
rect 7463 12615 7489 12641
rect 9479 12615 9505 12641
rect 9983 12615 10009 12641
rect 10935 12615 10961 12641
rect 12055 12615 12081 12641
rect 12111 12615 12137 12641
rect 13511 12615 13537 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 7239 12447 7265 12473
rect 10599 12447 10625 12473
rect 6623 12391 6649 12417
rect 9311 12391 9337 12417
rect 9815 12391 9841 12417
rect 9871 12391 9897 12417
rect 9927 12391 9953 12417
rect 13511 12391 13537 12417
rect 7015 12335 7041 12361
rect 9479 12335 9505 12361
rect 10487 12335 10513 12361
rect 10935 12335 10961 12361
rect 12671 12335 12697 12361
rect 13119 12335 13145 12361
rect 5559 12279 5585 12305
rect 11271 12279 11297 12305
rect 12335 12279 12361 12305
rect 14575 12279 14601 12305
rect 14799 12279 14825 12305
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 9983 12055 10009 12081
rect 967 11999 993 12025
rect 9479 11999 9505 12025
rect 10039 11999 10065 12025
rect 10263 11999 10289 12025
rect 11551 11999 11577 12025
rect 13343 11999 13369 12025
rect 2143 11943 2169 11969
rect 8079 11943 8105 11969
rect 9815 11943 9841 11969
rect 11439 11943 11465 11969
rect 11663 11943 11689 11969
rect 11943 11943 11969 11969
rect 13231 11943 13257 11969
rect 13399 11943 13425 11969
rect 6847 11887 6873 11913
rect 8415 11887 8441 11913
rect 11775 11887 11801 11913
rect 13287 11887 13313 11913
rect 6679 11831 6705 11857
rect 6791 11831 6817 11857
rect 9647 11831 9673 11857
rect 11495 11831 11521 11857
rect 13455 11831 13481 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 7127 11663 7153 11689
rect 7687 11663 7713 11689
rect 6791 11607 6817 11633
rect 6847 11607 6873 11633
rect 7575 11607 7601 11633
rect 11327 11607 11353 11633
rect 15023 11607 15049 11633
rect 2143 11551 2169 11577
rect 6623 11551 6649 11577
rect 7463 11551 7489 11577
rect 7743 11551 7769 11577
rect 9479 11551 9505 11577
rect 9703 11551 9729 11577
rect 11383 11551 11409 11577
rect 11495 11551 11521 11577
rect 11551 11551 11577 11577
rect 11719 11551 11745 11577
rect 13343 11551 13369 11577
rect 18831 11551 18857 11577
rect 5167 11495 5193 11521
rect 6231 11495 6257 11521
rect 7631 11495 7657 11521
rect 13735 11495 13761 11521
rect 14799 11495 14825 11521
rect 967 11439 993 11465
rect 6847 11439 6873 11465
rect 9703 11439 9729 11465
rect 20007 11439 20033 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 7407 11271 7433 11297
rect 7519 11271 7545 11297
rect 9759 11271 9785 11297
rect 10039 11271 10065 11297
rect 12111 11271 12137 11297
rect 967 11215 993 11241
rect 9927 11215 9953 11241
rect 12279 11215 12305 11241
rect 13567 11215 13593 11241
rect 20007 11215 20033 11241
rect 2143 11159 2169 11185
rect 7575 11159 7601 11185
rect 7799 11159 7825 11185
rect 7967 11159 7993 11185
rect 8919 11159 8945 11185
rect 9199 11159 9225 11185
rect 9479 11159 9505 11185
rect 11215 11159 11241 11185
rect 11383 11159 11409 11185
rect 11439 11159 11465 11185
rect 11495 11159 11521 11185
rect 13847 11159 13873 11185
rect 14015 11159 14041 11185
rect 18831 11159 18857 11185
rect 7351 11103 7377 11129
rect 8751 11103 8777 11129
rect 9143 11103 9169 11129
rect 9423 11103 9449 11129
rect 9535 11103 9561 11129
rect 11943 11103 11969 11129
rect 12223 11103 12249 11129
rect 14127 11103 14153 11129
rect 14183 11103 14209 11129
rect 7911 11047 7937 11073
rect 8807 11047 8833 11073
rect 9031 11047 9057 11073
rect 10207 11047 10233 11073
rect 11607 11047 11633 11073
rect 11775 11047 11801 11073
rect 13511 11047 13537 11073
rect 13623 11047 13649 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 7631 10879 7657 10905
rect 8863 10879 8889 10905
rect 10431 10879 10457 10905
rect 11047 10879 11073 10905
rect 11439 10879 11465 10905
rect 8695 10823 8721 10849
rect 9087 10823 9113 10849
rect 9591 10823 9617 10849
rect 10879 10823 10905 10849
rect 11887 10823 11913 10849
rect 13175 10823 13201 10849
rect 2143 10767 2169 10793
rect 7015 10767 7041 10793
rect 7407 10767 7433 10793
rect 9199 10767 9225 10793
rect 10039 10767 10065 10793
rect 10095 10767 10121 10793
rect 10263 10767 10289 10793
rect 10599 10767 10625 10793
rect 10991 10767 11017 10793
rect 11103 10767 11129 10793
rect 11271 10767 11297 10793
rect 11775 10767 11801 10793
rect 13063 10767 13089 10793
rect 13399 10767 13425 10793
rect 5951 10711 5977 10737
rect 10207 10711 10233 10737
rect 13791 10711 13817 10737
rect 14855 10711 14881 10737
rect 15079 10711 15105 10737
rect 967 10655 993 10681
rect 9535 10655 9561 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 6903 10487 6929 10513
rect 7015 10487 7041 10513
rect 10711 10431 10737 10457
rect 11439 10431 11465 10457
rect 13399 10431 13425 10457
rect 14631 10431 14657 10457
rect 7127 10375 7153 10401
rect 7407 10375 7433 10401
rect 10039 10375 10065 10401
rect 10767 10375 10793 10401
rect 11663 10375 11689 10401
rect 14575 10375 14601 10401
rect 14687 10375 14713 10401
rect 6847 10319 6873 10345
rect 7295 10319 7321 10345
rect 7575 10319 7601 10345
rect 7855 10319 7881 10345
rect 10655 10319 10681 10345
rect 10935 10319 10961 10345
rect 11159 10319 11185 10345
rect 11495 10319 11521 10345
rect 7463 10263 7489 10289
rect 11103 10263 11129 10289
rect 11383 10263 11409 10289
rect 14799 10263 14825 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 7855 10095 7881 10121
rect 8863 10095 8889 10121
rect 14295 10095 14321 10121
rect 14575 10095 14601 10121
rect 6903 10039 6929 10065
rect 7463 10039 7489 10065
rect 7631 10039 7657 10065
rect 9423 10039 9449 10065
rect 9479 10039 9505 10065
rect 11663 10039 11689 10065
rect 14239 10039 14265 10065
rect 2143 9983 2169 10009
rect 7295 9983 7321 10009
rect 8807 9983 8833 10009
rect 8975 9983 9001 10009
rect 9087 9983 9113 10009
rect 9703 9983 9729 10009
rect 12671 9983 12697 10009
rect 14407 9983 14433 10009
rect 18831 9983 18857 10009
rect 5839 9927 5865 9953
rect 8919 9927 8945 9953
rect 13007 9927 13033 9953
rect 14071 9927 14097 9953
rect 967 9871 993 9897
rect 9535 9871 9561 9897
rect 20007 9871 20033 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 7743 9647 7769 9673
rect 9983 9647 10009 9673
rect 12279 9647 12305 9673
rect 7183 9591 7209 9617
rect 9143 9591 9169 9617
rect 9703 9591 9729 9617
rect 9871 9591 9897 9617
rect 10935 9591 10961 9617
rect 11159 9591 11185 9617
rect 11495 9591 11521 9617
rect 12223 9591 12249 9617
rect 12335 9591 12361 9617
rect 13063 9591 13089 9617
rect 13343 9591 13369 9617
rect 6735 9535 6761 9561
rect 8807 9535 8833 9561
rect 9535 9535 9561 9561
rect 10039 9535 10065 9561
rect 11663 9535 11689 9561
rect 12055 9535 12081 9561
rect 13119 9535 13145 9561
rect 6791 9479 6817 9505
rect 6903 9479 6929 9505
rect 7015 9479 7041 9505
rect 10207 9479 10233 9505
rect 10375 9479 10401 9505
rect 10711 9479 10737 9505
rect 10823 9479 10849 9505
rect 10879 9479 10905 9505
rect 11327 9479 11353 9505
rect 13175 9479 13201 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 8807 9311 8833 9337
rect 9591 9311 9617 9337
rect 13623 9311 13649 9337
rect 7183 9255 7209 9281
rect 7463 9255 7489 9281
rect 7687 9255 7713 9281
rect 8863 9255 8889 9281
rect 11775 9255 11801 9281
rect 13567 9255 13593 9281
rect 2143 9199 2169 9225
rect 6455 9199 6481 9225
rect 6791 9199 6817 9225
rect 7295 9199 7321 9225
rect 8695 9199 8721 9225
rect 9311 9199 9337 9225
rect 11159 9199 11185 9225
rect 11551 9199 11577 9225
rect 12111 9199 12137 9225
rect 13735 9199 13761 9225
rect 5391 9143 5417 9169
rect 7239 9143 7265 9169
rect 10095 9143 10121 9169
rect 11719 9143 11745 9169
rect 967 9087 993 9113
rect 11887 9087 11913 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 6791 8919 6817 8945
rect 7239 8919 7265 8945
rect 9759 8919 9785 8945
rect 13903 8919 13929 8945
rect 967 8863 993 8889
rect 7071 8863 7097 8889
rect 13287 8863 13313 8889
rect 20007 8863 20033 8889
rect 2143 8807 2169 8833
rect 6847 8807 6873 8833
rect 8583 8807 8609 8833
rect 9647 8807 9673 8833
rect 10207 8807 10233 8833
rect 10319 8807 10345 8833
rect 11215 8807 11241 8833
rect 13231 8807 13257 8833
rect 13343 8807 13369 8833
rect 18831 8807 18857 8833
rect 6791 8751 6817 8777
rect 10935 8751 10961 8777
rect 11103 8751 11129 8777
rect 12895 8751 12921 8777
rect 13847 8751 13873 8777
rect 13903 8751 13929 8777
rect 7127 8695 7153 8721
rect 8639 8695 8665 8721
rect 8751 8695 8777 8721
rect 10767 8695 10793 8721
rect 12727 8695 12753 8721
rect 13119 8695 13145 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7575 8527 7601 8553
rect 8303 8527 8329 8553
rect 8919 8527 8945 8553
rect 9087 8527 9113 8553
rect 10655 8527 10681 8553
rect 11215 8527 11241 8553
rect 11383 8527 11409 8553
rect 15023 8527 15049 8553
rect 6959 8471 6985 8497
rect 8807 8471 8833 8497
rect 12839 8471 12865 8497
rect 13735 8471 13761 8497
rect 7351 8415 7377 8441
rect 9031 8415 9057 8441
rect 10151 8415 10177 8441
rect 12951 8415 12977 8441
rect 13399 8415 13425 8441
rect 5895 8359 5921 8385
rect 8975 8359 9001 8385
rect 9983 8359 10009 8385
rect 10095 8359 10121 8385
rect 10543 8359 10569 8385
rect 10599 8359 10625 8385
rect 14799 8359 14825 8385
rect 8247 8303 8273 8329
rect 8415 8303 8441 8329
rect 13119 8303 13145 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 10767 8135 10793 8161
rect 10879 8135 10905 8161
rect 7967 8079 7993 8105
rect 9031 8079 9057 8105
rect 9255 8079 9281 8105
rect 20007 8079 20033 8105
rect 7575 8023 7601 8049
rect 10655 8023 10681 8049
rect 12503 8023 12529 8049
rect 12839 8023 12865 8049
rect 13679 8023 13705 8049
rect 18831 8023 18857 8049
rect 10935 7967 10961 7993
rect 11159 7967 11185 7993
rect 13175 7967 13201 7993
rect 13231 7967 13257 7993
rect 11327 7911 11353 7937
rect 12615 7911 12641 7937
rect 12671 7911 12697 7937
rect 12727 7911 12753 7937
rect 13007 7911 13033 7937
rect 13063 7911 13089 7937
rect 13119 7911 13145 7937
rect 13511 7911 13537 7937
rect 13623 7911 13649 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 10207 7743 10233 7769
rect 11271 7743 11297 7769
rect 11607 7743 11633 7769
rect 11775 7743 11801 7769
rect 14407 7743 14433 7769
rect 8695 7687 8721 7713
rect 8807 7687 8833 7713
rect 9087 7687 9113 7713
rect 9199 7687 9225 7713
rect 9255 7687 9281 7713
rect 12279 7687 12305 7713
rect 8919 7631 8945 7657
rect 9031 7631 9057 7657
rect 9927 7631 9953 7657
rect 10095 7631 10121 7657
rect 11047 7631 11073 7657
rect 11439 7631 11465 7657
rect 12783 7631 12809 7657
rect 13119 7631 13145 7657
rect 18831 7631 18857 7657
rect 10151 7575 10177 7601
rect 11103 7575 11129 7601
rect 14183 7575 14209 7601
rect 20007 7575 20033 7601
rect 12335 7519 12361 7545
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 9815 7351 9841 7377
rect 7687 7295 7713 7321
rect 8751 7295 8777 7321
rect 8975 7295 9001 7321
rect 9647 7295 9673 7321
rect 11047 7295 11073 7321
rect 12111 7295 12137 7321
rect 12727 7295 12753 7321
rect 13791 7295 13817 7321
rect 14015 7295 14041 7321
rect 7351 7239 7377 7265
rect 10711 7239 10737 7265
rect 12335 7239 12361 7265
rect 9703 7183 9729 7209
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 12279 6959 12305 6985
rect 9311 6903 9337 6929
rect 8751 6847 8777 6873
rect 8975 6847 9001 6873
rect 10375 6791 10401 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 8863 2143 8889 2169
rect 9367 2031 9393 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 9311 1807 9337 1833
rect 8975 1751 9001 1777
rect 10375 1751 10401 1777
rect 10879 1639 10905 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 11088 20600 11144 21000
rect 11424 20600 11480 21000
rect 11760 20600 11816 21000
rect 12096 20600 12152 21000
rect 12432 20600 12488 21000
rect 12768 20600 12824 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 11102 19138 11130 20600
rect 11214 19138 11242 19143
rect 11102 19137 11242 19138
rect 11102 19111 11215 19137
rect 11241 19111 11242 19137
rect 11102 19110 11242 19111
rect 11214 19105 11242 19110
rect 11438 19082 11466 20600
rect 11774 19418 11802 20600
rect 11774 19390 12026 19418
rect 11438 19049 11466 19054
rect 10878 19025 10906 19031
rect 10878 18999 10879 19025
rect 10905 18999 10906 19025
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 966 13593 994 13599
rect 966 13567 967 13593
rect 993 13567 994 13593
rect 966 13146 994 13567
rect 9422 13594 9450 13599
rect 9422 13593 9506 13594
rect 9422 13567 9423 13593
rect 9449 13567 9506 13593
rect 9422 13566 9506 13567
rect 9422 13561 9450 13566
rect 966 13113 994 13118
rect 2030 13537 2058 13543
rect 2030 13511 2031 13537
rect 2057 13511 2058 13537
rect 2030 13090 2058 13511
rect 8022 13537 8050 13543
rect 8022 13511 8023 13537
rect 8049 13511 8050 13537
rect 2030 13057 2058 13062
rect 2086 13482 2114 13487
rect 966 13033 994 13039
rect 966 13007 967 13033
rect 993 13007 994 13033
rect 966 12810 994 13007
rect 966 12777 994 12782
rect 966 12025 994 12031
rect 966 11999 967 12025
rect 993 11999 994 12025
rect 966 11802 994 11999
rect 966 11769 994 11774
rect 966 11466 994 11471
rect 966 11419 994 11438
rect 966 11241 994 11247
rect 966 11215 967 11241
rect 993 11215 994 11241
rect 966 10794 994 11215
rect 966 10761 994 10766
rect 966 10681 994 10687
rect 966 10655 967 10681
rect 993 10655 994 10681
rect 966 10458 994 10655
rect 966 10425 994 10430
rect 2086 10010 2114 13454
rect 6846 13481 6874 13487
rect 6846 13455 6847 13481
rect 6873 13455 6874 13481
rect 2142 13146 2170 13151
rect 2142 13099 2170 13118
rect 5558 13146 5586 13151
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 5558 12754 5586 13118
rect 6006 13090 6034 13095
rect 6006 13043 6034 13062
rect 6846 12810 6874 13455
rect 8022 13454 8050 13511
rect 8358 13481 8386 13487
rect 8358 13455 8359 13481
rect 8385 13455 8386 13481
rect 8358 13454 8386 13455
rect 6902 13426 6930 13431
rect 8022 13426 8106 13454
rect 8358 13426 8442 13454
rect 6902 13425 7098 13426
rect 6902 13399 6903 13425
rect 6929 13399 7098 13425
rect 6902 13398 7098 13399
rect 6902 13393 6930 13398
rect 7070 13201 7098 13398
rect 7070 13175 7071 13201
rect 7097 13175 7098 13201
rect 7070 13169 7098 13175
rect 7462 13230 7658 13258
rect 7462 13146 7490 13230
rect 7294 13145 7490 13146
rect 7294 13119 7463 13145
rect 7489 13119 7490 13145
rect 7294 13118 7490 13119
rect 7630 13146 7658 13230
rect 7686 13146 7714 13151
rect 7630 13118 7686 13146
rect 6846 12777 6874 12782
rect 7238 13090 7266 13095
rect 5558 12305 5586 12726
rect 6902 12754 6930 12759
rect 7014 12754 7042 12759
rect 6902 12707 6930 12726
rect 6958 12753 7042 12754
rect 6958 12727 7015 12753
rect 7041 12727 7042 12753
rect 6958 12726 7042 12727
rect 6342 12698 6370 12703
rect 6342 12651 6370 12670
rect 6790 12697 6818 12703
rect 6790 12671 6791 12697
rect 6817 12671 6818 12697
rect 6398 12642 6426 12647
rect 6790 12642 6818 12671
rect 6846 12698 6874 12703
rect 6846 12651 6874 12670
rect 6398 12641 6650 12642
rect 6398 12615 6399 12641
rect 6425 12615 6650 12641
rect 6398 12614 6650 12615
rect 6398 12609 6426 12614
rect 6622 12417 6650 12614
rect 6622 12391 6623 12417
rect 6649 12391 6650 12417
rect 6622 12385 6650 12391
rect 5558 12279 5559 12305
rect 5585 12279 5586 12305
rect 5558 12273 5586 12279
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 2142 11970 2170 11975
rect 6790 11970 6818 12614
rect 6958 11970 6986 12726
rect 7014 12721 7042 12726
rect 7238 12753 7266 13062
rect 7238 12727 7239 12753
rect 7265 12727 7266 12753
rect 7238 12721 7266 12727
rect 7238 12474 7266 12479
rect 7294 12474 7322 13118
rect 7462 13113 7490 13118
rect 7686 13099 7714 13118
rect 8078 13146 8106 13426
rect 8414 13257 8442 13426
rect 8414 13231 8415 13257
rect 8441 13231 8442 13257
rect 8414 13225 8442 13231
rect 7350 12810 7378 12815
rect 7350 12754 7378 12782
rect 7406 12754 7434 12759
rect 7350 12753 7434 12754
rect 7350 12727 7407 12753
rect 7433 12727 7434 12753
rect 7350 12726 7434 12727
rect 7406 12721 7434 12726
rect 7574 12753 7602 12759
rect 7574 12727 7575 12753
rect 7601 12727 7602 12753
rect 7518 12698 7546 12703
rect 7462 12670 7518 12698
rect 7350 12642 7378 12647
rect 7462 12642 7490 12670
rect 7518 12665 7546 12670
rect 7350 12595 7378 12614
rect 7406 12641 7490 12642
rect 7406 12615 7463 12641
rect 7489 12615 7490 12641
rect 7406 12614 7490 12615
rect 7014 12473 7322 12474
rect 7014 12447 7239 12473
rect 7265 12447 7322 12473
rect 7014 12446 7322 12447
rect 7014 12361 7042 12446
rect 7014 12335 7015 12361
rect 7041 12335 7042 12361
rect 7014 12329 7042 12335
rect 6790 11942 6874 11970
rect 6958 11942 7042 11970
rect 2142 11923 2170 11942
rect 6846 11914 6874 11942
rect 6846 11913 6986 11914
rect 6846 11887 6847 11913
rect 6873 11887 6986 11913
rect 6846 11886 6986 11887
rect 6846 11881 6874 11886
rect 5166 11858 5194 11863
rect 2142 11578 2170 11583
rect 2142 11531 2170 11550
rect 5166 11521 5194 11830
rect 6678 11858 6706 11863
rect 6790 11858 6818 11863
rect 6678 11857 6762 11858
rect 6678 11831 6679 11857
rect 6705 11831 6762 11857
rect 6678 11830 6762 11831
rect 6678 11825 6706 11830
rect 6622 11690 6650 11695
rect 5166 11495 5167 11521
rect 5193 11495 5194 11521
rect 5166 11489 5194 11495
rect 5950 11578 5978 11583
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 2142 11186 2170 11191
rect 2142 11139 2170 11158
rect 5838 11186 5866 11191
rect 2142 10794 2170 10799
rect 2142 10747 2170 10766
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 2086 9977 2114 9982
rect 2142 10066 2170 10071
rect 2142 10009 2170 10038
rect 2142 9983 2143 10009
rect 2169 9983 2170 10009
rect 2142 9977 2170 9983
rect 5726 10066 5754 10071
rect 5726 9954 5754 10038
rect 5726 9921 5754 9926
rect 5838 10066 5866 11158
rect 5950 10737 5978 11550
rect 6622 11577 6650 11662
rect 6734 11634 6762 11830
rect 6790 11811 6818 11830
rect 6790 11634 6818 11639
rect 6734 11633 6818 11634
rect 6734 11607 6791 11633
rect 6817 11607 6818 11633
rect 6734 11606 6818 11607
rect 6790 11601 6818 11606
rect 6846 11634 6874 11639
rect 6846 11587 6874 11606
rect 6622 11551 6623 11577
rect 6649 11551 6650 11577
rect 6622 11545 6650 11551
rect 6230 11521 6258 11527
rect 6230 11495 6231 11521
rect 6257 11495 6258 11521
rect 6230 11466 6258 11495
rect 6230 11433 6258 11438
rect 6846 11466 6874 11471
rect 6846 11419 6874 11438
rect 5950 10711 5951 10737
rect 5977 10711 5978 10737
rect 5950 10705 5978 10711
rect 6902 10514 6930 10519
rect 6902 10467 6930 10486
rect 6846 10345 6874 10351
rect 6846 10319 6847 10345
rect 6873 10319 6874 10345
rect 6846 10066 6874 10319
rect 6958 10094 6986 11886
rect 7014 11298 7042 11942
rect 7014 11265 7042 11270
rect 7126 11690 7154 12446
rect 7238 12441 7266 12446
rect 7126 10906 7154 11662
rect 7406 11298 7434 12614
rect 7462 12609 7490 12614
rect 7574 12586 7602 12727
rect 7574 12553 7602 12558
rect 7686 12754 7714 12759
rect 7686 11689 7714 12726
rect 8022 12697 8050 12703
rect 8022 12671 8023 12697
rect 8049 12671 8050 12697
rect 8022 12586 8050 12671
rect 8022 11802 8050 12558
rect 8078 11969 8106 13118
rect 8302 13145 8330 13151
rect 8302 13119 8303 13145
rect 8329 13119 8330 13145
rect 8302 12865 8330 13119
rect 9478 12922 9506 13566
rect 10710 13482 10738 13487
rect 10710 13481 10850 13482
rect 10710 13455 10711 13481
rect 10737 13455 10850 13481
rect 10710 13454 10850 13455
rect 10710 13449 10738 13454
rect 9646 13425 9674 13431
rect 9646 13399 9647 13425
rect 9673 13399 9674 13425
rect 9534 13146 9562 13151
rect 9646 13146 9674 13399
rect 10654 13425 10682 13431
rect 10654 13399 10655 13425
rect 10681 13399 10682 13425
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 10094 13202 10122 13207
rect 10654 13202 10682 13399
rect 10094 13201 10682 13202
rect 10094 13175 10095 13201
rect 10121 13175 10682 13201
rect 10094 13174 10682 13175
rect 10094 13169 10122 13174
rect 9702 13146 9730 13151
rect 9534 13145 9702 13146
rect 9534 13119 9535 13145
rect 9561 13119 9702 13145
rect 9534 13118 9702 13119
rect 9534 13113 9562 13118
rect 9702 13099 9730 13118
rect 10038 13146 10066 13151
rect 9478 12894 9618 12922
rect 8302 12839 8303 12865
rect 8329 12839 8330 12865
rect 8302 12833 8330 12839
rect 8134 12754 8162 12759
rect 8134 12707 8162 12726
rect 9590 12754 9618 12894
rect 9814 12754 9842 12759
rect 9590 12753 9842 12754
rect 9590 12727 9591 12753
rect 9617 12727 9815 12753
rect 9841 12727 9842 12753
rect 9590 12726 9842 12727
rect 9590 12721 9618 12726
rect 9814 12721 9842 12726
rect 9478 12642 9506 12647
rect 9982 12642 10010 12647
rect 9506 12614 9562 12642
rect 9478 12595 9506 12614
rect 9310 12418 9338 12423
rect 9310 12417 9450 12418
rect 9310 12391 9311 12417
rect 9337 12391 9450 12417
rect 9310 12390 9450 12391
rect 9310 12385 9338 12390
rect 8078 11943 8079 11969
rect 8105 11943 8106 11969
rect 8078 11937 8106 11943
rect 8414 11913 8442 11919
rect 8414 11887 8415 11913
rect 8441 11887 8442 11913
rect 8414 11858 8442 11887
rect 8414 11825 8442 11830
rect 8022 11769 8050 11774
rect 8806 11802 8834 11807
rect 7686 11663 7687 11689
rect 7713 11663 7714 11689
rect 7686 11657 7714 11663
rect 7574 11634 7602 11639
rect 7574 11587 7602 11606
rect 7798 11634 7826 11639
rect 7462 11578 7490 11583
rect 7462 11531 7490 11550
rect 7742 11577 7770 11583
rect 7742 11551 7743 11577
rect 7769 11551 7770 11577
rect 7630 11521 7658 11527
rect 7630 11495 7631 11521
rect 7657 11495 7658 11521
rect 7630 11354 7658 11495
rect 7518 11326 7658 11354
rect 7406 11297 7490 11298
rect 7406 11271 7407 11297
rect 7433 11271 7490 11297
rect 7406 11270 7490 11271
rect 7406 11265 7434 11270
rect 7350 11130 7378 11135
rect 7126 10873 7154 10878
rect 7182 11129 7378 11130
rect 7182 11103 7351 11129
rect 7377 11103 7378 11129
rect 7182 11102 7378 11103
rect 7014 10794 7042 10799
rect 7182 10794 7210 11102
rect 7350 11097 7378 11102
rect 7406 10906 7434 10911
rect 7406 10794 7434 10878
rect 7014 10793 7210 10794
rect 7014 10767 7015 10793
rect 7041 10767 7210 10793
rect 7014 10766 7210 10767
rect 7350 10793 7434 10794
rect 7350 10767 7407 10793
rect 7433 10767 7434 10793
rect 7350 10766 7434 10767
rect 7014 10761 7042 10766
rect 7014 10626 7042 10631
rect 7014 10513 7042 10598
rect 7014 10487 7015 10513
rect 7041 10487 7042 10513
rect 7014 10481 7042 10487
rect 7126 10402 7154 10407
rect 7126 10355 7154 10374
rect 7294 10345 7322 10351
rect 7294 10319 7295 10345
rect 7321 10319 7322 10345
rect 7294 10094 7322 10319
rect 6902 10066 6930 10071
rect 6958 10066 7042 10094
rect 6846 10065 6930 10066
rect 6846 10039 6903 10065
rect 6929 10039 6930 10065
rect 6846 10038 6930 10039
rect 5838 9953 5866 10038
rect 6902 10033 6930 10038
rect 5838 9927 5839 9953
rect 5865 9927 5866 9953
rect 5838 9921 5866 9927
rect 966 9898 994 9903
rect 966 9851 994 9870
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 6734 9561 6762 9567
rect 6734 9535 6735 9561
rect 6761 9535 6762 9561
rect 6454 9506 6482 9511
rect 2142 9226 2170 9231
rect 2142 9179 2170 9198
rect 5894 9226 5922 9231
rect 5390 9170 5418 9175
rect 966 9114 994 9119
rect 966 9067 994 9086
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 966 8890 994 8895
rect 966 8843 994 8862
rect 2142 8834 2170 8839
rect 2142 8787 2170 8806
rect 5390 8778 5418 9142
rect 5390 8745 5418 8750
rect 5894 8834 5922 9198
rect 6454 9225 6482 9478
rect 6454 9199 6455 9225
rect 6481 9199 6482 9225
rect 6454 9193 6482 9199
rect 6734 8946 6762 9535
rect 6790 9506 6818 9511
rect 6902 9506 6930 9511
rect 6790 9505 6874 9506
rect 6790 9479 6791 9505
rect 6817 9479 6874 9505
rect 6790 9478 6874 9479
rect 6790 9473 6818 9478
rect 6846 9338 6874 9478
rect 6902 9459 6930 9478
rect 7014 9505 7042 10066
rect 7238 10066 7322 10094
rect 7350 10122 7378 10766
rect 7406 10761 7434 10766
rect 7406 10682 7434 10687
rect 7406 10401 7434 10654
rect 7462 10514 7490 11270
rect 7518 11297 7546 11326
rect 7518 11271 7519 11297
rect 7545 11271 7546 11297
rect 7518 11265 7546 11271
rect 7574 11185 7602 11191
rect 7574 11159 7575 11185
rect 7601 11159 7602 11185
rect 7462 10481 7490 10486
rect 7518 10794 7546 10799
rect 7406 10375 7407 10401
rect 7433 10375 7434 10401
rect 7406 10369 7434 10375
rect 7462 10402 7490 10407
rect 7462 10289 7490 10374
rect 7462 10263 7463 10289
rect 7489 10263 7490 10289
rect 7462 10257 7490 10263
rect 7518 10178 7546 10766
rect 7574 10626 7602 11159
rect 7742 11074 7770 11551
rect 7798 11185 7826 11606
rect 7798 11159 7799 11185
rect 7825 11159 7826 11185
rect 7798 11153 7826 11159
rect 7966 11186 7994 11191
rect 7966 11139 7994 11158
rect 8750 11129 8778 11135
rect 8750 11103 8751 11129
rect 8777 11103 8778 11129
rect 7910 11074 7938 11079
rect 7742 11073 7938 11074
rect 7742 11047 7911 11073
rect 7937 11047 7938 11073
rect 7742 11046 7938 11047
rect 7630 10906 7658 10911
rect 7630 10859 7658 10878
rect 7910 10850 7938 11046
rect 7630 10626 7658 10631
rect 7574 10598 7630 10626
rect 7630 10593 7658 10598
rect 7238 10033 7266 10038
rect 7294 10010 7322 10015
rect 7350 10010 7378 10094
rect 7462 10150 7546 10178
rect 7574 10346 7602 10351
rect 7462 10065 7490 10150
rect 7574 10094 7602 10318
rect 7462 10039 7463 10065
rect 7489 10039 7490 10065
rect 7462 10033 7490 10039
rect 7518 10066 7602 10094
rect 7854 10345 7882 10351
rect 7854 10319 7855 10345
rect 7881 10319 7882 10345
rect 7854 10122 7882 10319
rect 7910 10346 7938 10822
rect 8694 10850 8722 10855
rect 8694 10803 8722 10822
rect 7910 10313 7938 10318
rect 8526 10738 8554 10743
rect 7630 10066 7658 10071
rect 7294 10009 7378 10010
rect 7294 9983 7295 10009
rect 7321 9983 7378 10009
rect 7294 9982 7378 9983
rect 7294 9977 7322 9982
rect 7014 9479 7015 9505
rect 7041 9479 7042 9505
rect 6846 9310 6986 9338
rect 6790 9282 6818 9287
rect 6790 9225 6818 9254
rect 6790 9199 6791 9225
rect 6817 9199 6818 9225
rect 6790 9193 6818 9199
rect 6958 9170 6986 9310
rect 6958 9137 6986 9142
rect 7014 9002 7042 9479
rect 7182 9730 7210 9735
rect 7182 9617 7210 9702
rect 7182 9591 7183 9617
rect 7209 9591 7210 9617
rect 7182 9281 7210 9591
rect 7182 9255 7183 9281
rect 7209 9255 7210 9281
rect 7182 9249 7210 9255
rect 7462 9282 7490 9287
rect 7518 9282 7546 10066
rect 7630 10019 7658 10038
rect 7742 9898 7770 9903
rect 7742 9673 7770 9870
rect 7742 9647 7743 9673
rect 7769 9647 7770 9673
rect 7742 9641 7770 9647
rect 7686 9282 7714 9287
rect 7462 9281 7546 9282
rect 7462 9255 7463 9281
rect 7489 9255 7546 9281
rect 7462 9254 7546 9255
rect 7574 9254 7686 9282
rect 7462 9249 7490 9254
rect 7294 9226 7322 9231
rect 7294 9179 7322 9198
rect 6846 8974 7042 9002
rect 7238 9169 7266 9175
rect 7238 9143 7239 9169
rect 7265 9143 7266 9169
rect 6790 8946 6818 8951
rect 6734 8945 6818 8946
rect 6734 8919 6791 8945
rect 6817 8919 6818 8945
rect 6734 8918 6818 8919
rect 6790 8913 6818 8918
rect 5894 8385 5922 8806
rect 6846 8833 6874 8974
rect 7238 8945 7266 9143
rect 7238 8919 7239 8945
rect 7265 8919 7266 8945
rect 7238 8913 7266 8919
rect 7070 8890 7098 8895
rect 6846 8807 6847 8833
rect 6873 8807 6874 8833
rect 6846 8801 6874 8807
rect 6958 8889 7098 8890
rect 6958 8863 7071 8889
rect 7097 8863 7098 8889
rect 6958 8862 7098 8863
rect 6790 8778 6818 8783
rect 6790 8731 6818 8750
rect 6958 8497 6986 8862
rect 7070 8857 7098 8862
rect 6958 8471 6959 8497
rect 6985 8471 6986 8497
rect 6958 8465 6986 8471
rect 7126 8721 7154 8727
rect 7126 8695 7127 8721
rect 7153 8695 7154 8721
rect 5894 8359 5895 8385
rect 5921 8359 5922 8385
rect 5894 8353 5922 8359
rect 7126 8330 7154 8695
rect 7574 8553 7602 9254
rect 7686 9235 7714 9254
rect 7854 9282 7882 10094
rect 7854 9249 7882 9254
rect 7574 8527 7575 8553
rect 7601 8527 7602 8553
rect 7126 8297 7154 8302
rect 7350 8441 7378 8447
rect 7350 8415 7351 8441
rect 7377 8415 7378 8441
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 7350 8050 7378 8415
rect 7574 8050 7602 8527
rect 8302 9002 8330 9007
rect 8302 8554 8330 8974
rect 8526 8722 8554 10710
rect 8750 10682 8778 11103
rect 8750 10649 8778 10654
rect 8806 11073 8834 11774
rect 9422 11578 9450 12390
rect 9478 12361 9506 12367
rect 9478 12335 9479 12361
rect 9505 12335 9506 12361
rect 9478 12026 9506 12335
rect 9478 11979 9506 11998
rect 9478 11578 9506 11583
rect 9422 11577 9506 11578
rect 9422 11551 9479 11577
rect 9505 11551 9506 11577
rect 9422 11550 9506 11551
rect 9422 11466 9450 11550
rect 9478 11545 9506 11550
rect 9142 11438 9422 11466
rect 8918 11186 8946 11191
rect 9142 11186 9170 11438
rect 9422 11419 9450 11438
rect 9534 11354 9562 12614
rect 9814 12641 10010 12642
rect 9814 12615 9983 12641
rect 10009 12615 10010 12641
rect 9814 12614 10010 12615
rect 10038 12642 10066 13118
rect 10822 12809 10850 13454
rect 10822 12783 10823 12809
rect 10849 12783 10850 12809
rect 10822 12777 10850 12783
rect 10878 13090 10906 18999
rect 11998 18353 12026 19390
rect 12110 18746 12138 20600
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 12222 18746 12250 18751
rect 12110 18745 12250 18746
rect 12110 18719 12223 18745
rect 12249 18719 12250 18745
rect 12110 18718 12250 18719
rect 12222 18713 12250 18718
rect 11998 18327 11999 18353
rect 12025 18327 12026 18353
rect 11998 18321 12026 18327
rect 11270 13538 11298 13543
rect 10598 12754 10626 12759
rect 10430 12698 10458 12703
rect 10038 12614 10122 12642
rect 9814 12418 9842 12614
rect 9982 12609 10010 12614
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9702 12417 9842 12418
rect 9702 12391 9815 12417
rect 9841 12391 9842 12417
rect 9702 12390 9842 12391
rect 9702 11970 9730 12390
rect 9814 12385 9842 12390
rect 9870 12418 9898 12423
rect 9870 12371 9898 12390
rect 9926 12417 9954 12423
rect 9926 12391 9927 12417
rect 9953 12391 9954 12417
rect 9926 12082 9954 12391
rect 9982 12082 10010 12087
rect 9478 11326 9562 11354
rect 9590 11942 9730 11970
rect 9478 11242 9506 11326
rect 8918 11185 9170 11186
rect 8918 11159 8919 11185
rect 8945 11159 9170 11185
rect 8918 11158 9170 11159
rect 8918 11153 8946 11158
rect 9142 11129 9170 11158
rect 9198 11214 9506 11242
rect 9198 11185 9226 11214
rect 9198 11159 9199 11185
rect 9225 11159 9226 11185
rect 9198 11153 9226 11159
rect 9478 11185 9506 11214
rect 9478 11159 9479 11185
rect 9505 11159 9506 11185
rect 9478 11153 9506 11159
rect 9142 11103 9143 11129
rect 9169 11103 9170 11129
rect 9142 11097 9170 11103
rect 9422 11129 9450 11135
rect 9422 11103 9423 11129
rect 9449 11103 9450 11129
rect 8806 11047 8807 11073
rect 8833 11047 8834 11073
rect 8638 10178 8666 10183
rect 8582 8834 8610 8839
rect 8638 8834 8666 10150
rect 8806 10009 8834 11047
rect 9030 11073 9058 11079
rect 9030 11047 9031 11073
rect 9057 11047 9058 11073
rect 8862 10906 8890 10911
rect 8862 10859 8890 10878
rect 8862 10458 8890 10463
rect 8862 10121 8890 10430
rect 8862 10095 8863 10121
rect 8889 10095 8890 10121
rect 8862 10089 8890 10095
rect 8806 9983 8807 10009
rect 8833 9983 8834 10009
rect 8806 9977 8834 9983
rect 8974 10009 9002 10015
rect 8974 9983 8975 10009
rect 9001 9983 9002 10009
rect 8918 9953 8946 9959
rect 8918 9927 8919 9953
rect 8945 9927 8946 9953
rect 8806 9561 8834 9567
rect 8806 9535 8807 9561
rect 8833 9535 8834 9561
rect 8806 9337 8834 9535
rect 8806 9311 8807 9337
rect 8833 9311 8834 9337
rect 8806 9305 8834 9311
rect 8862 9282 8890 9287
rect 8918 9282 8946 9927
rect 8974 9898 9002 9983
rect 8974 9865 9002 9870
rect 8862 9281 8946 9282
rect 8862 9255 8863 9281
rect 8889 9255 8946 9281
rect 8862 9254 8946 9255
rect 8862 9249 8890 9254
rect 8694 9225 8722 9231
rect 9030 9226 9058 11047
rect 9086 10849 9114 10855
rect 9086 10823 9087 10849
rect 9113 10823 9114 10849
rect 9086 10626 9114 10823
rect 9198 10794 9226 10799
rect 9198 10747 9226 10766
rect 9366 10738 9394 10743
rect 9422 10738 9450 11103
rect 9534 11129 9562 11135
rect 9534 11103 9535 11129
rect 9561 11103 9562 11129
rect 9534 10906 9562 11103
rect 9394 10710 9450 10738
rect 9478 10878 9534 10906
rect 9366 10705 9394 10710
rect 9086 10178 9114 10598
rect 9086 10145 9114 10150
rect 9142 10122 9170 10127
rect 8694 9199 8695 9225
rect 8721 9199 8722 9225
rect 8694 9002 8722 9199
rect 8694 8969 8722 8974
rect 8918 9198 9058 9226
rect 9086 10009 9114 10015
rect 9086 9983 9087 10009
rect 9113 9983 9114 10009
rect 9086 9562 9114 9983
rect 9142 9618 9170 10094
rect 9422 10065 9450 10071
rect 9422 10039 9423 10065
rect 9449 10039 9450 10065
rect 9142 9617 9338 9618
rect 9142 9591 9143 9617
rect 9169 9591 9338 9617
rect 9142 9590 9338 9591
rect 9142 9585 9170 9590
rect 8582 8833 8834 8834
rect 8582 8807 8583 8833
rect 8609 8807 8834 8833
rect 8582 8806 8834 8807
rect 8582 8801 8610 8806
rect 8638 8722 8666 8727
rect 8526 8721 8666 8722
rect 8526 8695 8639 8721
rect 8665 8695 8666 8721
rect 8526 8694 8666 8695
rect 8638 8689 8666 8694
rect 8750 8721 8778 8727
rect 8750 8695 8751 8721
rect 8777 8695 8778 8721
rect 8302 8507 8330 8526
rect 8694 8554 8722 8559
rect 8246 8330 8274 8335
rect 7966 8329 8274 8330
rect 7966 8303 8247 8329
rect 8273 8303 8274 8329
rect 7966 8302 8274 8303
rect 7966 8105 7994 8302
rect 8246 8297 8274 8302
rect 8414 8329 8442 8335
rect 8414 8303 8415 8329
rect 8441 8303 8442 8329
rect 8414 8274 8442 8303
rect 8414 8241 8442 8246
rect 7966 8079 7967 8105
rect 7993 8079 7994 8105
rect 7966 8073 7994 8079
rect 7350 8049 7602 8050
rect 7350 8023 7575 8049
rect 7601 8023 7602 8049
rect 7350 8022 7602 8023
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 7350 7265 7378 8022
rect 7574 8003 7602 8022
rect 8694 7713 8722 8526
rect 8694 7687 8695 7713
rect 8721 7687 8722 7713
rect 8694 7681 8722 7687
rect 8750 7714 8778 8695
rect 8806 8497 8834 8806
rect 8806 8471 8807 8497
rect 8833 8471 8834 8497
rect 8806 8465 8834 8471
rect 8918 8553 8946 9198
rect 8918 8527 8919 8553
rect 8945 8527 8946 8553
rect 8918 8442 8946 8527
rect 9086 8554 9114 9534
rect 9310 9226 9338 9590
rect 9422 9282 9450 10039
rect 9478 10065 9506 10878
rect 9534 10873 9562 10878
rect 9590 10849 9618 11942
rect 9590 10823 9591 10849
rect 9617 10823 9618 10849
rect 9590 10817 9618 10823
rect 9646 11858 9674 11863
rect 9646 10738 9674 11830
rect 9702 11578 9730 11942
rect 9814 12081 10010 12082
rect 9814 12055 9983 12081
rect 10009 12055 10010 12081
rect 9814 12054 10010 12055
rect 9814 11969 9842 12054
rect 9982 12049 10010 12054
rect 10038 12026 10066 12031
rect 10094 12026 10122 12614
rect 10262 12026 10290 12031
rect 10094 12025 10290 12026
rect 10094 11999 10263 12025
rect 10289 11999 10290 12025
rect 10094 11998 10290 11999
rect 10038 11979 10066 11998
rect 10262 11993 10290 11998
rect 9814 11943 9815 11969
rect 9841 11943 9842 11969
rect 9814 11937 9842 11943
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9702 11577 10066 11578
rect 9702 11551 9703 11577
rect 9729 11551 10066 11577
rect 9702 11550 10066 11551
rect 9702 11545 9730 11550
rect 9702 11465 9730 11471
rect 9702 11439 9703 11465
rect 9729 11439 9730 11465
rect 9702 11410 9730 11439
rect 9702 11186 9730 11382
rect 9926 11466 9954 11471
rect 9758 11298 9786 11303
rect 9758 11251 9786 11270
rect 9926 11241 9954 11438
rect 10038 11297 10066 11550
rect 10038 11271 10039 11297
rect 10065 11271 10066 11297
rect 10038 11265 10066 11271
rect 9926 11215 9927 11241
rect 9953 11215 9954 11241
rect 9926 11209 9954 11215
rect 9702 11153 9730 11158
rect 10206 11074 10234 11079
rect 10206 11073 10346 11074
rect 10206 11047 10207 11073
rect 10233 11047 10346 11073
rect 10206 11046 10346 11047
rect 10206 11041 10234 11046
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 9646 10705 9674 10710
rect 10038 10850 10066 10855
rect 10038 10793 10066 10822
rect 10038 10767 10039 10793
rect 10065 10767 10066 10793
rect 9534 10682 9562 10687
rect 9534 10635 9562 10654
rect 10038 10514 10066 10767
rect 10094 10793 10122 10799
rect 10094 10767 10095 10793
rect 10121 10767 10122 10793
rect 10094 10738 10122 10767
rect 10262 10794 10290 10799
rect 10262 10747 10290 10766
rect 10094 10705 10122 10710
rect 10206 10737 10234 10743
rect 10206 10711 10207 10737
rect 10233 10711 10234 10737
rect 10206 10570 10234 10711
rect 10206 10537 10234 10542
rect 10038 10486 10178 10514
rect 10038 10402 10066 10407
rect 10038 10355 10066 10374
rect 9478 10039 9479 10065
rect 9505 10039 9506 10065
rect 9478 10033 9506 10039
rect 9814 10290 9842 10295
rect 9702 10010 9730 10015
rect 9590 9982 9702 10010
rect 9534 9898 9562 9903
rect 9534 9851 9562 9870
rect 9534 9562 9562 9567
rect 9534 9515 9562 9534
rect 9590 9337 9618 9982
rect 9702 9963 9730 9982
rect 9702 9842 9730 9847
rect 9702 9617 9730 9814
rect 9702 9591 9703 9617
rect 9729 9591 9730 9617
rect 9702 9585 9730 9591
rect 9814 9618 9842 10262
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 10094 9898 10122 9903
rect 9982 9730 10010 9735
rect 9982 9673 10010 9702
rect 9982 9647 9983 9673
rect 10009 9647 10010 9673
rect 9982 9641 10010 9647
rect 9870 9618 9898 9623
rect 9814 9617 9898 9618
rect 9814 9591 9871 9617
rect 9897 9591 9898 9617
rect 9814 9590 9898 9591
rect 9870 9585 9898 9590
rect 10038 9561 10066 9567
rect 10038 9535 10039 9561
rect 10065 9535 10066 9561
rect 10038 9506 10066 9535
rect 10038 9473 10066 9478
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9590 9311 9591 9337
rect 9617 9311 9618 9337
rect 9590 9305 9618 9311
rect 9422 9249 9450 9254
rect 9310 9225 9394 9226
rect 9310 9199 9311 9225
rect 9337 9199 9394 9225
rect 9310 9198 9394 9199
rect 9310 9193 9338 9198
rect 9086 8553 9170 8554
rect 9086 8527 9087 8553
rect 9113 8527 9170 8553
rect 9086 8526 9170 8527
rect 9086 8521 9114 8526
rect 9142 8498 9170 8526
rect 9142 8470 9338 8498
rect 8918 8409 8946 8414
rect 9030 8441 9058 8447
rect 9030 8415 9031 8441
rect 9057 8415 9058 8441
rect 8974 8385 9002 8391
rect 8974 8359 8975 8385
rect 9001 8359 9002 8385
rect 8974 8274 9002 8359
rect 8974 8241 9002 8246
rect 9030 8106 9058 8415
rect 9254 8106 9282 8111
rect 8974 8105 9058 8106
rect 8974 8079 9031 8105
rect 9057 8079 9058 8105
rect 8974 8078 9058 8079
rect 8806 7714 8834 7719
rect 8750 7713 8834 7714
rect 8750 7687 8807 7713
rect 8833 7687 8834 7713
rect 8750 7686 8834 7687
rect 8806 7681 8834 7686
rect 8862 7714 8890 7719
rect 7686 7658 7714 7663
rect 7686 7321 7714 7630
rect 8862 7574 8890 7686
rect 8918 7658 8946 7663
rect 8918 7611 8946 7630
rect 8750 7546 8890 7574
rect 8974 7574 9002 8078
rect 9030 8073 9058 8078
rect 9142 8078 9254 8106
rect 9086 7714 9114 7719
rect 9030 7713 9114 7714
rect 9030 7687 9087 7713
rect 9113 7687 9114 7713
rect 9030 7686 9114 7687
rect 9030 7657 9058 7686
rect 9086 7681 9114 7686
rect 9030 7631 9031 7657
rect 9057 7631 9058 7657
rect 9030 7625 9058 7631
rect 9142 7658 9170 8078
rect 9254 8059 9282 8078
rect 9198 7714 9226 7719
rect 9198 7667 9226 7686
rect 9254 7714 9282 7719
rect 9310 7714 9338 8470
rect 9366 8106 9394 9198
rect 9646 9170 9674 9175
rect 9646 8833 9674 9142
rect 10094 9169 10122 9870
rect 10094 9143 10095 9169
rect 10121 9143 10122 9169
rect 10094 9137 10122 9143
rect 10150 9058 10178 10486
rect 10318 10122 10346 11046
rect 10430 10905 10458 12670
rect 10598 12473 10626 12726
rect 10766 12754 10794 12759
rect 10766 12707 10794 12726
rect 10878 12753 10906 13062
rect 10878 12727 10879 12753
rect 10905 12727 10906 12753
rect 10878 12721 10906 12727
rect 10990 13537 11298 13538
rect 10990 13511 11271 13537
rect 11297 13511 11298 13537
rect 10990 13510 11298 13511
rect 10654 12698 10682 12703
rect 10654 12651 10682 12670
rect 10934 12641 10962 12647
rect 10934 12615 10935 12641
rect 10961 12615 10962 12641
rect 10934 12474 10962 12615
rect 10598 12447 10599 12473
rect 10625 12447 10626 12473
rect 10486 12418 10514 12423
rect 10486 12361 10514 12390
rect 10486 12335 10487 12361
rect 10513 12335 10514 12361
rect 10486 12329 10514 12335
rect 10598 11186 10626 12447
rect 10878 12446 10962 12474
rect 10878 12250 10906 12446
rect 10934 12362 10962 12367
rect 10990 12362 11018 13510
rect 11270 13505 11298 13510
rect 11662 13482 11690 13487
rect 11606 13481 11690 13482
rect 11606 13455 11663 13481
rect 11689 13455 11690 13481
rect 11606 13454 11690 13455
rect 11494 13426 11634 13454
rect 11662 13449 11690 13454
rect 11158 13090 11186 13095
rect 11158 13043 11186 13062
rect 11494 12809 11522 13426
rect 11494 12783 11495 12809
rect 11521 12783 11522 12809
rect 11494 12777 11522 12783
rect 11662 12810 11690 12815
rect 11662 12763 11690 12782
rect 12110 12810 12138 12815
rect 12110 12763 12138 12782
rect 11606 12753 11634 12759
rect 11606 12727 11607 12753
rect 11633 12727 11634 12753
rect 11438 12697 11466 12703
rect 11438 12671 11439 12697
rect 11465 12671 11466 12697
rect 11438 12586 11466 12671
rect 10934 12361 10990 12362
rect 10934 12335 10935 12361
rect 10961 12335 10990 12361
rect 10934 12334 10990 12335
rect 10934 12329 10962 12334
rect 10990 12315 11018 12334
rect 11214 12558 11466 12586
rect 11606 12642 11634 12727
rect 10878 12222 10962 12250
rect 10598 11153 10626 11158
rect 10430 10879 10431 10905
rect 10457 10879 10458 10905
rect 10430 10873 10458 10879
rect 10934 10906 10962 12222
rect 11214 11690 11242 12558
rect 11438 12474 11466 12479
rect 11214 11522 11242 11662
rect 11270 12305 11298 12311
rect 11270 12279 11271 12305
rect 11297 12279 11298 12305
rect 11270 11634 11298 12279
rect 11438 11969 11466 12446
rect 11550 12418 11578 12423
rect 11550 12025 11578 12390
rect 11550 11999 11551 12025
rect 11577 11999 11578 12025
rect 11550 11993 11578 11999
rect 11438 11943 11439 11969
rect 11465 11943 11466 11969
rect 11438 11774 11466 11943
rect 11382 11746 11466 11774
rect 11494 11857 11522 11863
rect 11494 11831 11495 11857
rect 11521 11831 11522 11857
rect 11494 11802 11522 11831
rect 11494 11746 11578 11802
rect 11382 11713 11410 11718
rect 11494 11713 11522 11718
rect 11270 11601 11298 11606
rect 11326 11690 11354 11695
rect 11326 11633 11354 11662
rect 11326 11607 11327 11633
rect 11353 11607 11354 11633
rect 11326 11601 11354 11607
rect 11550 11634 11578 11639
rect 11382 11578 11410 11583
rect 11382 11531 11410 11550
rect 11494 11577 11522 11583
rect 11494 11551 11495 11577
rect 11521 11551 11522 11577
rect 11214 11494 11354 11522
rect 11214 11186 11242 11191
rect 11214 11139 11242 11158
rect 10934 10873 10962 10878
rect 11046 11130 11074 11135
rect 11046 10905 11074 11102
rect 11046 10879 11047 10905
rect 11073 10879 11074 10905
rect 11046 10873 11074 10879
rect 10878 10849 10906 10855
rect 10878 10823 10879 10849
rect 10905 10823 10906 10849
rect 10318 10089 10346 10094
rect 10598 10793 10626 10799
rect 10598 10767 10599 10793
rect 10625 10767 10626 10793
rect 10598 9618 10626 10767
rect 10710 10794 10738 10799
rect 10710 10457 10738 10766
rect 10710 10431 10711 10457
rect 10737 10431 10738 10457
rect 10710 10425 10738 10431
rect 10766 10682 10794 10687
rect 10766 10401 10794 10654
rect 10878 10458 10906 10823
rect 10990 10793 11018 10799
rect 10990 10767 10991 10793
rect 11017 10767 11018 10793
rect 10990 10682 11018 10767
rect 11102 10794 11130 10799
rect 11102 10793 11242 10794
rect 11102 10767 11103 10793
rect 11129 10767 11242 10793
rect 11102 10766 11242 10767
rect 11102 10761 11130 10766
rect 10990 10649 11018 10654
rect 10878 10430 11018 10458
rect 10766 10375 10767 10401
rect 10793 10375 10794 10401
rect 10766 10369 10794 10375
rect 10654 10345 10682 10351
rect 10654 10319 10655 10345
rect 10681 10319 10682 10345
rect 10654 10290 10682 10319
rect 10654 10257 10682 10262
rect 10934 10345 10962 10351
rect 10934 10319 10935 10345
rect 10961 10319 10962 10345
rect 10934 9842 10962 10319
rect 10990 10290 11018 10430
rect 11158 10345 11186 10351
rect 11158 10319 11159 10345
rect 11185 10319 11186 10345
rect 11102 10290 11130 10295
rect 10990 10289 11130 10290
rect 10990 10263 11103 10289
rect 11129 10263 11130 10289
rect 10990 10262 11130 10263
rect 10934 9809 10962 9814
rect 10990 10122 11018 10127
rect 10990 9674 11018 10094
rect 10598 9585 10626 9590
rect 10934 9646 11018 9674
rect 10934 9617 10962 9646
rect 10934 9591 10935 9617
rect 10961 9591 10962 9617
rect 10934 9585 10962 9591
rect 10206 9505 10234 9511
rect 10206 9479 10207 9505
rect 10233 9479 10234 9505
rect 10206 9114 10234 9479
rect 10374 9506 10402 9511
rect 10374 9459 10402 9478
rect 10710 9505 10738 9511
rect 10710 9479 10711 9505
rect 10737 9479 10738 9505
rect 10318 9114 10346 9119
rect 10206 9086 10318 9114
rect 10094 9030 10178 9058
rect 9758 9002 9786 9007
rect 9758 8945 9786 8974
rect 9758 8919 9759 8945
rect 9785 8919 9786 8945
rect 9758 8913 9786 8919
rect 9646 8807 9647 8833
rect 9673 8807 9674 8833
rect 9646 8778 9674 8807
rect 9646 8745 9674 8750
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 10094 8554 10122 9030
rect 10206 8834 10234 8839
rect 10206 8787 10234 8806
rect 10318 8833 10346 9086
rect 10318 8807 10319 8833
rect 10345 8807 10346 8833
rect 10318 8801 10346 8807
rect 10654 8834 10682 8839
rect 10654 8554 10682 8806
rect 10710 8778 10738 9479
rect 10822 9505 10850 9511
rect 10822 9479 10823 9505
rect 10849 9479 10850 9505
rect 10822 9114 10850 9479
rect 10878 9505 10906 9511
rect 10878 9479 10879 9505
rect 10905 9479 10906 9505
rect 10878 9226 10906 9479
rect 11102 9506 11130 10262
rect 11158 9898 11186 10319
rect 11214 10290 11242 10766
rect 11214 10257 11242 10262
rect 11270 10793 11298 10799
rect 11270 10767 11271 10793
rect 11297 10767 11298 10793
rect 11158 9865 11186 9870
rect 11214 10122 11242 10127
rect 11158 9618 11186 9623
rect 11158 9571 11186 9590
rect 10878 9193 10906 9198
rect 10934 9282 10962 9287
rect 10822 9081 10850 9086
rect 10710 8722 10738 8750
rect 10878 9058 10906 9063
rect 10766 8722 10794 8727
rect 10710 8721 10794 8722
rect 10710 8695 10767 8721
rect 10793 8695 10794 8721
rect 10710 8694 10794 8695
rect 10766 8689 10794 8694
rect 10094 8526 10514 8554
rect 9982 8386 10010 8391
rect 9982 8339 10010 8358
rect 10094 8385 10122 8526
rect 10150 8442 10178 8447
rect 10150 8441 10234 8442
rect 10150 8415 10151 8441
rect 10177 8415 10234 8441
rect 10150 8414 10234 8415
rect 10150 8409 10178 8414
rect 10094 8359 10095 8385
rect 10121 8359 10122 8385
rect 10094 8353 10122 8359
rect 9366 8073 9394 8078
rect 9702 8330 9730 8335
rect 9254 7713 9310 7714
rect 9254 7687 9255 7713
rect 9281 7687 9310 7713
rect 9254 7686 9310 7687
rect 9254 7681 9282 7686
rect 9310 7667 9338 7686
rect 9142 7625 9170 7630
rect 8974 7546 9170 7574
rect 8750 7322 8778 7546
rect 9030 7490 9058 7495
rect 7686 7295 7687 7321
rect 7713 7295 7714 7321
rect 7686 7289 7714 7295
rect 8694 7321 8778 7322
rect 8694 7295 8751 7321
rect 8777 7295 8778 7321
rect 8694 7294 8778 7295
rect 7350 7239 7351 7265
rect 7377 7239 7378 7265
rect 7350 7233 7378 7239
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 8694 2170 8722 7294
rect 8750 7289 8778 7294
rect 8974 7462 9030 7490
rect 8974 7321 9002 7462
rect 8974 7295 8975 7321
rect 9001 7295 9002 7321
rect 8974 7289 9002 7295
rect 8750 6874 8778 6879
rect 8974 6874 9002 6879
rect 9030 6874 9058 7462
rect 8750 6873 9058 6874
rect 8750 6847 8751 6873
rect 8777 6847 8975 6873
rect 9001 6847 9058 6873
rect 8750 6846 9058 6847
rect 8750 6841 8778 6846
rect 8974 6841 9002 6846
rect 9142 5894 9170 7546
rect 9646 7322 9674 7327
rect 9310 7321 9674 7322
rect 9310 7295 9647 7321
rect 9673 7295 9674 7321
rect 9310 7294 9674 7295
rect 9310 6929 9338 7294
rect 9646 7289 9674 7294
rect 9702 7209 9730 8302
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 10206 7770 10234 8414
rect 10486 8218 10514 8526
rect 10654 8507 10682 8526
rect 10542 8386 10570 8391
rect 10542 8339 10570 8358
rect 10598 8385 10626 8391
rect 10598 8359 10599 8385
rect 10625 8359 10626 8385
rect 10598 8330 10626 8359
rect 10626 8302 10794 8330
rect 10598 8297 10626 8302
rect 10486 8190 10682 8218
rect 10654 8049 10682 8190
rect 10766 8161 10794 8302
rect 10766 8135 10767 8161
rect 10793 8135 10794 8161
rect 10766 8129 10794 8135
rect 10878 8161 10906 9030
rect 10934 8778 10962 9254
rect 10934 8777 11018 8778
rect 10934 8751 10935 8777
rect 10961 8751 11018 8777
rect 10934 8750 11018 8751
rect 10934 8745 10962 8750
rect 10990 8554 11018 8750
rect 11102 8777 11130 9478
rect 11158 9226 11186 9231
rect 11158 9179 11186 9198
rect 11214 8834 11242 10094
rect 11270 9730 11298 10767
rect 11326 10458 11354 11494
rect 11494 11466 11522 11551
rect 11550 11577 11578 11606
rect 11550 11551 11551 11577
rect 11577 11551 11578 11577
rect 11550 11545 11578 11551
rect 11606 11466 11634 12614
rect 11718 12753 11746 12759
rect 11718 12727 11719 12753
rect 11745 12727 11746 12753
rect 11662 11969 11690 11975
rect 11662 11943 11663 11969
rect 11689 11943 11690 11969
rect 11662 11746 11690 11943
rect 11662 11713 11690 11718
rect 11718 11578 11746 12727
rect 11494 11438 11634 11466
rect 11662 11577 11746 11578
rect 11662 11551 11719 11577
rect 11745 11551 11746 11577
rect 11662 11550 11746 11551
rect 11494 11298 11522 11303
rect 11382 11186 11410 11191
rect 11382 11139 11410 11158
rect 11438 11185 11466 11191
rect 11438 11159 11439 11185
rect 11465 11159 11466 11185
rect 11438 11018 11466 11159
rect 11494 11185 11522 11270
rect 11494 11159 11495 11185
rect 11521 11159 11522 11185
rect 11494 11153 11522 11159
rect 11606 11074 11634 11079
rect 11606 11027 11634 11046
rect 11382 10990 11466 11018
rect 11382 10850 11410 10990
rect 11438 10906 11466 10911
rect 11438 10859 11466 10878
rect 11382 10817 11410 10822
rect 11326 10425 11354 10430
rect 11438 10514 11466 10519
rect 11662 10514 11690 11550
rect 11718 11545 11746 11550
rect 11774 12754 11802 12759
rect 11774 11913 11802 12726
rect 12222 12754 12250 12759
rect 12222 12707 12250 12726
rect 12054 12641 12082 12647
rect 12054 12615 12055 12641
rect 12081 12615 12082 12641
rect 12054 12418 12082 12615
rect 12110 12641 12138 12647
rect 12110 12615 12111 12641
rect 12137 12615 12138 12641
rect 12110 12474 12138 12615
rect 12110 12441 12138 12446
rect 12054 12385 12082 12390
rect 12278 12306 12306 18999
rect 12446 18746 12474 20600
rect 12782 19138 12810 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 12782 19105 12810 19110
rect 14686 19138 14714 19143
rect 14686 19091 14714 19110
rect 12838 19082 12866 19087
rect 12838 19035 12866 19054
rect 14294 19025 14322 19031
rect 14294 18999 14295 19025
rect 14321 18999 14322 19025
rect 12446 18713 12474 18718
rect 13118 18746 13146 18751
rect 13118 18699 13146 18718
rect 12838 18634 12866 18639
rect 12838 18633 12922 18634
rect 12838 18607 12839 18633
rect 12865 18607 12922 18633
rect 12838 18606 12922 18607
rect 12838 18601 12866 18606
rect 12726 13593 12754 13599
rect 12726 13567 12727 13593
rect 12753 13567 12754 13593
rect 12726 13454 12754 13567
rect 12894 13481 12922 18606
rect 12894 13455 12895 13481
rect 12921 13455 12922 13481
rect 12670 13426 12866 13454
rect 12894 13449 12922 13455
rect 12950 18241 12978 18247
rect 12950 18215 12951 18241
rect 12977 18215 12978 18241
rect 12950 13538 12978 18215
rect 13006 13538 13034 13543
rect 12950 13537 13034 13538
rect 12950 13511 13007 13537
rect 13033 13511 13034 13537
rect 12950 13510 13034 13511
rect 12334 13146 12362 13151
rect 12334 12753 12362 13118
rect 12670 13146 12698 13426
rect 12838 13370 12866 13426
rect 12950 13370 12978 13510
rect 13006 13505 13034 13510
rect 13286 13481 13314 13487
rect 13286 13455 13287 13481
rect 13313 13455 13314 13481
rect 13286 13454 13314 13455
rect 12838 13342 12978 13370
rect 13118 13426 13314 13454
rect 12782 13258 12810 13263
rect 12782 13211 12810 13230
rect 12670 13099 12698 13118
rect 12334 12727 12335 12753
rect 12361 12727 12362 12753
rect 12334 12721 12362 12727
rect 12670 12362 12698 12367
rect 12670 12315 12698 12334
rect 13118 12362 13146 13426
rect 14294 13258 14322 18999
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 20118 18129 20146 18135
rect 20118 18103 20119 18129
rect 20145 18103 20146 18129
rect 20118 17850 20146 18103
rect 20118 17817 20146 17822
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 14294 13225 14322 13230
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 20006 12809 20034 12815
rect 20006 12783 20007 12809
rect 20033 12783 20034 12809
rect 18830 12753 18858 12759
rect 18830 12727 18831 12753
rect 18857 12727 18858 12753
rect 13454 12698 13482 12703
rect 12334 12306 12362 12311
rect 11942 12305 12362 12306
rect 11942 12279 12335 12305
rect 12361 12279 12362 12305
rect 11942 12278 12362 12279
rect 11942 11969 11970 12278
rect 12334 12273 12362 12278
rect 11942 11943 11943 11969
rect 11969 11943 11970 11969
rect 11942 11937 11970 11943
rect 11774 11887 11775 11913
rect 11801 11887 11802 11913
rect 11774 11242 11802 11887
rect 13118 11802 13146 12334
rect 13342 12697 13482 12698
rect 13342 12671 13455 12697
rect 13481 12671 13482 12697
rect 13342 12670 13482 12671
rect 13342 12025 13370 12670
rect 13454 12665 13482 12670
rect 13510 12641 13538 12647
rect 13510 12615 13511 12641
rect 13537 12615 13538 12641
rect 13510 12417 13538 12615
rect 13510 12391 13511 12417
rect 13537 12391 13538 12417
rect 13510 12385 13538 12391
rect 13342 11999 13343 12025
rect 13369 11999 13370 12025
rect 13342 11993 13370 11999
rect 13398 12306 13426 12311
rect 13118 11769 13146 11774
rect 13230 11969 13258 11975
rect 13230 11943 13231 11969
rect 13257 11943 13258 11969
rect 11830 11690 11858 11695
rect 11830 11298 11858 11662
rect 11830 11265 11858 11270
rect 12110 11298 12138 11303
rect 12110 11251 12138 11270
rect 11718 11214 11802 11242
rect 12278 11242 12306 11247
rect 12278 11241 12362 11242
rect 12278 11215 12279 11241
rect 12305 11215 12362 11241
rect 12278 11214 12362 11215
rect 11718 11130 11746 11214
rect 12278 11209 12306 11214
rect 11718 11097 11746 11102
rect 11942 11186 11970 11191
rect 11942 11129 11970 11158
rect 11942 11103 11943 11129
rect 11969 11103 11970 11129
rect 11942 11097 11970 11103
rect 12222 11186 12250 11191
rect 12222 11129 12250 11158
rect 12222 11103 12223 11129
rect 12249 11103 12250 11129
rect 12222 11097 12250 11103
rect 11438 10457 11466 10486
rect 11438 10431 11439 10457
rect 11465 10431 11466 10457
rect 11438 10425 11466 10431
rect 11606 10486 11690 10514
rect 11774 11073 11802 11079
rect 11774 11047 11775 11073
rect 11801 11047 11802 11073
rect 11774 10793 11802 11047
rect 11774 10767 11775 10793
rect 11801 10767 11802 10793
rect 11774 10514 11802 10767
rect 11494 10345 11522 10351
rect 11494 10319 11495 10345
rect 11521 10319 11522 10345
rect 11270 9697 11298 9702
rect 11382 10290 11410 10295
rect 11326 9506 11354 9511
rect 11270 9505 11354 9506
rect 11270 9479 11327 9505
rect 11353 9479 11354 9505
rect 11270 9478 11354 9479
rect 11270 9450 11298 9478
rect 11326 9473 11354 9478
rect 11270 9058 11298 9422
rect 11382 9394 11410 10262
rect 11494 9898 11522 10319
rect 11494 9617 11522 9870
rect 11494 9591 11495 9617
rect 11521 9591 11522 9617
rect 11494 9585 11522 9591
rect 11606 9450 11634 10486
rect 11774 10481 11802 10486
rect 11886 10849 11914 10855
rect 11886 10823 11887 10849
rect 11913 10823 11914 10849
rect 11886 10794 11914 10823
rect 11886 10458 11914 10766
rect 11886 10425 11914 10430
rect 11662 10402 11690 10407
rect 11662 10065 11690 10374
rect 11662 10039 11663 10065
rect 11689 10039 11690 10065
rect 11662 10033 11690 10039
rect 12278 9954 12306 9959
rect 11662 9842 11690 9847
rect 11662 9561 11690 9814
rect 12278 9673 12306 9926
rect 12278 9647 12279 9673
rect 12305 9647 12306 9673
rect 12278 9641 12306 9647
rect 11662 9535 11663 9561
rect 11689 9535 11690 9561
rect 11662 9529 11690 9535
rect 11718 9618 11746 9623
rect 11606 9417 11634 9422
rect 11270 9025 11298 9030
rect 11326 9366 11410 9394
rect 11214 8833 11298 8834
rect 11214 8807 11215 8833
rect 11241 8807 11298 8833
rect 11214 8806 11298 8807
rect 11214 8801 11242 8806
rect 11102 8751 11103 8777
rect 11129 8751 11130 8777
rect 11102 8745 11130 8751
rect 11214 8554 11242 8559
rect 10990 8553 11242 8554
rect 10990 8527 11215 8553
rect 11241 8527 11242 8553
rect 10990 8526 11242 8527
rect 10878 8135 10879 8161
rect 10905 8135 10906 8161
rect 10878 8129 10906 8135
rect 10654 8023 10655 8049
rect 10681 8023 10682 8049
rect 10654 8017 10682 8023
rect 10206 7723 10234 7742
rect 10934 7993 10962 7999
rect 10934 7967 10935 7993
rect 10961 7967 10962 7993
rect 9926 7714 9954 7719
rect 9926 7657 9954 7686
rect 9926 7631 9927 7657
rect 9953 7631 9954 7657
rect 9926 7625 9954 7631
rect 10094 7657 10122 7663
rect 10094 7631 10095 7657
rect 10121 7631 10122 7657
rect 9814 7602 9842 7607
rect 9814 7377 9842 7574
rect 9814 7351 9815 7377
rect 9841 7351 9842 7377
rect 9814 7345 9842 7351
rect 9702 7183 9703 7209
rect 9729 7183 9730 7209
rect 9702 7177 9730 7183
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9310 6903 9311 6929
rect 9337 6903 9338 6929
rect 9310 6897 9338 6903
rect 10094 6818 10122 7631
rect 10150 7602 10178 7621
rect 10150 7569 10178 7574
rect 10934 7574 10962 7967
rect 11102 7882 11130 8526
rect 11214 8521 11242 8526
rect 11270 8442 11298 8806
rect 11214 8414 11298 8442
rect 11214 8386 11242 8414
rect 11326 8386 11354 9366
rect 11550 9226 11578 9231
rect 11550 9179 11578 9198
rect 11718 9169 11746 9590
rect 12222 9617 12250 9623
rect 12222 9591 12223 9617
rect 12249 9591 12250 9617
rect 12054 9561 12082 9567
rect 12054 9535 12055 9561
rect 12081 9535 12082 9561
rect 12054 9450 12082 9535
rect 12222 9562 12250 9591
rect 12334 9617 12362 11214
rect 12838 10850 12866 10855
rect 12334 9591 12335 9617
rect 12361 9591 12362 9617
rect 12334 9585 12362 9591
rect 12670 10122 12698 10127
rect 12670 10009 12698 10094
rect 12670 9983 12671 10009
rect 12697 9983 12698 10009
rect 12222 9529 12250 9534
rect 12054 9417 12082 9422
rect 11774 9282 11802 9287
rect 11774 9235 11802 9254
rect 12110 9226 12138 9231
rect 12110 9179 12138 9198
rect 12670 9226 12698 9983
rect 12698 9198 12810 9226
rect 12670 9193 12698 9198
rect 11718 9143 11719 9169
rect 11745 9143 11746 9169
rect 11718 9137 11746 9143
rect 11886 9114 11914 9119
rect 11886 8722 11914 9086
rect 11886 8689 11914 8694
rect 12726 8721 12754 8727
rect 12726 8695 12727 8721
rect 12753 8695 12754 8721
rect 11382 8554 11410 8559
rect 11382 8507 11410 8526
rect 12726 8554 12754 8695
rect 12726 8521 12754 8526
rect 11214 8353 11242 8358
rect 11270 8358 11354 8386
rect 12502 8386 12530 8391
rect 11158 7994 11186 7999
rect 11270 7994 11298 8358
rect 12502 8049 12530 8358
rect 12502 8023 12503 8049
rect 12529 8023 12530 8049
rect 12502 8017 12530 8023
rect 11158 7993 11298 7994
rect 11158 7967 11159 7993
rect 11185 7967 11298 7993
rect 11158 7966 11298 7967
rect 11158 7961 11186 7966
rect 11326 7937 11354 7943
rect 11326 7911 11327 7937
rect 11353 7911 11354 7937
rect 11102 7854 11298 7882
rect 11270 7769 11298 7854
rect 11270 7743 11271 7769
rect 11297 7743 11298 7769
rect 11270 7737 11298 7743
rect 11326 7770 11354 7911
rect 12614 7937 12642 7943
rect 12614 7911 12615 7937
rect 12641 7911 12642 7937
rect 11606 7770 11634 7775
rect 11326 7769 11634 7770
rect 11326 7743 11607 7769
rect 11633 7743 11634 7769
rect 11326 7742 11634 7743
rect 11046 7657 11074 7663
rect 11046 7631 11047 7657
rect 11073 7631 11074 7657
rect 10934 7546 11018 7574
rect 10990 7322 11018 7546
rect 11046 7546 11074 7631
rect 11102 7602 11130 7607
rect 11326 7602 11354 7742
rect 11606 7737 11634 7742
rect 11774 7770 11802 7775
rect 11774 7723 11802 7742
rect 12614 7770 12642 7911
rect 12614 7737 12642 7742
rect 12670 7937 12698 7943
rect 12670 7911 12671 7937
rect 12697 7911 12698 7937
rect 12278 7714 12306 7719
rect 12278 7667 12306 7686
rect 11102 7601 11354 7602
rect 11102 7575 11103 7601
rect 11129 7575 11354 7601
rect 11102 7574 11354 7575
rect 11438 7657 11466 7663
rect 11438 7631 11439 7657
rect 11465 7631 11466 7657
rect 11102 7569 11130 7574
rect 11046 7513 11074 7518
rect 11438 7546 11466 7631
rect 12670 7658 12698 7911
rect 12726 7938 12754 7943
rect 12726 7891 12754 7910
rect 12670 7625 12698 7630
rect 12782 7657 12810 9198
rect 12838 8666 12866 10822
rect 13174 10850 13202 10855
rect 13174 10803 13202 10822
rect 13062 10793 13090 10799
rect 13062 10767 13063 10793
rect 13089 10767 13090 10793
rect 13006 9954 13034 9959
rect 13006 9907 13034 9926
rect 13062 9842 13090 10767
rect 13230 10794 13258 11943
rect 13398 11969 13426 12278
rect 14574 12306 14602 12311
rect 14798 12306 14826 12311
rect 14574 12259 14602 12278
rect 14742 12305 14826 12306
rect 14742 12279 14799 12305
rect 14825 12279 14826 12305
rect 14742 12278 14826 12279
rect 13398 11943 13399 11969
rect 13425 11943 13426 11969
rect 13398 11937 13426 11943
rect 13230 10761 13258 10766
rect 13286 11913 13314 11919
rect 13286 11887 13287 11913
rect 13313 11887 13314 11913
rect 13286 11410 13314 11887
rect 13454 11857 13482 11863
rect 13454 11831 13455 11857
rect 13481 11831 13482 11857
rect 13062 9617 13090 9814
rect 13062 9591 13063 9617
rect 13089 9591 13090 9617
rect 13062 9585 13090 9591
rect 13118 9562 13146 9567
rect 13118 9515 13146 9534
rect 13174 9505 13202 9511
rect 13174 9479 13175 9505
rect 13201 9479 13202 9505
rect 13174 8834 13202 9479
rect 13286 9506 13314 11382
rect 13342 11802 13370 11807
rect 13342 11577 13370 11774
rect 13342 11551 13343 11577
rect 13369 11551 13370 11577
rect 13342 10794 13370 11551
rect 13454 10906 13482 11831
rect 14742 11634 14770 12278
rect 14798 12273 14826 12278
rect 18830 12306 18858 12727
rect 20006 12474 20034 12783
rect 20006 12441 20034 12446
rect 18830 12273 18858 12278
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 15022 11634 15050 11639
rect 14742 11633 15050 11634
rect 14742 11607 15023 11633
rect 15049 11607 15050 11633
rect 14742 11606 15050 11607
rect 13734 11522 13762 11527
rect 13566 11521 13762 11522
rect 13566 11495 13735 11521
rect 13761 11495 13762 11521
rect 13566 11494 13762 11495
rect 13566 11241 13594 11494
rect 13734 11489 13762 11494
rect 14126 11522 14154 11527
rect 13566 11215 13567 11241
rect 13593 11215 13594 11241
rect 13566 11209 13594 11215
rect 13846 11186 13874 11191
rect 14014 11186 14042 11191
rect 13846 11185 14042 11186
rect 13846 11159 13847 11185
rect 13873 11159 14015 11185
rect 14041 11159 14042 11185
rect 13846 11158 14042 11159
rect 13846 11153 13874 11158
rect 14014 11153 14042 11158
rect 14126 11129 14154 11494
rect 14126 11103 14127 11129
rect 14153 11103 14154 11129
rect 14126 11097 14154 11103
rect 14182 11129 14210 11135
rect 14182 11103 14183 11129
rect 14209 11103 14210 11129
rect 13510 11074 13538 11079
rect 13510 11027 13538 11046
rect 13622 11073 13650 11079
rect 13622 11047 13623 11073
rect 13649 11047 13650 11073
rect 13454 10873 13482 10878
rect 13622 10850 13650 11047
rect 13398 10794 13426 10799
rect 13342 10793 13426 10794
rect 13342 10767 13399 10793
rect 13425 10767 13426 10793
rect 13342 10766 13426 10767
rect 13398 10457 13426 10766
rect 13398 10431 13399 10457
rect 13425 10431 13426 10457
rect 13398 10122 13426 10431
rect 13622 10402 13650 10822
rect 14182 10906 14210 11103
rect 13790 10738 13818 10743
rect 13790 10691 13818 10710
rect 13622 10369 13650 10374
rect 13342 9954 13370 9959
rect 13342 9617 13370 9926
rect 13342 9591 13343 9617
rect 13369 9591 13370 9617
rect 13342 9585 13370 9591
rect 13286 9478 13370 9506
rect 13286 9282 13314 9287
rect 13286 8889 13314 9254
rect 13286 8863 13287 8889
rect 13313 8863 13314 8889
rect 13286 8857 13314 8863
rect 13230 8834 13258 8839
rect 12894 8806 13230 8834
rect 12894 8777 12922 8806
rect 13230 8787 13258 8806
rect 13342 8833 13370 9478
rect 13342 8807 13343 8833
rect 13369 8807 13370 8833
rect 12894 8751 12895 8777
rect 12921 8751 12922 8777
rect 12894 8745 12922 8751
rect 13118 8722 13146 8727
rect 13118 8675 13146 8694
rect 13342 8666 13370 8807
rect 12838 8638 12922 8666
rect 12838 8554 12866 8559
rect 12838 8497 12866 8526
rect 12838 8471 12839 8497
rect 12865 8471 12866 8497
rect 12838 8465 12866 8471
rect 12838 8050 12866 8055
rect 12894 8050 12922 8638
rect 13174 8638 13370 8666
rect 13174 8610 13202 8638
rect 12950 8582 13202 8610
rect 12950 8441 12978 8582
rect 12950 8415 12951 8441
rect 12977 8415 12978 8441
rect 12950 8409 12978 8415
rect 13398 8441 13426 10094
rect 14182 10094 14210 10878
rect 14630 10738 14658 10743
rect 14294 10682 14322 10687
rect 14294 10121 14322 10654
rect 14574 10570 14602 10575
rect 14574 10401 14602 10542
rect 14630 10457 14658 10710
rect 14630 10431 14631 10457
rect 14657 10431 14658 10457
rect 14630 10425 14658 10431
rect 14574 10375 14575 10401
rect 14601 10375 14602 10401
rect 14574 10369 14602 10375
rect 14686 10402 14714 10407
rect 14686 10355 14714 10374
rect 14742 10290 14770 11606
rect 15022 11601 15050 11606
rect 18830 11578 18858 11583
rect 18830 11531 18858 11550
rect 14798 11522 14826 11527
rect 14798 11475 14826 11494
rect 20006 11466 20034 11471
rect 20006 11419 20034 11438
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 18830 11185 18858 11191
rect 18830 11159 18831 11185
rect 18857 11159 18858 11185
rect 14854 10738 14882 10743
rect 15078 10738 15106 10743
rect 14854 10691 14882 10710
rect 15022 10737 15106 10738
rect 15022 10711 15079 10737
rect 15105 10711 15106 10737
rect 15022 10710 15106 10711
rect 14686 10262 14770 10290
rect 14798 10289 14826 10295
rect 14798 10263 14799 10289
rect 14825 10263 14826 10289
rect 14294 10095 14295 10121
rect 14321 10095 14322 10121
rect 14182 10066 14266 10094
rect 14294 10089 14322 10095
rect 14574 10122 14602 10141
rect 14686 10122 14714 10262
rect 14602 10094 14714 10122
rect 14798 10094 14826 10263
rect 14574 10089 14602 10094
rect 14742 10066 14826 10094
rect 15022 10122 15050 10710
rect 15078 10705 15106 10710
rect 18830 10738 18858 11159
rect 20006 10794 20034 11215
rect 20006 10761 20034 10766
rect 18830 10705 18858 10710
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 14238 10065 14266 10066
rect 14238 10039 14239 10065
rect 14265 10039 14266 10065
rect 14238 10033 14266 10039
rect 14630 10038 14770 10066
rect 14406 10010 14434 10015
rect 14630 10010 14658 10038
rect 14406 10009 14658 10010
rect 14406 9983 14407 10009
rect 14433 9983 14658 10009
rect 14406 9982 14658 9983
rect 14406 9977 14434 9982
rect 14070 9954 14098 9959
rect 14070 9907 14098 9926
rect 13622 9338 13650 9343
rect 13622 9337 13930 9338
rect 13622 9311 13623 9337
rect 13649 9311 13930 9337
rect 13622 9310 13930 9311
rect 13622 9305 13650 9310
rect 13566 9282 13594 9287
rect 13566 9235 13594 9254
rect 13734 9225 13762 9231
rect 13734 9199 13735 9225
rect 13761 9199 13762 9225
rect 13734 8497 13762 9199
rect 13902 8945 13930 9310
rect 13902 8919 13903 8945
rect 13929 8919 13930 8945
rect 13902 8913 13930 8919
rect 13902 8834 13930 8839
rect 13734 8471 13735 8497
rect 13761 8471 13762 8497
rect 13734 8465 13762 8471
rect 13846 8778 13874 8783
rect 13398 8415 13399 8441
rect 13425 8415 13426 8441
rect 13398 8409 13426 8415
rect 13118 8330 13146 8335
rect 13118 8329 13258 8330
rect 13118 8303 13119 8329
rect 13145 8303 13258 8329
rect 13118 8302 13258 8303
rect 13118 8297 13146 8302
rect 12838 8049 13202 8050
rect 12838 8023 12839 8049
rect 12865 8023 13202 8049
rect 12838 8022 13202 8023
rect 12838 8017 12866 8022
rect 13174 7993 13202 8022
rect 13174 7967 13175 7993
rect 13201 7967 13202 7993
rect 13174 7961 13202 7967
rect 13230 7993 13258 8302
rect 13678 8050 13706 8055
rect 13846 8050 13874 8750
rect 13902 8777 13930 8806
rect 13902 8751 13903 8777
rect 13929 8751 13930 8777
rect 13902 8745 13930 8751
rect 15022 8554 15050 10094
rect 18830 10010 18858 10015
rect 18830 9963 18858 9982
rect 20006 9897 20034 9903
rect 20006 9871 20007 9897
rect 20033 9871 20034 9897
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 20006 9786 20034 9871
rect 20006 9753 20034 9758
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 13678 8049 13874 8050
rect 13678 8023 13679 8049
rect 13705 8023 13874 8049
rect 13678 8022 13874 8023
rect 14406 8553 15050 8554
rect 14406 8527 15023 8553
rect 15049 8527 15050 8553
rect 14406 8526 15050 8527
rect 13678 8017 13706 8022
rect 13230 7967 13231 7993
rect 13257 7967 13258 7993
rect 13230 7961 13258 7967
rect 13006 7937 13034 7943
rect 13006 7911 13007 7937
rect 13033 7911 13034 7937
rect 13006 7770 13034 7911
rect 13006 7737 13034 7742
rect 13062 7937 13090 7943
rect 13062 7911 13063 7937
rect 13089 7911 13090 7937
rect 13062 7714 13090 7911
rect 13118 7937 13146 7943
rect 13118 7911 13119 7937
rect 13145 7911 13146 7937
rect 13118 7770 13146 7911
rect 13510 7938 13538 7943
rect 13510 7891 13538 7910
rect 13622 7938 13650 7943
rect 13622 7891 13650 7910
rect 14182 7938 14210 7943
rect 13118 7737 13146 7742
rect 13062 7681 13090 7686
rect 12782 7631 12783 7657
rect 12809 7631 12810 7657
rect 11046 7322 11074 7327
rect 10990 7321 11074 7322
rect 10990 7295 11047 7321
rect 11073 7295 11074 7321
rect 10990 7294 11074 7295
rect 11046 7289 11074 7294
rect 11438 7322 11466 7518
rect 12334 7546 12362 7551
rect 12334 7499 12362 7518
rect 12726 7546 12754 7551
rect 11438 7289 11466 7294
rect 12110 7322 12138 7327
rect 12110 7275 12138 7294
rect 12726 7321 12754 7518
rect 12726 7295 12727 7321
rect 12753 7295 12754 7321
rect 12726 7289 12754 7295
rect 10710 7266 10738 7271
rect 12334 7266 12362 7271
rect 10710 7219 10738 7238
rect 12278 7238 12334 7266
rect 12278 6985 12306 7238
rect 12334 7219 12362 7238
rect 12782 7266 12810 7631
rect 13118 7658 13146 7663
rect 13118 7611 13146 7630
rect 13790 7658 13818 7663
rect 13790 7321 13818 7630
rect 14182 7601 14210 7910
rect 14406 7770 14434 8526
rect 15022 8521 15050 8526
rect 15078 8834 15106 8839
rect 15078 8442 15106 8806
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 14798 8414 15106 8442
rect 14798 8385 14826 8414
rect 14798 8359 14799 8385
rect 14825 8359 14826 8385
rect 14798 8353 14826 8359
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 20006 8105 20034 8111
rect 20006 8079 20007 8105
rect 20033 8079 20034 8105
rect 18830 8050 18858 8055
rect 18830 8003 18858 8022
rect 14182 7575 14183 7601
rect 14209 7575 14210 7601
rect 14182 7569 14210 7575
rect 14294 7769 14434 7770
rect 14294 7743 14407 7769
rect 14433 7743 14434 7769
rect 14294 7742 14434 7743
rect 14294 7546 14322 7742
rect 14406 7737 14434 7742
rect 20006 7770 20034 8079
rect 20006 7737 20034 7742
rect 18830 7658 18858 7663
rect 18830 7611 18858 7630
rect 14238 7518 14322 7546
rect 20006 7601 20034 7607
rect 20006 7575 20007 7601
rect 20033 7575 20034 7601
rect 14238 7490 14266 7518
rect 13790 7295 13791 7321
rect 13817 7295 13818 7321
rect 13790 7289 13818 7295
rect 14014 7462 14266 7490
rect 17598 7462 17730 7467
rect 14014 7321 14042 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 20006 7434 20034 7575
rect 20006 7401 20034 7406
rect 14014 7295 14015 7321
rect 14041 7295 14042 7321
rect 14014 7289 14042 7295
rect 12782 7233 12810 7238
rect 12278 6959 12279 6985
rect 12305 6959 12306 6985
rect 12278 6953 12306 6959
rect 10374 6818 10402 6823
rect 10094 6817 10402 6818
rect 10094 6791 10375 6817
rect 10401 6791 10402 6817
rect 10094 6790 10402 6791
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9086 5866 9170 5894
rect 8862 2170 8890 2175
rect 8694 2169 8890 2170
rect 8694 2143 8863 2169
rect 8889 2143 8890 2169
rect 8694 2142 8890 2143
rect 8862 2137 8890 2142
rect 8750 2058 8778 2063
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8750 400 8778 2030
rect 8974 1778 9002 1783
rect 9086 1778 9114 5866
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9366 2058 9394 2063
rect 9366 2011 9394 2030
rect 8974 1777 9114 1778
rect 8974 1751 8975 1777
rect 9001 1751 9114 1777
rect 8974 1750 9114 1751
rect 9310 1833 9338 1839
rect 9310 1807 9311 1833
rect 9337 1807 9338 1833
rect 8974 1745 9002 1750
rect 9310 1694 9338 1807
rect 10374 1777 10402 6790
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 10374 1751 10375 1777
rect 10401 1751 10402 1777
rect 10374 1745 10402 1751
rect 9086 1666 9338 1694
rect 10094 1722 10122 1727
rect 9086 400 9114 1666
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10094 400 10122 1694
rect 10878 1722 10906 1727
rect 10878 1665 10906 1694
rect 10878 1639 10879 1665
rect 10905 1639 10906 1665
rect 10878 1633 10906 1639
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 10080 0 10136 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 11438 19054 11466 19082
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 966 13118 994 13146
rect 2030 13062 2058 13090
rect 2086 13454 2114 13482
rect 966 12782 994 12810
rect 966 11774 994 11802
rect 966 11465 994 11466
rect 966 11439 967 11465
rect 967 11439 993 11465
rect 993 11439 994 11465
rect 966 11438 994 11439
rect 966 10766 994 10794
rect 966 10430 994 10458
rect 2142 13145 2170 13146
rect 2142 13119 2143 13145
rect 2143 13119 2169 13145
rect 2169 13119 2170 13145
rect 2142 13118 2170 13119
rect 5558 13118 5586 13146
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 6006 13089 6034 13090
rect 6006 13063 6007 13089
rect 6007 13063 6033 13089
rect 6033 13063 6034 13089
rect 6006 13062 6034 13063
rect 7686 13145 7714 13146
rect 7686 13119 7687 13145
rect 7687 13119 7713 13145
rect 7713 13119 7714 13145
rect 7686 13118 7714 13119
rect 6846 12782 6874 12810
rect 7238 13062 7266 13090
rect 5558 12726 5586 12754
rect 6902 12753 6930 12754
rect 6902 12727 6903 12753
rect 6903 12727 6929 12753
rect 6929 12727 6930 12753
rect 6902 12726 6930 12727
rect 6342 12697 6370 12698
rect 6342 12671 6343 12697
rect 6343 12671 6369 12697
rect 6369 12671 6370 12697
rect 6342 12670 6370 12671
rect 6846 12697 6874 12698
rect 6846 12671 6847 12697
rect 6847 12671 6873 12697
rect 6873 12671 6874 12697
rect 6846 12670 6874 12671
rect 6790 12614 6818 12642
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 2142 11969 2170 11970
rect 2142 11943 2143 11969
rect 2143 11943 2169 11969
rect 2169 11943 2170 11969
rect 2142 11942 2170 11943
rect 8078 13118 8106 13146
rect 7350 12782 7378 12810
rect 7518 12670 7546 12698
rect 7350 12641 7378 12642
rect 7350 12615 7351 12641
rect 7351 12615 7377 12641
rect 7377 12615 7378 12641
rect 7350 12614 7378 12615
rect 5166 11830 5194 11858
rect 2142 11577 2170 11578
rect 2142 11551 2143 11577
rect 2143 11551 2169 11577
rect 2169 11551 2170 11577
rect 2142 11550 2170 11551
rect 6622 11662 6650 11690
rect 5950 11550 5978 11578
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 2142 11185 2170 11186
rect 2142 11159 2143 11185
rect 2143 11159 2169 11185
rect 2169 11159 2170 11185
rect 2142 11158 2170 11159
rect 5838 11158 5866 11186
rect 2142 10793 2170 10794
rect 2142 10767 2143 10793
rect 2143 10767 2169 10793
rect 2169 10767 2170 10793
rect 2142 10766 2170 10767
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 2086 9982 2114 10010
rect 2142 10038 2170 10066
rect 5726 10038 5754 10066
rect 5726 9926 5754 9954
rect 6790 11857 6818 11858
rect 6790 11831 6791 11857
rect 6791 11831 6817 11857
rect 6817 11831 6818 11857
rect 6790 11830 6818 11831
rect 6846 11633 6874 11634
rect 6846 11607 6847 11633
rect 6847 11607 6873 11633
rect 6873 11607 6874 11633
rect 6846 11606 6874 11607
rect 6230 11438 6258 11466
rect 6846 11465 6874 11466
rect 6846 11439 6847 11465
rect 6847 11439 6873 11465
rect 6873 11439 6874 11465
rect 6846 11438 6874 11439
rect 6902 10513 6930 10514
rect 6902 10487 6903 10513
rect 6903 10487 6929 10513
rect 6929 10487 6930 10513
rect 6902 10486 6930 10487
rect 5838 10038 5866 10066
rect 7014 11270 7042 11298
rect 7126 11689 7154 11690
rect 7126 11663 7127 11689
rect 7127 11663 7153 11689
rect 7153 11663 7154 11689
rect 7126 11662 7154 11663
rect 7574 12558 7602 12586
rect 7686 12726 7714 12754
rect 8022 12558 8050 12586
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9702 13145 9730 13146
rect 9702 13119 9703 13145
rect 9703 13119 9729 13145
rect 9729 13119 9730 13145
rect 9702 13118 9730 13119
rect 10038 13118 10066 13146
rect 8134 12753 8162 12754
rect 8134 12727 8135 12753
rect 8135 12727 8161 12753
rect 8161 12727 8162 12753
rect 8134 12726 8162 12727
rect 9478 12641 9506 12642
rect 9478 12615 9479 12641
rect 9479 12615 9505 12641
rect 9505 12615 9506 12641
rect 9478 12614 9506 12615
rect 8414 11830 8442 11858
rect 8022 11774 8050 11802
rect 8806 11774 8834 11802
rect 7574 11633 7602 11634
rect 7574 11607 7575 11633
rect 7575 11607 7601 11633
rect 7601 11607 7602 11633
rect 7574 11606 7602 11607
rect 7798 11606 7826 11634
rect 7462 11577 7490 11578
rect 7462 11551 7463 11577
rect 7463 11551 7489 11577
rect 7489 11551 7490 11577
rect 7462 11550 7490 11551
rect 7126 10878 7154 10906
rect 7406 10878 7434 10906
rect 7014 10598 7042 10626
rect 7126 10401 7154 10402
rect 7126 10375 7127 10401
rect 7127 10375 7153 10401
rect 7153 10375 7154 10401
rect 7126 10374 7154 10375
rect 966 9897 994 9898
rect 966 9871 967 9897
rect 967 9871 993 9897
rect 993 9871 994 9897
rect 966 9870 994 9871
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 6454 9478 6482 9506
rect 2142 9225 2170 9226
rect 2142 9199 2143 9225
rect 2143 9199 2169 9225
rect 2169 9199 2170 9225
rect 2142 9198 2170 9199
rect 5894 9198 5922 9226
rect 5390 9169 5418 9170
rect 5390 9143 5391 9169
rect 5391 9143 5417 9169
rect 5417 9143 5418 9169
rect 5390 9142 5418 9143
rect 966 9113 994 9114
rect 966 9087 967 9113
rect 967 9087 993 9113
rect 993 9087 994 9113
rect 966 9086 994 9087
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 966 8889 994 8890
rect 966 8863 967 8889
rect 967 8863 993 8889
rect 993 8863 994 8889
rect 966 8862 994 8863
rect 2142 8833 2170 8834
rect 2142 8807 2143 8833
rect 2143 8807 2169 8833
rect 2169 8807 2170 8833
rect 2142 8806 2170 8807
rect 5390 8750 5418 8778
rect 6902 9505 6930 9506
rect 6902 9479 6903 9505
rect 6903 9479 6929 9505
rect 6929 9479 6930 9505
rect 6902 9478 6930 9479
rect 7406 10654 7434 10682
rect 7462 10486 7490 10514
rect 7518 10766 7546 10794
rect 7462 10374 7490 10402
rect 7966 11185 7994 11186
rect 7966 11159 7967 11185
rect 7967 11159 7993 11185
rect 7993 11159 7994 11185
rect 7966 11158 7994 11159
rect 7630 10905 7658 10906
rect 7630 10879 7631 10905
rect 7631 10879 7657 10905
rect 7657 10879 7658 10905
rect 7630 10878 7658 10879
rect 7910 10822 7938 10850
rect 7630 10598 7658 10626
rect 7350 10094 7378 10122
rect 7238 10038 7266 10066
rect 7574 10345 7602 10346
rect 7574 10319 7575 10345
rect 7575 10319 7601 10345
rect 7601 10319 7602 10345
rect 7574 10318 7602 10319
rect 8694 10849 8722 10850
rect 8694 10823 8695 10849
rect 8695 10823 8721 10849
rect 8721 10823 8722 10849
rect 8694 10822 8722 10823
rect 7910 10318 7938 10346
rect 8526 10710 8554 10738
rect 7854 10121 7882 10122
rect 7854 10095 7855 10121
rect 7855 10095 7881 10121
rect 7881 10095 7882 10121
rect 7854 10094 7882 10095
rect 6790 9254 6818 9282
rect 6958 9142 6986 9170
rect 7182 9702 7210 9730
rect 7630 10065 7658 10066
rect 7630 10039 7631 10065
rect 7631 10039 7657 10065
rect 7657 10039 7658 10065
rect 7630 10038 7658 10039
rect 7742 9870 7770 9898
rect 7686 9281 7714 9282
rect 7686 9255 7687 9281
rect 7687 9255 7713 9281
rect 7713 9255 7714 9281
rect 7686 9254 7714 9255
rect 7294 9225 7322 9226
rect 7294 9199 7295 9225
rect 7295 9199 7321 9225
rect 7321 9199 7322 9225
rect 7294 9198 7322 9199
rect 5894 8806 5922 8834
rect 6790 8777 6818 8778
rect 6790 8751 6791 8777
rect 6791 8751 6817 8777
rect 6817 8751 6818 8777
rect 6790 8750 6818 8751
rect 7854 9254 7882 9282
rect 7126 8302 7154 8330
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 8302 8974 8330 9002
rect 8750 10654 8778 10682
rect 9478 12025 9506 12026
rect 9478 11999 9479 12025
rect 9479 11999 9505 12025
rect 9505 11999 9506 12025
rect 9478 11998 9506 11999
rect 9422 11438 9450 11466
rect 10878 13062 10906 13090
rect 10598 12726 10626 12754
rect 10430 12670 10458 12698
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9870 12417 9898 12418
rect 9870 12391 9871 12417
rect 9871 12391 9897 12417
rect 9897 12391 9898 12417
rect 9870 12390 9898 12391
rect 8638 10150 8666 10178
rect 8862 10905 8890 10906
rect 8862 10879 8863 10905
rect 8863 10879 8889 10905
rect 8889 10879 8890 10905
rect 8862 10878 8890 10879
rect 8862 10430 8890 10458
rect 8974 9870 9002 9898
rect 9198 10793 9226 10794
rect 9198 10767 9199 10793
rect 9199 10767 9225 10793
rect 9225 10767 9226 10793
rect 9198 10766 9226 10767
rect 9366 10710 9394 10738
rect 9534 10878 9562 10906
rect 9086 10598 9114 10626
rect 9086 10150 9114 10178
rect 9142 10094 9170 10122
rect 8694 8974 8722 9002
rect 9086 9534 9114 9562
rect 8302 8553 8330 8554
rect 8302 8527 8303 8553
rect 8303 8527 8329 8553
rect 8329 8527 8330 8553
rect 8302 8526 8330 8527
rect 8694 8526 8722 8554
rect 8414 8246 8442 8274
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 9646 11857 9674 11858
rect 9646 11831 9647 11857
rect 9647 11831 9673 11857
rect 9673 11831 9674 11857
rect 9646 11830 9674 11831
rect 10038 12025 10066 12026
rect 10038 11999 10039 12025
rect 10039 11999 10065 12025
rect 10065 11999 10066 12025
rect 10038 11998 10066 11999
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 9702 11382 9730 11410
rect 9926 11438 9954 11466
rect 9758 11297 9786 11298
rect 9758 11271 9759 11297
rect 9759 11271 9785 11297
rect 9785 11271 9786 11297
rect 9758 11270 9786 11271
rect 9702 11158 9730 11186
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 9646 10710 9674 10738
rect 10038 10822 10066 10850
rect 9534 10681 9562 10682
rect 9534 10655 9535 10681
rect 9535 10655 9561 10681
rect 9561 10655 9562 10681
rect 9534 10654 9562 10655
rect 10262 10793 10290 10794
rect 10262 10767 10263 10793
rect 10263 10767 10289 10793
rect 10289 10767 10290 10793
rect 10262 10766 10290 10767
rect 10094 10710 10122 10738
rect 10206 10542 10234 10570
rect 10038 10401 10066 10402
rect 10038 10375 10039 10401
rect 10039 10375 10065 10401
rect 10065 10375 10066 10401
rect 10038 10374 10066 10375
rect 9814 10262 9842 10290
rect 9702 10009 9730 10010
rect 9702 9983 9703 10009
rect 9703 9983 9729 10009
rect 9729 9983 9730 10009
rect 9702 9982 9730 9983
rect 9534 9897 9562 9898
rect 9534 9871 9535 9897
rect 9535 9871 9561 9897
rect 9561 9871 9562 9897
rect 9534 9870 9562 9871
rect 9534 9561 9562 9562
rect 9534 9535 9535 9561
rect 9535 9535 9561 9561
rect 9561 9535 9562 9561
rect 9534 9534 9562 9535
rect 9702 9814 9730 9842
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 10094 9870 10122 9898
rect 9982 9702 10010 9730
rect 10038 9478 10066 9506
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9422 9254 9450 9282
rect 8918 8414 8946 8442
rect 8974 8246 9002 8274
rect 8862 7686 8890 7714
rect 7686 7630 7714 7658
rect 8918 7657 8946 7658
rect 8918 7631 8919 7657
rect 8919 7631 8945 7657
rect 8945 7631 8946 7657
rect 8918 7630 8946 7631
rect 9254 8105 9282 8106
rect 9254 8079 9255 8105
rect 9255 8079 9281 8105
rect 9281 8079 9282 8105
rect 9254 8078 9282 8079
rect 9198 7713 9226 7714
rect 9198 7687 9199 7713
rect 9199 7687 9225 7713
rect 9225 7687 9226 7713
rect 9198 7686 9226 7687
rect 9646 9142 9674 9170
rect 10766 12753 10794 12754
rect 10766 12727 10767 12753
rect 10767 12727 10793 12753
rect 10793 12727 10794 12753
rect 10766 12726 10794 12727
rect 10654 12697 10682 12698
rect 10654 12671 10655 12697
rect 10655 12671 10681 12697
rect 10681 12671 10682 12697
rect 10654 12670 10682 12671
rect 10486 12390 10514 12418
rect 11158 13089 11186 13090
rect 11158 13063 11159 13089
rect 11159 13063 11185 13089
rect 11185 13063 11186 13089
rect 11158 13062 11186 13063
rect 11662 12809 11690 12810
rect 11662 12783 11663 12809
rect 11663 12783 11689 12809
rect 11689 12783 11690 12809
rect 11662 12782 11690 12783
rect 12110 12809 12138 12810
rect 12110 12783 12111 12809
rect 12111 12783 12137 12809
rect 12137 12783 12138 12809
rect 12110 12782 12138 12783
rect 10990 12334 11018 12362
rect 11606 12614 11634 12642
rect 10598 11158 10626 11186
rect 11438 12446 11466 12474
rect 11214 11662 11242 11690
rect 11550 12390 11578 12418
rect 11382 11718 11410 11746
rect 11494 11718 11522 11746
rect 11270 11606 11298 11634
rect 11326 11662 11354 11690
rect 11550 11606 11578 11634
rect 11382 11577 11410 11578
rect 11382 11551 11383 11577
rect 11383 11551 11409 11577
rect 11409 11551 11410 11577
rect 11382 11550 11410 11551
rect 11214 11185 11242 11186
rect 11214 11159 11215 11185
rect 11215 11159 11241 11185
rect 11241 11159 11242 11185
rect 11214 11158 11242 11159
rect 10934 10878 10962 10906
rect 11046 11102 11074 11130
rect 10318 10094 10346 10122
rect 10710 10766 10738 10794
rect 10766 10654 10794 10682
rect 10990 10654 11018 10682
rect 10654 10262 10682 10290
rect 10934 9814 10962 9842
rect 10990 10094 11018 10122
rect 10598 9590 10626 9618
rect 10374 9505 10402 9506
rect 10374 9479 10375 9505
rect 10375 9479 10401 9505
rect 10401 9479 10402 9505
rect 10374 9478 10402 9479
rect 10318 9086 10346 9114
rect 9758 8974 9786 9002
rect 9646 8750 9674 8778
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 10206 8833 10234 8834
rect 10206 8807 10207 8833
rect 10207 8807 10233 8833
rect 10233 8807 10234 8833
rect 10206 8806 10234 8807
rect 10654 8806 10682 8834
rect 11214 10262 11242 10290
rect 11158 9870 11186 9898
rect 11214 10094 11242 10122
rect 11158 9617 11186 9618
rect 11158 9591 11159 9617
rect 11159 9591 11185 9617
rect 11185 9591 11186 9617
rect 11158 9590 11186 9591
rect 11102 9478 11130 9506
rect 10878 9198 10906 9226
rect 10934 9254 10962 9282
rect 10822 9086 10850 9114
rect 10710 8750 10738 8778
rect 10878 9030 10906 9058
rect 9982 8385 10010 8386
rect 9982 8359 9983 8385
rect 9983 8359 10009 8385
rect 10009 8359 10010 8385
rect 9982 8358 10010 8359
rect 9366 8078 9394 8106
rect 9702 8302 9730 8330
rect 9310 7686 9338 7714
rect 9142 7630 9170 7658
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 9030 7462 9058 7490
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 10654 8553 10682 8554
rect 10654 8527 10655 8553
rect 10655 8527 10681 8553
rect 10681 8527 10682 8553
rect 10654 8526 10682 8527
rect 10542 8385 10570 8386
rect 10542 8359 10543 8385
rect 10543 8359 10569 8385
rect 10569 8359 10570 8385
rect 10542 8358 10570 8359
rect 10598 8302 10626 8330
rect 11158 9225 11186 9226
rect 11158 9199 11159 9225
rect 11159 9199 11185 9225
rect 11185 9199 11186 9225
rect 11158 9198 11186 9199
rect 11662 11718 11690 11746
rect 11494 11270 11522 11298
rect 11382 11185 11410 11186
rect 11382 11159 11383 11185
rect 11383 11159 11409 11185
rect 11409 11159 11410 11185
rect 11382 11158 11410 11159
rect 11606 11073 11634 11074
rect 11606 11047 11607 11073
rect 11607 11047 11633 11073
rect 11633 11047 11634 11073
rect 11606 11046 11634 11047
rect 11438 10905 11466 10906
rect 11438 10879 11439 10905
rect 11439 10879 11465 10905
rect 11465 10879 11466 10905
rect 11438 10878 11466 10879
rect 11382 10822 11410 10850
rect 11326 10430 11354 10458
rect 11774 12726 11802 12754
rect 12222 12753 12250 12754
rect 12222 12727 12223 12753
rect 12223 12727 12249 12753
rect 12249 12727 12250 12753
rect 12222 12726 12250 12727
rect 12110 12446 12138 12474
rect 12054 12390 12082 12418
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 12782 19110 12810 19138
rect 14686 19137 14714 19138
rect 14686 19111 14687 19137
rect 14687 19111 14713 19137
rect 14713 19111 14714 19137
rect 14686 19110 14714 19111
rect 12838 19081 12866 19082
rect 12838 19055 12839 19081
rect 12839 19055 12865 19081
rect 12865 19055 12866 19081
rect 12838 19054 12866 19055
rect 12446 18718 12474 18746
rect 13118 18745 13146 18746
rect 13118 18719 13119 18745
rect 13119 18719 13145 18745
rect 13145 18719 13146 18745
rect 13118 18718 13146 18719
rect 12334 13118 12362 13146
rect 12782 13257 12810 13258
rect 12782 13231 12783 13257
rect 12783 13231 12809 13257
rect 12809 13231 12810 13257
rect 12782 13230 12810 13231
rect 12670 13145 12698 13146
rect 12670 13119 12671 13145
rect 12671 13119 12697 13145
rect 12697 13119 12698 13145
rect 12670 13118 12698 13119
rect 12670 12361 12698 12362
rect 12670 12335 12671 12361
rect 12671 12335 12697 12361
rect 12697 12335 12698 12361
rect 12670 12334 12698 12335
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 20118 17822 20146 17850
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 14294 13230 14322 13258
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 13118 12361 13146 12362
rect 13118 12335 13119 12361
rect 13119 12335 13145 12361
rect 13145 12335 13146 12361
rect 13118 12334 13146 12335
rect 13398 12278 13426 12306
rect 13118 11774 13146 11802
rect 11830 11662 11858 11690
rect 11830 11270 11858 11298
rect 12110 11297 12138 11298
rect 12110 11271 12111 11297
rect 12111 11271 12137 11297
rect 12137 11271 12138 11297
rect 12110 11270 12138 11271
rect 11718 11102 11746 11130
rect 11942 11158 11970 11186
rect 12222 11158 12250 11186
rect 11438 10486 11466 10514
rect 11774 10486 11802 10514
rect 11270 9702 11298 9730
rect 11382 10289 11410 10290
rect 11382 10263 11383 10289
rect 11383 10263 11409 10289
rect 11409 10263 11410 10289
rect 11382 10262 11410 10263
rect 11270 9422 11298 9450
rect 11494 9870 11522 9898
rect 11886 10766 11914 10794
rect 11886 10430 11914 10458
rect 11662 10401 11690 10402
rect 11662 10375 11663 10401
rect 11663 10375 11689 10401
rect 11689 10375 11690 10401
rect 11662 10374 11690 10375
rect 12278 9926 12306 9954
rect 11662 9814 11690 9842
rect 11718 9590 11746 9618
rect 11606 9422 11634 9450
rect 11270 9030 11298 9058
rect 10206 7769 10234 7770
rect 10206 7743 10207 7769
rect 10207 7743 10233 7769
rect 10233 7743 10234 7769
rect 10206 7742 10234 7743
rect 9926 7686 9954 7714
rect 9814 7574 9842 7602
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 10150 7601 10178 7602
rect 10150 7575 10151 7601
rect 10151 7575 10177 7601
rect 10177 7575 10178 7601
rect 10150 7574 10178 7575
rect 11550 9225 11578 9226
rect 11550 9199 11551 9225
rect 11551 9199 11577 9225
rect 11577 9199 11578 9225
rect 11550 9198 11578 9199
rect 12838 10822 12866 10850
rect 12670 10094 12698 10122
rect 12222 9534 12250 9562
rect 12054 9422 12082 9450
rect 11774 9281 11802 9282
rect 11774 9255 11775 9281
rect 11775 9255 11801 9281
rect 11801 9255 11802 9281
rect 11774 9254 11802 9255
rect 12110 9225 12138 9226
rect 12110 9199 12111 9225
rect 12111 9199 12137 9225
rect 12137 9199 12138 9225
rect 12110 9198 12138 9199
rect 12670 9198 12698 9226
rect 11886 9113 11914 9114
rect 11886 9087 11887 9113
rect 11887 9087 11913 9113
rect 11913 9087 11914 9113
rect 11886 9086 11914 9087
rect 11886 8694 11914 8722
rect 11382 8553 11410 8554
rect 11382 8527 11383 8553
rect 11383 8527 11409 8553
rect 11409 8527 11410 8553
rect 11382 8526 11410 8527
rect 12726 8526 12754 8554
rect 11214 8358 11242 8386
rect 12502 8358 12530 8386
rect 11774 7769 11802 7770
rect 11774 7743 11775 7769
rect 11775 7743 11801 7769
rect 11801 7743 11802 7769
rect 11774 7742 11802 7743
rect 12614 7742 12642 7770
rect 12278 7713 12306 7714
rect 12278 7687 12279 7713
rect 12279 7687 12305 7713
rect 12305 7687 12306 7713
rect 12278 7686 12306 7687
rect 11046 7518 11074 7546
rect 12726 7937 12754 7938
rect 12726 7911 12727 7937
rect 12727 7911 12753 7937
rect 12753 7911 12754 7937
rect 12726 7910 12754 7911
rect 12670 7630 12698 7658
rect 13174 10849 13202 10850
rect 13174 10823 13175 10849
rect 13175 10823 13201 10849
rect 13201 10823 13202 10849
rect 13174 10822 13202 10823
rect 13006 9953 13034 9954
rect 13006 9927 13007 9953
rect 13007 9927 13033 9953
rect 13033 9927 13034 9953
rect 13006 9926 13034 9927
rect 14574 12305 14602 12306
rect 14574 12279 14575 12305
rect 14575 12279 14601 12305
rect 14601 12279 14602 12305
rect 14574 12278 14602 12279
rect 13230 10766 13258 10794
rect 13286 11382 13314 11410
rect 13062 9814 13090 9842
rect 13118 9561 13146 9562
rect 13118 9535 13119 9561
rect 13119 9535 13145 9561
rect 13145 9535 13146 9561
rect 13118 9534 13146 9535
rect 13342 11774 13370 11802
rect 20006 12446 20034 12474
rect 18830 12278 18858 12306
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 14126 11494 14154 11522
rect 13510 11073 13538 11074
rect 13510 11047 13511 11073
rect 13511 11047 13537 11073
rect 13537 11047 13538 11073
rect 13510 11046 13538 11047
rect 13454 10878 13482 10906
rect 13622 10822 13650 10850
rect 14182 10878 14210 10906
rect 13790 10737 13818 10738
rect 13790 10711 13791 10737
rect 13791 10711 13817 10737
rect 13817 10711 13818 10737
rect 13790 10710 13818 10711
rect 13622 10374 13650 10402
rect 13398 10094 13426 10122
rect 13342 9926 13370 9954
rect 13286 9254 13314 9282
rect 13230 8833 13258 8834
rect 13230 8807 13231 8833
rect 13231 8807 13257 8833
rect 13257 8807 13258 8833
rect 13230 8806 13258 8807
rect 13118 8721 13146 8722
rect 13118 8695 13119 8721
rect 13119 8695 13145 8721
rect 13145 8695 13146 8721
rect 13118 8694 13146 8695
rect 12838 8526 12866 8554
rect 14630 10710 14658 10738
rect 14294 10654 14322 10682
rect 14574 10542 14602 10570
rect 14686 10401 14714 10402
rect 14686 10375 14687 10401
rect 14687 10375 14713 10401
rect 14713 10375 14714 10401
rect 14686 10374 14714 10375
rect 18830 11577 18858 11578
rect 18830 11551 18831 11577
rect 18831 11551 18857 11577
rect 18857 11551 18858 11577
rect 18830 11550 18858 11551
rect 14798 11521 14826 11522
rect 14798 11495 14799 11521
rect 14799 11495 14825 11521
rect 14825 11495 14826 11521
rect 14798 11494 14826 11495
rect 20006 11465 20034 11466
rect 20006 11439 20007 11465
rect 20007 11439 20033 11465
rect 20033 11439 20034 11465
rect 20006 11438 20034 11439
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 14854 10737 14882 10738
rect 14854 10711 14855 10737
rect 14855 10711 14881 10737
rect 14881 10711 14882 10737
rect 14854 10710 14882 10711
rect 14574 10121 14602 10122
rect 14574 10095 14575 10121
rect 14575 10095 14601 10121
rect 14601 10095 14602 10121
rect 14574 10094 14602 10095
rect 20006 10766 20034 10794
rect 18830 10710 18858 10738
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 15022 10094 15050 10122
rect 14070 9953 14098 9954
rect 14070 9927 14071 9953
rect 14071 9927 14097 9953
rect 14097 9927 14098 9953
rect 14070 9926 14098 9927
rect 13566 9281 13594 9282
rect 13566 9255 13567 9281
rect 13567 9255 13593 9281
rect 13593 9255 13594 9281
rect 13566 9254 13594 9255
rect 13902 8806 13930 8834
rect 13846 8777 13874 8778
rect 13846 8751 13847 8777
rect 13847 8751 13873 8777
rect 13873 8751 13874 8777
rect 13846 8750 13874 8751
rect 18830 10009 18858 10010
rect 18830 9983 18831 10009
rect 18831 9983 18857 10009
rect 18857 9983 18858 10009
rect 18830 9982 18858 9983
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 20006 9758 20034 9786
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 13006 7742 13034 7770
rect 13510 7937 13538 7938
rect 13510 7911 13511 7937
rect 13511 7911 13537 7937
rect 13537 7911 13538 7937
rect 13510 7910 13538 7911
rect 13622 7937 13650 7938
rect 13622 7911 13623 7937
rect 13623 7911 13649 7937
rect 13649 7911 13650 7937
rect 13622 7910 13650 7911
rect 14182 7910 14210 7938
rect 13118 7742 13146 7770
rect 13062 7686 13090 7714
rect 11438 7518 11466 7546
rect 12334 7545 12362 7546
rect 12334 7519 12335 7545
rect 12335 7519 12361 7545
rect 12361 7519 12362 7545
rect 12334 7518 12362 7519
rect 12726 7518 12754 7546
rect 11438 7294 11466 7322
rect 12110 7321 12138 7322
rect 12110 7295 12111 7321
rect 12111 7295 12137 7321
rect 12137 7295 12138 7321
rect 12110 7294 12138 7295
rect 10710 7265 10738 7266
rect 10710 7239 10711 7265
rect 10711 7239 10737 7265
rect 10737 7239 10738 7265
rect 10710 7238 10738 7239
rect 12334 7265 12362 7266
rect 12334 7239 12335 7265
rect 12335 7239 12361 7265
rect 12361 7239 12362 7265
rect 12334 7238 12362 7239
rect 13118 7657 13146 7658
rect 13118 7631 13119 7657
rect 13119 7631 13145 7657
rect 13145 7631 13146 7657
rect 13118 7630 13146 7631
rect 13790 7630 13818 7658
rect 15078 8806 15106 8834
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 20006 8750 20034 8778
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 18830 8049 18858 8050
rect 18830 8023 18831 8049
rect 18831 8023 18857 8049
rect 18857 8023 18858 8049
rect 18830 8022 18858 8023
rect 20006 7742 20034 7770
rect 18830 7657 18858 7658
rect 18830 7631 18831 7657
rect 18831 7631 18857 7657
rect 18857 7631 18858 7657
rect 18830 7630 18858 7631
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 20006 7406 20034 7434
rect 12782 7238 12810 7266
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 8750 2030 8778 2058
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9366 2057 9394 2058
rect 9366 2031 9367 2057
rect 9367 2031 9393 2057
rect 9393 2031 9394 2057
rect 9366 2030 9394 2031
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 10094 1694 10122 1722
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 10878 1694 10906 1722
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 12777 19110 12782 19138
rect 12810 19110 14686 19138
rect 14714 19110 14719 19138
rect 11433 19054 11438 19082
rect 11466 19054 12838 19082
rect 12866 19054 12871 19082
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 12441 18718 12446 18746
rect 12474 18718 13118 18746
rect 13146 18718 13151 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 20600 17850 21000 17864
rect 20113 17822 20118 17850
rect 20146 17822 21000 17850
rect 20600 17808 21000 17822
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 0 13482 400 13496
rect 0 13454 2086 13482
rect 2114 13454 2119 13482
rect 0 13440 400 13454
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 12777 13230 12782 13258
rect 12810 13230 14294 13258
rect 14322 13230 14327 13258
rect 0 13146 400 13160
rect 0 13118 966 13146
rect 994 13118 999 13146
rect 2137 13118 2142 13146
rect 2170 13118 5558 13146
rect 5586 13118 5591 13146
rect 7681 13118 7686 13146
rect 7714 13118 8078 13146
rect 8106 13118 9702 13146
rect 9730 13118 10038 13146
rect 10066 13118 10071 13146
rect 12329 13118 12334 13146
rect 12362 13118 12670 13146
rect 12698 13118 12703 13146
rect 0 13104 400 13118
rect 2025 13062 2030 13090
rect 2058 13062 6006 13090
rect 6034 13062 7238 13090
rect 7266 13062 7271 13090
rect 10873 13062 10878 13090
rect 10906 13062 11158 13090
rect 11186 13062 11191 13090
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 0 12810 400 12824
rect 0 12782 966 12810
rect 994 12782 999 12810
rect 6841 12782 6846 12810
rect 6874 12782 7350 12810
rect 7378 12782 7383 12810
rect 11657 12782 11662 12810
rect 11690 12782 12110 12810
rect 12138 12782 12143 12810
rect 0 12768 400 12782
rect 5553 12726 5558 12754
rect 5586 12726 6902 12754
rect 6930 12726 6935 12754
rect 7681 12726 7686 12754
rect 7714 12726 8134 12754
rect 8162 12726 10598 12754
rect 10626 12726 10766 12754
rect 10794 12726 10799 12754
rect 11769 12726 11774 12754
rect 11802 12726 12222 12754
rect 12250 12726 12255 12754
rect 6337 12670 6342 12698
rect 6370 12670 6846 12698
rect 6874 12670 6879 12698
rect 7513 12670 7518 12698
rect 7546 12670 10430 12698
rect 10458 12670 10654 12698
rect 10682 12670 10687 12698
rect 6785 12614 6790 12642
rect 6818 12614 7350 12642
rect 7378 12614 7383 12642
rect 9473 12614 9478 12642
rect 9506 12614 11606 12642
rect 11634 12614 11639 12642
rect 7569 12558 7574 12586
rect 7602 12558 8022 12586
rect 8050 12558 8055 12586
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 20600 12474 21000 12488
rect 11433 12446 11438 12474
rect 11466 12446 12110 12474
rect 12138 12446 12143 12474
rect 20001 12446 20006 12474
rect 20034 12446 21000 12474
rect 20600 12432 21000 12446
rect 9865 12390 9870 12418
rect 9898 12390 10486 12418
rect 10514 12390 11550 12418
rect 11578 12390 12054 12418
rect 12082 12390 12087 12418
rect 10985 12334 10990 12362
rect 11018 12334 12670 12362
rect 12698 12334 13118 12362
rect 13146 12334 13151 12362
rect 13393 12278 13398 12306
rect 13426 12278 14574 12306
rect 14602 12278 18830 12306
rect 18858 12278 18863 12306
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 9473 11998 9478 12026
rect 9506 11998 10038 12026
rect 10066 11998 10071 12026
rect 2137 11942 2142 11970
rect 2170 11942 4214 11970
rect 4186 11858 4214 11942
rect 4186 11830 5166 11858
rect 5194 11830 6790 11858
rect 6818 11830 6823 11858
rect 8409 11830 8414 11858
rect 8442 11830 9646 11858
rect 9674 11830 9679 11858
rect 0 11802 400 11816
rect 0 11774 966 11802
rect 994 11774 999 11802
rect 8017 11774 8022 11802
rect 8050 11774 8806 11802
rect 8834 11774 8839 11802
rect 13113 11774 13118 11802
rect 13146 11774 13342 11802
rect 13370 11774 13375 11802
rect 0 11760 400 11774
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 11363 11718 11382 11746
rect 11410 11718 11415 11746
rect 11489 11718 11494 11746
rect 11522 11718 11527 11746
rect 11657 11718 11662 11746
rect 11690 11718 11695 11746
rect 6617 11662 6622 11690
rect 6650 11662 7126 11690
rect 7154 11662 7159 11690
rect 11209 11662 11214 11690
rect 11242 11662 11326 11690
rect 11354 11662 11359 11690
rect 11494 11634 11522 11718
rect 11662 11690 11690 11718
rect 11662 11662 11830 11690
rect 11858 11662 11863 11690
rect 6841 11606 6846 11634
rect 6874 11606 7574 11634
rect 7602 11606 7798 11634
rect 7826 11606 7831 11634
rect 11265 11606 11270 11634
rect 11298 11606 11303 11634
rect 11494 11606 11550 11634
rect 11578 11606 11583 11634
rect 11270 11578 11298 11606
rect 2137 11550 2142 11578
rect 2170 11550 5950 11578
rect 5978 11550 7462 11578
rect 7490 11550 7495 11578
rect 11270 11550 11382 11578
rect 11410 11550 11415 11578
rect 15946 11550 18830 11578
rect 18858 11550 18863 11578
rect 15946 11522 15974 11550
rect 14121 11494 14126 11522
rect 14154 11494 14798 11522
rect 14826 11494 15974 11522
rect 0 11466 400 11480
rect 20600 11466 21000 11480
rect 0 11438 966 11466
rect 994 11438 999 11466
rect 6225 11438 6230 11466
rect 6258 11438 6846 11466
rect 6874 11438 6879 11466
rect 9417 11438 9422 11466
rect 9450 11438 9926 11466
rect 9954 11438 9959 11466
rect 20001 11438 20006 11466
rect 20034 11438 21000 11466
rect 0 11424 400 11438
rect 20600 11424 21000 11438
rect 9697 11382 9702 11410
rect 9730 11382 13286 11410
rect 13314 11382 13319 11410
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 7009 11270 7014 11298
rect 7042 11270 9758 11298
rect 9786 11270 11494 11298
rect 11522 11270 11830 11298
rect 11858 11270 12110 11298
rect 12138 11270 12143 11298
rect 2137 11158 2142 11186
rect 2170 11158 5838 11186
rect 5866 11158 5871 11186
rect 7961 11158 7966 11186
rect 7994 11158 9702 11186
rect 9730 11158 9735 11186
rect 10593 11158 10598 11186
rect 10626 11158 11214 11186
rect 11242 11158 11247 11186
rect 11363 11158 11382 11186
rect 11410 11158 11942 11186
rect 11970 11158 12222 11186
rect 12250 11158 12255 11186
rect 11041 11102 11046 11130
rect 11074 11102 11718 11130
rect 11746 11102 11751 11130
rect 11601 11046 11606 11074
rect 11634 11046 13510 11074
rect 13538 11046 13543 11074
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 7121 10878 7126 10906
rect 7154 10878 7406 10906
rect 7434 10878 7630 10906
rect 7658 10878 7663 10906
rect 8857 10878 8862 10906
rect 8890 10878 9534 10906
rect 9562 10878 9567 10906
rect 10929 10878 10934 10906
rect 10962 10878 11438 10906
rect 11466 10878 13454 10906
rect 13482 10878 14182 10906
rect 14210 10878 14215 10906
rect 7905 10822 7910 10850
rect 7938 10822 8694 10850
rect 8722 10822 8727 10850
rect 10033 10822 10038 10850
rect 10066 10822 11382 10850
rect 11410 10822 11415 10850
rect 12833 10822 12838 10850
rect 12866 10822 13174 10850
rect 13202 10822 13622 10850
rect 13650 10822 13655 10850
rect 0 10794 400 10808
rect 20600 10794 21000 10808
rect 0 10766 966 10794
rect 994 10766 999 10794
rect 2137 10766 2142 10794
rect 2170 10766 7518 10794
rect 7546 10766 7551 10794
rect 9193 10766 9198 10794
rect 9226 10766 10262 10794
rect 10290 10766 10710 10794
rect 10738 10766 10743 10794
rect 11881 10766 11886 10794
rect 11914 10766 13230 10794
rect 13258 10766 13263 10794
rect 20001 10766 20006 10794
rect 20034 10766 21000 10794
rect 0 10752 400 10766
rect 20600 10752 21000 10766
rect 8521 10710 8526 10738
rect 8554 10710 9366 10738
rect 9394 10710 9646 10738
rect 9674 10710 10094 10738
rect 10122 10710 10127 10738
rect 13785 10710 13790 10738
rect 13818 10710 14630 10738
rect 14658 10710 14663 10738
rect 14849 10710 14854 10738
rect 14882 10710 18830 10738
rect 18858 10710 18863 10738
rect 14854 10682 14882 10710
rect 7401 10654 7406 10682
rect 7434 10654 8750 10682
rect 8778 10654 9534 10682
rect 9562 10654 10766 10682
rect 10794 10654 10990 10682
rect 11018 10654 11023 10682
rect 14289 10654 14294 10682
rect 14322 10654 14882 10682
rect 7009 10598 7014 10626
rect 7042 10598 7630 10626
rect 7658 10598 9086 10626
rect 9114 10598 9119 10626
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 10201 10542 10206 10570
rect 10234 10542 14574 10570
rect 14602 10542 14607 10570
rect 6897 10486 6902 10514
rect 6930 10486 7462 10514
rect 7490 10486 7495 10514
rect 11433 10486 11438 10514
rect 11466 10486 11774 10514
rect 11802 10486 11807 10514
rect 0 10458 400 10472
rect 0 10430 966 10458
rect 994 10430 999 10458
rect 8857 10430 8862 10458
rect 8890 10430 11326 10458
rect 11354 10430 11886 10458
rect 11914 10430 11919 10458
rect 0 10416 400 10430
rect 7121 10374 7126 10402
rect 7154 10374 7462 10402
rect 7490 10374 7495 10402
rect 10033 10374 10038 10402
rect 10066 10374 11662 10402
rect 11690 10374 11695 10402
rect 13617 10374 13622 10402
rect 13650 10374 14686 10402
rect 14714 10374 14719 10402
rect 7569 10318 7574 10346
rect 7602 10318 7910 10346
rect 7938 10318 7943 10346
rect 9809 10262 9814 10290
rect 9842 10262 10654 10290
rect 10682 10262 11214 10290
rect 11242 10262 11382 10290
rect 11410 10262 11415 10290
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 8633 10150 8638 10178
rect 8666 10150 9086 10178
rect 9114 10150 9119 10178
rect 7345 10094 7350 10122
rect 7378 10094 7854 10122
rect 7882 10094 9142 10122
rect 9170 10094 9175 10122
rect 10313 10094 10318 10122
rect 10346 10094 10990 10122
rect 11018 10094 11214 10122
rect 11242 10094 11247 10122
rect 12665 10094 12670 10122
rect 12698 10094 13398 10122
rect 13426 10094 14574 10122
rect 14602 10094 15022 10122
rect 15050 10094 15055 10122
rect 2137 10038 2142 10066
rect 2170 10038 5726 10066
rect 5754 10038 5759 10066
rect 5833 10038 5838 10066
rect 5866 10038 7238 10066
rect 7266 10038 7630 10066
rect 7658 10038 7663 10066
rect 2081 9982 2086 10010
rect 2114 9982 9702 10010
rect 9730 9982 9735 10010
rect 15946 9982 18830 10010
rect 18858 9982 18863 10010
rect 15946 9954 15974 9982
rect 5721 9926 5726 9954
rect 5754 9926 7574 9954
rect 12273 9926 12278 9954
rect 12306 9926 13006 9954
rect 13034 9926 13039 9954
rect 13337 9926 13342 9954
rect 13370 9926 14070 9954
rect 14098 9926 15974 9954
rect 7546 9898 7574 9926
rect 961 9870 966 9898
rect 994 9870 999 9898
rect 7546 9870 7742 9898
rect 7770 9870 8974 9898
rect 9002 9870 9007 9898
rect 9529 9870 9534 9898
rect 9562 9870 10094 9898
rect 10122 9870 11158 9898
rect 11186 9870 11494 9898
rect 11522 9870 11527 9898
rect 0 9786 400 9800
rect 966 9786 994 9870
rect 9697 9814 9702 9842
rect 9730 9814 10934 9842
rect 10962 9814 11662 9842
rect 11690 9814 13062 9842
rect 13090 9814 13095 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 20600 9786 21000 9800
rect 0 9758 994 9786
rect 20001 9758 20006 9786
rect 20034 9758 21000 9786
rect 0 9744 400 9758
rect 20600 9744 21000 9758
rect 7177 9702 7182 9730
rect 7210 9702 9982 9730
rect 10010 9702 11270 9730
rect 11298 9702 11303 9730
rect 10593 9590 10598 9618
rect 10626 9590 11158 9618
rect 11186 9590 11718 9618
rect 11746 9590 11751 9618
rect 9081 9534 9086 9562
rect 9114 9534 9534 9562
rect 9562 9534 9567 9562
rect 12217 9534 12222 9562
rect 12250 9534 13118 9562
rect 13146 9534 13151 9562
rect 6449 9478 6454 9506
rect 6482 9478 6902 9506
rect 6930 9478 6935 9506
rect 10033 9478 10038 9506
rect 10066 9478 10374 9506
rect 10402 9478 11102 9506
rect 11130 9478 11135 9506
rect 11265 9422 11270 9450
rect 11298 9422 11606 9450
rect 11634 9422 12054 9450
rect 12082 9422 12087 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 6785 9254 6790 9282
rect 6818 9254 7686 9282
rect 7714 9254 7854 9282
rect 7882 9254 7887 9282
rect 9417 9254 9422 9282
rect 9450 9254 10934 9282
rect 10962 9254 11774 9282
rect 11802 9254 11807 9282
rect 13281 9254 13286 9282
rect 13314 9254 13566 9282
rect 13594 9254 13599 9282
rect 2137 9198 2142 9226
rect 2170 9198 4214 9226
rect 5889 9198 5894 9226
rect 5922 9198 7294 9226
rect 7322 9198 7327 9226
rect 10873 9198 10878 9226
rect 10906 9198 11158 9226
rect 11186 9198 11191 9226
rect 11545 9198 11550 9226
rect 11578 9198 12110 9226
rect 12138 9198 12670 9226
rect 12698 9198 12703 9226
rect 4186 9170 4214 9198
rect 4186 9142 5390 9170
rect 5418 9142 5423 9170
rect 6953 9142 6958 9170
rect 6986 9142 9646 9170
rect 9674 9142 9679 9170
rect 0 9114 400 9128
rect 0 9086 966 9114
rect 994 9086 999 9114
rect 10313 9086 10318 9114
rect 10346 9086 10822 9114
rect 10850 9086 11886 9114
rect 11914 9086 11919 9114
rect 0 9072 400 9086
rect 10873 9030 10878 9058
rect 10906 9030 11270 9058
rect 11298 9030 11303 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 8297 8974 8302 9002
rect 8330 8974 8694 9002
rect 8722 8974 9758 9002
rect 9786 8974 9791 9002
rect 961 8862 966 8890
rect 994 8862 999 8890
rect 0 8778 400 8792
rect 966 8778 994 8862
rect 2137 8806 2142 8834
rect 2170 8806 5894 8834
rect 5922 8806 5927 8834
rect 10201 8806 10206 8834
rect 10234 8806 10654 8834
rect 10682 8806 10687 8834
rect 13225 8806 13230 8834
rect 13258 8806 13454 8834
rect 13897 8806 13902 8834
rect 13930 8806 15078 8834
rect 15106 8806 18830 8834
rect 18858 8806 18863 8834
rect 13426 8778 13454 8806
rect 20600 8778 21000 8792
rect 0 8750 994 8778
rect 5385 8750 5390 8778
rect 5418 8750 6790 8778
rect 6818 8750 6823 8778
rect 9641 8750 9646 8778
rect 9674 8750 10710 8778
rect 10738 8750 10743 8778
rect 13426 8750 13846 8778
rect 13874 8750 13879 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 0 8736 400 8750
rect 20600 8736 21000 8750
rect 11881 8694 11886 8722
rect 11914 8694 13118 8722
rect 13146 8694 13151 8722
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 8297 8526 8302 8554
rect 8330 8526 8694 8554
rect 8722 8526 8727 8554
rect 10649 8526 10654 8554
rect 10682 8526 11382 8554
rect 11410 8526 12726 8554
rect 12754 8526 12838 8554
rect 12866 8526 12871 8554
rect 8913 8414 8918 8442
rect 8946 8414 8951 8442
rect 8918 8386 8946 8414
rect 8918 8358 9982 8386
rect 10010 8358 10015 8386
rect 10537 8358 10542 8386
rect 10570 8358 11214 8386
rect 11242 8358 12502 8386
rect 12530 8358 12535 8386
rect 7121 8302 7126 8330
rect 7154 8302 9702 8330
rect 9730 8302 10598 8330
rect 10626 8302 10631 8330
rect 8409 8246 8414 8274
rect 8442 8246 8974 8274
rect 9002 8246 9007 8274
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 9249 8078 9254 8106
rect 9282 8078 9366 8106
rect 9394 8078 9399 8106
rect 15946 8022 18830 8050
rect 18858 8022 18863 8050
rect 15946 7938 15974 8022
rect 12721 7910 12726 7938
rect 12754 7910 13510 7938
rect 13538 7910 13543 7938
rect 13617 7910 13622 7938
rect 13650 7910 14182 7938
rect 14210 7910 15974 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 20600 7770 21000 7784
rect 10201 7742 10206 7770
rect 10234 7742 11774 7770
rect 11802 7742 12614 7770
rect 12642 7742 13006 7770
rect 13034 7742 13039 7770
rect 13113 7742 13118 7770
rect 13146 7742 13454 7770
rect 20001 7742 20006 7770
rect 20034 7742 21000 7770
rect 8857 7686 8862 7714
rect 8890 7686 9198 7714
rect 9226 7686 9231 7714
rect 9305 7686 9310 7714
rect 9338 7686 9926 7714
rect 9954 7686 9959 7714
rect 12273 7686 12278 7714
rect 12306 7686 13062 7714
rect 13090 7686 13095 7714
rect 13426 7658 13454 7742
rect 20600 7728 21000 7742
rect 7681 7630 7686 7658
rect 7714 7630 8918 7658
rect 8946 7630 8951 7658
rect 9030 7630 9142 7658
rect 9170 7630 9175 7658
rect 12665 7630 12670 7658
rect 12698 7630 13118 7658
rect 13146 7630 13151 7658
rect 13426 7630 13790 7658
rect 13818 7630 18830 7658
rect 18858 7630 18863 7658
rect 9030 7490 9058 7630
rect 9809 7574 9814 7602
rect 9842 7574 10150 7602
rect 10178 7574 10183 7602
rect 11041 7518 11046 7546
rect 11074 7518 11438 7546
rect 11466 7518 11471 7546
rect 12329 7518 12334 7546
rect 12362 7518 12726 7546
rect 12754 7518 12759 7546
rect 9025 7462 9030 7490
rect 9058 7462 9063 7490
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 20600 7434 21000 7448
rect 20001 7406 20006 7434
rect 20034 7406 21000 7434
rect 20600 7392 21000 7406
rect 11433 7294 11438 7322
rect 11466 7294 12110 7322
rect 12138 7294 12143 7322
rect 10705 7238 10710 7266
rect 10738 7238 12334 7266
rect 12362 7238 12782 7266
rect 12810 7238 12815 7266
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 8745 2030 8750 2058
rect 8778 2030 9366 2058
rect 9394 2030 9399 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 10089 1694 10094 1722
rect 10122 1694 10878 1722
rect 10906 1694 10911 1722
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 11382 11718 11410 11746
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 11382 11158 11410 11186
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 9904 10990 10064 11746
rect 11382 11746 11410 11751
rect 11382 11186 11410 11718
rect 11382 11153 11410 11158
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _095_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11536 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _096_
timestamp 1698175906
transform 1 0 11144 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _097_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11256 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _098_
timestamp 1698175906
transform -1 0 10472 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _099_
timestamp 1698175906
transform -1 0 9576 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _100_
timestamp 1698175906
transform 1 0 9744 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _101_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9856 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10640 0 1 8624
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9632 0 1 8624
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11424 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1698175906
transform -1 0 9800 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10976 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _107_
timestamp 1698175906
transform -1 0 11424 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11592 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_
timestamp 1698175906
transform 1 0 11648 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _110_
timestamp 1698175906
transform -1 0 9688 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _111_
timestamp 1698175906
transform 1 0 8680 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8680 0 -1 10192
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _113_
timestamp 1698175906
transform -1 0 8960 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _114_
timestamp 1698175906
transform -1 0 10136 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform -1 0 7280 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 6944 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _117_
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698175906
transform -1 0 9744 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform 1 0 11704 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _120_
timestamp 1698175906
transform -1 0 10136 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _121_
timestamp 1698175906
transform 1 0 9744 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11200 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _123_
timestamp 1698175906
transform -1 0 12432 0 1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _124_
timestamp 1698175906
transform -1 0 11984 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform 1 0 11088 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11368 0 1 12544
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _127_
timestamp 1698175906
transform 1 0 11200 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _128_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9296 0 -1 11760
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _129_
timestamp 1698175906
transform 1 0 13104 0 1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _130_
timestamp 1698175906
transform 1 0 13384 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform -1 0 9912 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform 1 0 10360 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7952 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _134_
timestamp 1698175906
transform 1 0 8176 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _135_
timestamp 1698175906
transform 1 0 10472 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _136_
timestamp 1698175906
transform 1 0 11536 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _137_
timestamp 1698175906
transform -1 0 9296 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _138_
timestamp 1698175906
transform 1 0 9912 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _139_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _140_
timestamp 1698175906
transform -1 0 11032 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _141_
timestamp 1698175906
transform -1 0 9632 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _142_
timestamp 1698175906
transform -1 0 8960 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _143_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7112 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _144_
timestamp 1698175906
transform -1 0 7336 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _145_
timestamp 1698175906
transform 1 0 12936 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _146_
timestamp 1698175906
transform 1 0 12768 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _147_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12936 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _148_
timestamp 1698175906
transform 1 0 12208 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _149_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9296 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _150_
timestamp 1698175906
transform 1 0 6720 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _151_
timestamp 1698175906
transform 1 0 6272 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _152_
timestamp 1698175906
transform -1 0 10696 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _153_
timestamp 1698175906
transform -1 0 8064 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _154_
timestamp 1698175906
transform 1 0 7392 0 -1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _155_
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _156_
timestamp 1698175906
transform -1 0 9352 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _157_
timestamp 1698175906
transform -1 0 7728 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698175906
transform -1 0 6944 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _159_
timestamp 1698175906
transform 1 0 6720 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform 1 0 8512 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _161_
timestamp 1698175906
transform -1 0 9352 0 -1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _162_
timestamp 1698175906
transform -1 0 9072 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _163_
timestamp 1698175906
transform 1 0 8736 0 -1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _164_
timestamp 1698175906
transform -1 0 8512 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _165_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11984 0 1 11760
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _166_
timestamp 1698175906
transform 1 0 11256 0 -1 11760
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _167_
timestamp 1698175906
transform -1 0 7672 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _168_
timestamp 1698175906
transform -1 0 7224 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _169_
timestamp 1698175906
transform 1 0 7168 0 1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _170_
timestamp 1698175906
transform 1 0 6776 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _171_
timestamp 1698175906
transform -1 0 10304 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _172_
timestamp 1698175906
transform -1 0 9912 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _173_
timestamp 1698175906
transform -1 0 10360 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _174_
timestamp 1698175906
transform 1 0 14168 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _175_
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _176_
timestamp 1698175906
transform 1 0 12656 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform 1 0 13776 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _178_
timestamp 1698175906
transform -1 0 13440 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _179_
timestamp 1698175906
transform 1 0 13496 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _180_
timestamp 1698175906
transform 1 0 11144 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _181_
timestamp 1698175906
transform -1 0 14280 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _182_
timestamp 1698175906
transform 1 0 13440 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _183_
timestamp 1698175906
transform 1 0 12992 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _184_
timestamp 1698175906
transform 1 0 12040 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _185_
timestamp 1698175906
transform -1 0 12432 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _186_
timestamp 1698175906
transform -1 0 13776 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _187_
timestamp 1698175906
transform -1 0 12936 0 1 7840
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _188_
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _189_
timestamp 1698175906
transform -1 0 10808 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _190_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9296 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _191_
timestamp 1698175906
transform -1 0 6944 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _192_
timestamp 1698175906
transform 1 0 11200 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _193_
timestamp 1698175906
transform 1 0 13048 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_
timestamp 1698175906
transform 1 0 7952 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1698175906
transform 1 0 7896 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _196_
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _197_
timestamp 1698175906
transform -1 0 11648 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _198_
timestamp 1698175906
transform -1 0 7448 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _199_
timestamp 1698175906
transform 1 0 12264 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _200_
timestamp 1698175906
transform -1 0 7112 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1698175906
transform -1 0 7504 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_
timestamp 1698175906
transform -1 0 6720 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform 1 0 7224 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform 1 0 7504 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform 1 0 10808 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform -1 0 7392 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform -1 0 7560 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform 1 0 8848 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform 1 0 13328 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 13272 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 13272 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 12656 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 9632 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _217_
timestamp 1698175906
transform -1 0 13160 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _218_
timestamp 1698175906
transform -1 0 7728 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _219_
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9296 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__CLK
timestamp 1698175906
transform 1 0 7672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__CLK
timestamp 1698175906
transform 1 0 13272 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__CLK
timestamp 1698175906
transform 1 0 14784 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__CLK
timestamp 1698175906
transform 1 0 10248 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1698175906
transform 1 0 9632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__CLK
timestamp 1698175906
transform -1 0 12320 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__CLK
timestamp 1698175906
transform 1 0 12096 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__CLK
timestamp 1698175906
transform 1 0 7560 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__CLK
timestamp 1698175906
transform 1 0 14000 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__CLK
timestamp 1698175906
transform 1 0 7224 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__CLK
timestamp 1698175906
transform 1 0 7616 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK
timestamp 1698175906
transform 1 0 7112 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1698175906
transform 1 0 8960 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform 1 0 9240 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 7840 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 7672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 8736 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 15064 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 15008 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 15008 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 14560 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 14392 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 9520 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 9632 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9632 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 11592 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_198
timestamp 1698175906
transform 1 0 11760 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_202
timestamp 1698175906
transform 1 0 11984 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_144
timestamp 1698175906
transform 1 0 8736 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_171
timestamp 1698175906
transform 1 0 10248 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_203
timestamp 1698175906
transform 1 0 12040 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 12264 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 16128 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 10248 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_175 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10472 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_191 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11368 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_199
timestamp 1698175906
transform 1 0 11816 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_203
timestamp 1698175906
transform 1 0 12040 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_205
timestamp 1698175906
transform 1 0 12152 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698175906
transform 1 0 12320 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_115
timestamp 1698175906
transform 1 0 7112 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_146
timestamp 1698175906
transform 1 0 8848 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_150
timestamp 1698175906
transform 1 0 9072 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_158
timestamp 1698175906
transform 1 0 9520 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_165
timestamp 1698175906
transform 1 0 9912 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698175906
transform 1 0 10360 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_206
timestamp 1698175906
transform 1 0 12208 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_236
timestamp 1698175906
transform 1 0 13888 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_240
timestamp 1698175906
transform 1 0 14112 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 14336 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 8288 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_155
timestamp 1698175906
transform 1 0 9352 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_163
timestamp 1698175906
transform 1 0 9800 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_172
timestamp 1698175906
transform 1 0 10304 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_180
timestamp 1698175906
transform 1 0 10752 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_200
timestamp 1698175906
transform 1 0 11872 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_204
timestamp 1698175906
transform 1 0 12096 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_243
timestamp 1698175906
transform 1 0 14280 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_247
timestamp 1698175906
transform 1 0 14504 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 16296 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_314
timestamp 1698175906
transform 1 0 18256 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_322
timestamp 1698175906
transform 1 0 18704 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_115
timestamp 1698175906
transform 1 0 7112 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_119
timestamp 1698175906
transform 1 0 7336 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_121
timestamp 1698175906
transform 1 0 7448 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_151
timestamp 1698175906
transform 1 0 9128 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_155
timestamp 1698175906
transform 1 0 9352 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698175906
transform 1 0 10248 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_185
timestamp 1698175906
transform 1 0 11032 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_192
timestamp 1698175906
transform 1 0 11424 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_208
timestamp 1698175906
transform 1 0 12320 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_234
timestamp 1698175906
transform 1 0 13776 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698175906
transform 1 0 14224 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 14336 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 18648 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_88
timestamp 1698175906
transform 1 0 5600 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_121
timestamp 1698175906
transform 1 0 7448 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_125
timestamp 1698175906
transform 1 0 7672 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_133
timestamp 1698175906
transform 1 0 8120 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_153
timestamp 1698175906
transform 1 0 9240 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_161
timestamp 1698175906
transform 1 0 9688 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_171
timestamp 1698175906
transform 1 0 10248 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_181
timestamp 1698175906
transform 1 0 10808 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_185
timestamp 1698175906
transform 1 0 11032 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_193
timestamp 1698175906
transform 1 0 11480 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 12376 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_224
timestamp 1698175906
transform 1 0 13216 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_254
timestamp 1698175906
transform 1 0 14896 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_258
timestamp 1698175906
transform 1 0 15120 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_274
timestamp 1698175906
transform 1 0 16016 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698175906
transform 1 0 16240 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 20048 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 20160 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_112
timestamp 1698175906
transform 1 0 6944 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_119
timestamp 1698175906
transform 1 0 7336 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_135
timestamp 1698175906
transform 1 0 8232 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_139
timestamp 1698175906
transform 1 0 8456 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_145
timestamp 1698175906
transform 1 0 8792 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_153
timestamp 1698175906
transform 1 0 9240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_157
timestamp 1698175906
transform 1 0 9464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_159
timestamp 1698175906
transform 1 0 9576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_177
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_191
timestamp 1698175906
transform 1 0 11368 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_207
timestamp 1698175906
transform 1 0 12264 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_211
timestamp 1698175906
transform 1 0 12488 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_213
timestamp 1698175906
transform 1 0 12600 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_228
timestamp 1698175906
transform 1 0 13440 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_232
timestamp 1698175906
transform 1 0 13664 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_239
timestamp 1698175906
transform 1 0 14056 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698175906
transform 1 0 14280 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 2240 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 4032 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 4480 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_80
timestamp 1698175906
transform 1 0 5152 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_82
timestamp 1698175906
transform 1 0 5264 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_112
timestamp 1698175906
transform 1 0 6944 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_114
timestamp 1698175906
transform 1 0 7056 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_123
timestamp 1698175906
transform 1 0 7560 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_127
timestamp 1698175906
transform 1 0 7784 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_135
timestamp 1698175906
transform 1 0 8232 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 8456 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_148
timestamp 1698175906
transform 1 0 8960 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_152
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_156
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_160
timestamp 1698175906
transform 1 0 9632 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_164
timestamp 1698175906
transform 1 0 9856 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_166
timestamp 1698175906
transform 1 0 9968 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_202
timestamp 1698175906
transform 1 0 11984 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698175906
transform 1 0 12208 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_228
timestamp 1698175906
transform 1 0 13440 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_234
timestamp 1698175906
transform 1 0 13776 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_266
timestamp 1698175906
transform 1 0 15568 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_274
timestamp 1698175906
transform 1 0 16016 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 16240 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 20048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 20160 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_118
timestamp 1698175906
transform 1 0 7280 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_122
timestamp 1698175906
transform 1 0 7504 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_124
timestamp 1698175906
transform 1 0 7616 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_154
timestamp 1698175906
transform 1 0 9296 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_156
timestamp 1698175906
transform 1 0 9408 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_185
timestamp 1698175906
transform 1 0 11032 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_198
timestamp 1698175906
transform 1 0 11760 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_210
timestamp 1698175906
transform 1 0 12432 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_218
timestamp 1698175906
transform 1 0 12880 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_228
timestamp 1698175906
transform 1 0 13440 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 14336 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 2240 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 4032 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 4480 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_88
timestamp 1698175906
transform 1 0 5600 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_90
timestamp 1698175906
transform 1 0 5712 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_126
timestamp 1698175906
transform 1 0 7728 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_130
timestamp 1698175906
transform 1 0 7952 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_138
timestamp 1698175906
transform 1 0 8400 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_142
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_152
timestamp 1698175906
transform 1 0 9184 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_246
timestamp 1698175906
transform 1 0 14448 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_250
timestamp 1698175906
transform 1 0 14672 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_266
timestamp 1698175906
transform 1 0 15568 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_274
timestamp 1698175906
transform 1 0 16016 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 16240 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 18256 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 18704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_255
timestamp 1698175906
transform 1 0 14952 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_287
timestamp 1698175906
transform 1 0 16744 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_303
timestamp 1698175906
transform 1 0 17640 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 2240 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 4032 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 4480 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_88
timestamp 1698175906
transform 1 0 5600 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_92
timestamp 1698175906
transform 1 0 5824 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_122
timestamp 1698175906
transform 1 0 7504 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_126
timestamp 1698175906
transform 1 0 7728 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_134
timestamp 1698175906
transform 1 0 8176 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_138
timestamp 1698175906
transform 1 0 8400 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_148
timestamp 1698175906
transform 1 0 8960 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_155
timestamp 1698175906
transform 1 0 9352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_161
timestamp 1698175906
transform 1 0 9688 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_179
timestamp 1698175906
transform 1 0 10696 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_194
timestamp 1698175906
transform 1 0 11536 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_202
timestamp 1698175906
transform 1 0 11984 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_216
timestamp 1698175906
transform 1 0 12768 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_218
timestamp 1698175906
transform 1 0 12880 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_225
timestamp 1698175906
transform 1 0 13272 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_255
timestamp 1698175906
transform 1 0 14952 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_259
timestamp 1698175906
transform 1 0 15176 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_275
timestamp 1698175906
transform 1 0 16072 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 16296 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 20048 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 20160 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 2240 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 2464 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_115
timestamp 1698175906
transform 1 0 7112 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_117
timestamp 1698175906
transform 1 0 7224 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_126
timestamp 1698175906
transform 1 0 7728 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_132
timestamp 1698175906
transform 1 0 8064 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_140
timestamp 1698175906
transform 1 0 8512 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_142
timestamp 1698175906
transform 1 0 8624 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698175906
transform 1 0 10304 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 10416 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_177
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_185
timestamp 1698175906
transform 1 0 11032 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_209
timestamp 1698175906
transform 1 0 12376 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_225
timestamp 1698175906
transform 1 0 13272 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_227
timestamp 1698175906
transform 1 0 13384 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_236
timestamp 1698175906
transform 1 0 13888 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698175906
transform 1 0 14280 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 2240 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 4032 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 4480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_76
timestamp 1698175906
transform 1 0 4928 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_78
timestamp 1698175906
transform 1 0 5040 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_113
timestamp 1698175906
transform 1 0 7000 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_117
timestamp 1698175906
transform 1 0 7224 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_119
timestamp 1698175906
transform 1 0 7336 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_129
timestamp 1698175906
transform 1 0 7896 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698175906
transform 1 0 8344 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 8456 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_150
timestamp 1698175906
transform 1 0 9072 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_164
timestamp 1698175906
transform 1 0 9856 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_180
timestamp 1698175906
transform 1 0 10752 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_188
timestamp 1698175906
transform 1 0 11200 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_199
timestamp 1698175906
transform 1 0 11816 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698175906
transform 1 0 12264 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_220
timestamp 1698175906
transform 1 0 12992 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_224
timestamp 1698175906
transform 1 0 13216 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_254
timestamp 1698175906
transform 1 0 14896 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_258
timestamp 1698175906
transform 1 0 15120 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_274
timestamp 1698175906
transform 1 0 16016 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698175906
transform 1 0 16240 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 2240 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 2464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_112
timestamp 1698175906
transform 1 0 6944 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_128
timestamp 1698175906
transform 1 0 7840 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_169
timestamp 1698175906
transform 1 0 10136 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_173
timestamp 1698175906
transform 1 0 10360 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_185
timestamp 1698175906
transform 1 0 11032 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_189
timestamp 1698175906
transform 1 0 11256 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_202
timestamp 1698175906
transform 1 0 11984 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_218
timestamp 1698175906
transform 1 0 12880 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_231
timestamp 1698175906
transform 1 0 13608 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_239
timestamp 1698175906
transform 1 0 14056 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 14280 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698175906
transform 1 0 5152 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_84
timestamp 1698175906
transform 1 0 5376 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_115
timestamp 1698175906
transform 1 0 7112 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_119
timestamp 1698175906
transform 1 0 7336 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_135
timestamp 1698175906
transform 1 0 8232 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 8456 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_150
timestamp 1698175906
transform 1 0 9072 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_152
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_159
timestamp 1698175906
transform 1 0 9576 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_161
timestamp 1698175906
transform 1 0 9688 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_168
timestamp 1698175906
transform 1 0 10080 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_172
timestamp 1698175906
transform 1 0 10304 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_179
timestamp 1698175906
transform 1 0 10696 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_216
timestamp 1698175906
transform 1 0 12768 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_220
timestamp 1698175906
transform 1 0 12992 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_250
timestamp 1698175906
transform 1 0 14672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_254
timestamp 1698175906
transform 1 0 14896 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_270
timestamp 1698175906
transform 1 0 15792 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698175906
transform 1 0 16240 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_69
timestamp 1698175906
transform 1 0 4536 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_85
timestamp 1698175906
transform 1 0 5432 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_93
timestamp 1698175906
transform 1 0 5880 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_97
timestamp 1698175906
transform 1 0 6104 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_99
timestamp 1698175906
transform 1 0 6216 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698175906
transform 1 0 6496 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_125
timestamp 1698175906
transform 1 0 7672 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_129
timestamp 1698175906
transform 1 0 7896 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_138
timestamp 1698175906
transform 1 0 8400 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_154
timestamp 1698175906
transform 1 0 9296 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_168
timestamp 1698175906
transform 1 0 10080 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698175906
transform 1 0 10304 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 10416 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_186
timestamp 1698175906
transform 1 0 11088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_190
timestamp 1698175906
transform 1 0 11312 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_210
timestamp 1698175906
transform 1 0 12432 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_226
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_231
timestamp 1698175906
transform 1 0 13608 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_239
timestamp 1698175906
transform 1 0 14056 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698175906
transform 1 0 14280 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 18648 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 2240 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 4032 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 4480 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_88
timestamp 1698175906
transform 1 0 5600 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_92
timestamp 1698175906
transform 1 0 5824 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_123
timestamp 1698175906
transform 1 0 7560 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_127
timestamp 1698175906
transform 1 0 7784 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_131
timestamp 1698175906
transform 1 0 8008 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_133
timestamp 1698175906
transform 1 0 8120 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_189
timestamp 1698175906
transform 1 0 11256 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_205
timestamp 1698175906
transform 1 0 12152 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 12376 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_218
timestamp 1698175906
transform 1 0 12880 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_250
timestamp 1698175906
transform 1 0 14672 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_266
timestamp 1698175906
transform 1 0 15568 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_274
timestamp 1698175906
transform 1 0 16016 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698175906
transform 1 0 16240 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 20048 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 20160 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 2240 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 2464 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_113
timestamp 1698175906
transform 1 0 7000 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_158
timestamp 1698175906
transform 1 0 9520 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_162
timestamp 1698175906
transform 1 0 9744 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_170
timestamp 1698175906
transform 1 0 10192 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698175906
transform 1 0 10416 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_181
timestamp 1698175906
transform 1 0 10808 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_185
timestamp 1698175906
transform 1 0 11032 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_187
timestamp 1698175906
transform 1 0 11144 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_223
timestamp 1698175906
transform 1 0 13160 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_227
timestamp 1698175906
transform 1 0 13384 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698175906
transform 1 0 14280 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698175906
transform 1 0 12208 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_193
timestamp 1698175906
transform 1 0 11480 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_197
timestamp 1698175906
transform 1 0 11704 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_225
timestamp 1698175906
transform 1 0 13272 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_333
timestamp 1698175906
transform 1 0 19320 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_341
timestamp 1698175906
transform 1 0 19768 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_174
timestamp 1698175906
transform 1 0 10416 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_190
timestamp 1698175906
transform 1 0 11312 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_198
timestamp 1698175906
transform 1 0 11760 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_202
timestamp 1698175906
transform 1 0 11984 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_204
timestamp 1698175906
transform 1 0 12096 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 14000 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 15792 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 16240 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_266
timestamp 1698175906
transform 1 0 15568 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_270
timestamp 1698175906
transform 1 0 15792 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita31_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19992 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita31_26
timestamp 1698175906
transform -1 0 12376 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 18760 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 18760 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 18760 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 2240 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 13272 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 2240 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 8792 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 8736 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform -1 0 2240 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 2240 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 2240 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 2240 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 18760 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 2240 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 2240 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 18760 0 -1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 10640 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13440 400 13496 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 12432 20600 12488 21000 0 FreeSans 224 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 20600 9744 21000 9800 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 20600 7728 21000 7784 0 FreeSans 224 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 0 10416 400 10472 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 20600 17808 21000 17864 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 11760 20600 11816 21000 0 FreeSans 224 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 0 10752 400 10808 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 12096 20600 12152 21000 0 FreeSans 224 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 20600 10752 21000 10808 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 8736 0 8792 400 0 FreeSans 224 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 11424 20600 11480 21000 0 FreeSans 224 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 11760 400 11816 0 FreeSans 224 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 13104 400 13160 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 10080 0 10136 400 0 FreeSans 224 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 0 11424 400 11480 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 0 12768 400 12824 0 FreeSans 224 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 0 8736 400 8792 0 FreeSans 224 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 20600 12432 21000 12488 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 12768 20600 12824 21000 0 FreeSans 224 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 0 9744 400 9800 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 9072 400 9128 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 20600 7392 21000 7448 0 FreeSans 224 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal3 12908 7644 12908 7644 0 _000_
rlabel metal2 10668 13300 10668 13300 0 _001_
rlabel metal2 8820 9436 8820 9436 0 _002_
rlabel metal2 6468 9352 6468 9352 0 _003_
rlabel metal2 11648 13468 11648 13468 0 _004_
rlabel metal2 13524 12516 13524 12516 0 _005_
rlabel metal2 9436 10920 9436 10920 0 _006_
rlabel metal2 8372 13454 8372 13454 0 _007_
rlabel metal2 10948 7770 10948 7770 0 _008_
rlabel metal3 11032 9212 11032 9212 0 _009_
rlabel metal2 6972 8680 6972 8680 0 _010_
rlabel metal3 12544 7532 12544 7532 0 _011_
rlabel metal2 6636 12516 6636 12516 0 _012_
rlabel metal2 7112 10780 7112 10780 0 _013_
rlabel metal2 6244 11480 6244 11480 0 _014_
rlabel metal3 8316 7644 8316 7644 0 _015_
rlabel metal2 7980 8204 7980 8204 0 _016_
rlabel metal3 11284 11592 11284 11592 0 _017_
rlabel metal2 6888 10052 6888 10052 0 _018_
rlabel metal2 7084 13300 7084 13300 0 _019_
rlabel metal2 9324 7112 9324 7112 0 _020_
rlabel metal2 14644 10584 14644 10584 0 _021_
rlabel metal2 13748 8848 13748 8848 0 _022_
rlabel metal2 13580 11368 13580 11368 0 _023_
rlabel metal2 12292 9800 12292 9800 0 _024_
rlabel metal2 13636 10724 13636 10724 0 _025_
rlabel metal2 13244 8148 13244 8148 0 _026_
rlabel metal3 12684 7700 12684 7700 0 _027_
rlabel metal2 7000 11956 7000 11956 0 _028_
rlabel metal3 6608 12684 6608 12684 0 _029_
rlabel metal2 7476 12656 7476 12656 0 _030_
rlabel metal2 7812 11396 7812 11396 0 _031_
rlabel metal2 7532 11312 7532 11312 0 _032_
rlabel metal3 9744 10780 9744 10780 0 _033_
rlabel metal2 7028 10556 7028 10556 0 _034_
rlabel metal2 6776 11620 6776 11620 0 _035_
rlabel metal2 8792 7700 8792 7700 0 _036_
rlabel metal2 9044 7672 9044 7672 0 _037_
rlabel metal2 8428 8288 8428 8288 0 _038_
rlabel metal2 11536 11788 11536 11788 0 _039_
rlabel metal2 7476 10332 7476 10332 0 _040_
rlabel metal2 7392 12740 7392 12740 0 _041_
rlabel metal3 9996 7588 9996 7588 0 _042_
rlabel metal2 14588 10472 14588 10472 0 _043_
rlabel metal2 14812 10178 14812 10178 0 _044_
rlabel metal2 13860 8400 13860 8400 0 _045_
rlabel metal2 13916 9128 13916 9128 0 _046_
rlabel metal2 13300 9072 13300 9072 0 _047_
rlabel metal3 12572 11060 12572 11060 0 _048_
rlabel metal2 13944 11172 13944 11172 0 _049_
rlabel metal2 12236 9576 12236 9576 0 _050_
rlabel metal2 12348 10416 12348 10416 0 _051_
rlabel metal3 13132 7924 13132 7924 0 _052_
rlabel metal2 10780 13468 10780 13468 0 _053_
rlabel metal2 10948 9016 10948 9016 0 _054_
rlabel metal2 10668 8680 10668 8680 0 _055_
rlabel metal3 10752 9492 10752 9492 0 _056_
rlabel metal2 11900 8904 11900 8904 0 _057_
rlabel metal2 9464 11564 9464 11564 0 _058_
rlabel metal2 9828 12516 9828 12516 0 _059_
rlabel metal2 10948 9632 10948 9632 0 _060_
rlabel metal2 6972 9240 6972 9240 0 _061_
rlabel metal2 8708 9100 8708 9100 0 _062_
rlabel metal2 10948 10080 10948 10080 0 _063_
rlabel metal3 9324 9548 9324 9548 0 _064_
rlabel metal2 11340 7840 11340 7840 0 _065_
rlabel metal2 11396 9828 11396 9828 0 _066_
rlabel metal2 11788 10920 11788 10920 0 _067_
rlabel metal2 11900 10640 11900 10640 0 _068_
rlabel metal2 7420 10528 7420 10528 0 _069_
rlabel metal2 8820 10528 8820 10528 0 _070_
rlabel metal2 8904 9268 8904 9268 0 _071_
rlabel metal2 7196 9660 7196 9660 0 _072_
rlabel metal2 6916 11900 6916 11900 0 _073_
rlabel metal2 6776 8932 6776 8932 0 _074_
rlabel metal3 10556 12628 10556 12628 0 _075_
rlabel metal2 11452 12208 11452 12208 0 _076_
rlabel metal2 9968 12068 9968 12068 0 _077_
rlabel metal2 11564 12208 11564 12208 0 _078_
rlabel metal2 11788 11564 11788 11564 0 _079_
rlabel metal3 11900 12796 11900 12796 0 _080_
rlabel metal3 10892 9604 10892 9604 0 _081_
rlabel metal2 12068 9492 12068 9492 0 _082_
rlabel metal2 13468 11368 13468 11368 0 _083_
rlabel metal2 9716 11312 9716 11312 0 _084_
rlabel metal2 13356 12348 13356 12348 0 _085_
rlabel metal3 7924 12740 7924 12740 0 _086_
rlabel metal2 8316 12992 8316 12992 0 _087_
rlabel metal2 7140 8512 7140 8512 0 _088_
rlabel metal2 10220 8092 10220 8092 0 _089_
rlabel metal2 8932 8876 8932 8876 0 _090_
rlabel metal2 10052 10808 10052 10808 0 _091_
rlabel metal3 9212 10892 9212 10892 0 _092_
rlabel metal2 7532 9674 7532 9674 0 _093_
rlabel metal2 7252 9044 7252 9044 0 _094_
rlabel metal3 1239 13468 1239 13468 0 clk
rlabel metal2 11676 10220 11676 10220 0 clknet_0_clk
rlabel metal2 7476 13188 7476 13188 0 clknet_1_0__leaf_clk
rlabel metal2 11144 13524 11144 13524 0 clknet_1_1__leaf_clk
rlabel metal3 9772 12012 9772 12012 0 dut31.count\[0\]
rlabel metal2 9464 13580 9464 13580 0 dut31.count\[1\]
rlabel metal3 11788 7308 11788 7308 0 dut31.count\[2\]
rlabel metal2 10108 9520 10108 9520 0 dut31.count\[3\]
rlabel metal2 12880 18620 12880 18620 0 net1
rlabel metal3 9044 7700 9044 7700 0 net10
rlabel metal2 12320 12292 12320 12292 0 net11
rlabel metal2 9044 1764 9044 1764 0 net12
rlabel metal3 3178 11956 3178 11956 0 net13
rlabel metal2 2044 13300 2044 13300 0 net14
rlabel metal2 10388 4284 10388 4284 0 net15
rlabel metal2 5964 11144 5964 11144 0 net16
rlabel metal2 5572 12712 5572 12712 0 net17
rlabel metal2 5908 8792 5908 8792 0 net18
rlabel metal2 18844 12516 18844 12516 0 net19
rlabel metal2 14812 8400 14812 8400 0 net2
rlabel metal2 14308 16128 14308 16128 0 net20
rlabel metal2 2156 10024 2156 10024 0 net21
rlabel metal3 3178 9212 3178 9212 0 net22
rlabel metal2 13804 7476 13804 7476 0 net23
rlabel metal3 11032 13076 11032 13076 0 net24
rlabel metal2 20132 17976 20132 17976 0 net25
rlabel metal2 12180 18732 12180 18732 0 net26
rlabel metal2 14140 11312 14140 11312 0 net3
rlabel metal3 15022 9940 15022 9940 0 net4
rlabel metal2 14196 7756 14196 7756 0 net5
rlabel metal2 7532 10472 7532 10472 0 net6
rlabel metal2 12992 13524 12992 13524 0 net7
rlabel metal3 4004 11172 4004 11172 0 net8
rlabel metal2 14308 10388 14308 10388 0 net9
rlabel metal2 12460 19677 12460 19677 0 segm[0]
rlabel metal2 20020 8820 20020 8820 0 segm[10]
rlabel metal3 20321 11452 20321 11452 0 segm[11]
rlabel metal2 20020 9828 20020 9828 0 segm[12]
rlabel metal2 20020 7924 20020 7924 0 segm[13]
rlabel metal3 679 10444 679 10444 0 segm[1]
rlabel metal2 12012 18872 12012 18872 0 segm[3]
rlabel metal3 679 10780 679 10780 0 segm[4]
rlabel metal2 20020 11004 20020 11004 0 segm[6]
rlabel metal3 9072 2044 9072 2044 0 segm[7]
rlabel metal2 11452 19845 11452 19845 0 segm[8]
rlabel metal2 9100 1029 9100 1029 0 segm[9]
rlabel metal3 679 11788 679 11788 0 sel[0]
rlabel metal3 679 13132 679 13132 0 sel[10]
rlabel metal3 10500 1708 10500 1708 0 sel[11]
rlabel metal3 679 11452 679 11452 0 sel[1]
rlabel metal3 679 12796 679 12796 0 sel[2]
rlabel metal3 679 8764 679 8764 0 sel[3]
rlabel metal2 20020 12628 20020 12628 0 sel[4]
rlabel metal2 12796 19873 12796 19873 0 sel[5]
rlabel metal3 679 9772 679 9772 0 sel[6]
rlabel metal3 679 9100 679 9100 0 sel[7]
rlabel metal2 20020 7504 20020 7504 0 sel[8]
rlabel metal2 11116 19873 11116 19873 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
