magic
tech gf180mcuD
magscale 1 5
timestamp 1699643023
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 9417 19055 9423 19081
rect 9449 19055 9455 19081
rect 11097 19055 11103 19081
rect 11129 19055 11135 19081
rect 9865 18999 9871 19025
rect 9897 18999 9903 19025
rect 11993 18999 11999 19025
rect 12025 18999 12031 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 10375 18745 10401 18751
rect 10375 18713 10401 18719
rect 9865 18607 9871 18633
rect 9897 18607 9903 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 9591 18353 9617 18359
rect 9591 18321 9617 18327
rect 9193 18215 9199 18241
rect 9225 18215 9231 18241
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 9921 13903 9927 13929
rect 9953 13903 9959 13929
rect 18937 13903 18943 13929
rect 18969 13903 18975 13929
rect 11607 13873 11633 13879
rect 10257 13847 10263 13873
rect 10289 13847 10295 13873
rect 11321 13847 11327 13873
rect 11353 13847 11359 13873
rect 19945 13847 19951 13873
rect 19977 13847 19983 13873
rect 11607 13841 11633 13847
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 10711 13593 10737 13599
rect 9865 13567 9871 13593
rect 9897 13567 9903 13593
rect 10711 13561 10737 13567
rect 20007 13593 20033 13599
rect 20007 13561 20033 13567
rect 11047 13537 11073 13543
rect 8465 13511 8471 13537
rect 8497 13511 8503 13537
rect 10929 13511 10935 13537
rect 10961 13511 10967 13537
rect 18825 13511 18831 13537
rect 18857 13511 18863 13537
rect 11047 13505 11073 13511
rect 10767 13481 10793 13487
rect 8801 13455 8807 13481
rect 8833 13455 8839 13481
rect 10767 13449 10793 13455
rect 11159 13481 11185 13487
rect 11159 13449 11185 13455
rect 11215 13481 11241 13487
rect 11215 13449 11241 13455
rect 13175 13481 13201 13487
rect 13175 13449 13201 13455
rect 13231 13481 13257 13487
rect 13231 13449 13257 13455
rect 10095 13425 10121 13431
rect 10095 13393 10121 13399
rect 10655 13425 10681 13431
rect 10655 13393 10681 13399
rect 12559 13425 12585 13431
rect 12559 13393 12585 13399
rect 13343 13425 13369 13431
rect 13343 13393 13369 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 7519 13257 7545 13263
rect 7519 13225 7545 13231
rect 9087 13257 9113 13263
rect 9087 13225 9113 13231
rect 9759 13257 9785 13263
rect 9759 13225 9785 13231
rect 9143 13201 9169 13207
rect 9143 13169 9169 13175
rect 9815 13201 9841 13207
rect 14513 13175 14519 13201
rect 14545 13175 14551 13201
rect 9815 13169 9841 13175
rect 8639 13145 8665 13151
rect 7289 13119 7295 13145
rect 7321 13119 7327 13145
rect 8639 13113 8665 13119
rect 8863 13145 8889 13151
rect 8863 13113 8889 13119
rect 8975 13145 9001 13151
rect 9423 13145 9449 13151
rect 9249 13119 9255 13145
rect 9281 13119 9287 13145
rect 10481 13119 10487 13145
rect 10513 13119 10519 13145
rect 12721 13119 12727 13145
rect 12753 13119 12759 13145
rect 14401 13119 14407 13145
rect 14433 13119 14439 13145
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 8975 13113 9001 13119
rect 9423 13113 9449 13119
rect 8919 13089 8945 13095
rect 12111 13089 12137 13095
rect 5833 13063 5839 13089
rect 5865 13063 5871 13089
rect 6897 13063 6903 13089
rect 6929 13063 6935 13089
rect 10817 13063 10823 13089
rect 10849 13063 10855 13089
rect 11881 13063 11887 13089
rect 11913 13063 11919 13089
rect 8919 13057 8945 13063
rect 12111 13057 12137 13063
rect 12335 13089 12361 13095
rect 13113 13063 13119 13089
rect 13145 13063 13151 13089
rect 14177 13063 14183 13089
rect 14209 13063 14215 13089
rect 19945 13063 19951 13089
rect 19977 13063 19983 13089
rect 12335 13057 12361 13063
rect 9759 13033 9785 13039
rect 9759 13001 9785 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 967 12809 993 12815
rect 9871 12809 9897 12815
rect 20007 12809 20033 12815
rect 8241 12783 8247 12809
rect 8273 12783 8279 12809
rect 9305 12783 9311 12809
rect 9337 12783 9343 12809
rect 13729 12783 13735 12809
rect 13761 12783 13767 12809
rect 967 12777 993 12783
rect 9871 12777 9897 12783
rect 20007 12777 20033 12783
rect 7463 12753 7489 12759
rect 9479 12753 9505 12759
rect 2137 12727 2143 12753
rect 2169 12727 2175 12753
rect 7905 12727 7911 12753
rect 7937 12727 7943 12753
rect 7463 12721 7489 12727
rect 9479 12721 9505 12727
rect 11047 12753 11073 12759
rect 11047 12721 11073 12727
rect 11327 12753 11353 12759
rect 11327 12721 11353 12727
rect 11439 12753 11465 12759
rect 11439 12721 11465 12727
rect 11607 12753 11633 12759
rect 12273 12727 12279 12753
rect 12305 12727 12311 12753
rect 13953 12727 13959 12753
rect 13985 12727 13991 12753
rect 18825 12727 18831 12753
rect 18857 12727 18863 12753
rect 11607 12721 11633 12727
rect 9641 12671 9647 12697
rect 9673 12671 9679 12697
rect 11937 12671 11943 12697
rect 11969 12671 11975 12697
rect 12665 12671 12671 12697
rect 12697 12671 12703 12697
rect 7519 12641 7545 12647
rect 7519 12609 7545 12615
rect 7631 12641 7657 12647
rect 7631 12609 7657 12615
rect 10991 12641 11017 12647
rect 10991 12609 11017 12615
rect 11103 12641 11129 12647
rect 11103 12609 11129 12615
rect 11551 12641 11577 12647
rect 11551 12609 11577 12615
rect 12111 12641 12137 12647
rect 14065 12615 14071 12641
rect 14097 12615 14103 12641
rect 12111 12609 12137 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 7687 12473 7713 12479
rect 7687 12441 7713 12447
rect 8135 12473 8161 12479
rect 9199 12473 9225 12479
rect 8969 12447 8975 12473
rect 9001 12447 9007 12473
rect 8135 12441 8161 12447
rect 9199 12441 9225 12447
rect 12671 12473 12697 12479
rect 12671 12441 12697 12447
rect 13063 12473 13089 12479
rect 13063 12441 13089 12447
rect 13119 12473 13145 12479
rect 13119 12441 13145 12447
rect 13567 12473 13593 12479
rect 13567 12441 13593 12447
rect 7799 12417 7825 12423
rect 7799 12385 7825 12391
rect 13511 12417 13537 12423
rect 13511 12385 13537 12391
rect 13679 12417 13705 12423
rect 13679 12385 13705 12391
rect 7575 12361 7601 12367
rect 2137 12335 2143 12361
rect 2169 12335 2175 12361
rect 7401 12335 7407 12361
rect 7433 12335 7439 12361
rect 7575 12329 7601 12335
rect 7911 12361 7937 12367
rect 7911 12329 7937 12335
rect 8695 12361 8721 12367
rect 8695 12329 8721 12335
rect 8807 12361 8833 12367
rect 8807 12329 8833 12335
rect 9087 12361 9113 12367
rect 9087 12329 9113 12335
rect 9255 12361 9281 12367
rect 12615 12361 12641 12367
rect 9753 12335 9759 12361
rect 9785 12335 9791 12361
rect 9255 12329 9281 12335
rect 12615 12329 12641 12335
rect 12727 12361 12753 12367
rect 12727 12329 12753 12335
rect 12951 12361 12977 12367
rect 12951 12329 12977 12335
rect 13175 12361 13201 12367
rect 13337 12335 13343 12361
rect 13369 12335 13375 12361
rect 18937 12335 18943 12361
rect 18969 12335 18975 12361
rect 13175 12329 13201 12335
rect 6001 12279 6007 12305
rect 6033 12279 6039 12305
rect 7065 12279 7071 12305
rect 7097 12279 7103 12305
rect 12217 12279 12223 12305
rect 12249 12279 12255 12305
rect 967 12249 993 12255
rect 967 12217 993 12223
rect 20007 12249 20033 12255
rect 20007 12217 20033 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 20007 12025 20033 12031
rect 20007 11993 20033 11999
rect 7463 11969 7489 11975
rect 7463 11937 7489 11943
rect 7575 11969 7601 11975
rect 7575 11937 7601 11943
rect 7687 11969 7713 11975
rect 7687 11937 7713 11943
rect 7911 11969 7937 11975
rect 8801 11943 8807 11969
rect 8833 11943 8839 11969
rect 18825 11943 18831 11969
rect 18857 11943 18863 11969
rect 7911 11937 7937 11943
rect 7295 11913 7321 11919
rect 7295 11881 7321 11887
rect 7351 11913 7377 11919
rect 7351 11881 7377 11887
rect 7743 11857 7769 11863
rect 7743 11825 7769 11831
rect 8695 11857 8721 11863
rect 8695 11825 8721 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 9647 11689 9673 11695
rect 9137 11663 9143 11689
rect 9169 11663 9175 11689
rect 9647 11657 9673 11663
rect 7799 11633 7825 11639
rect 9591 11633 9617 11639
rect 8969 11607 8975 11633
rect 9001 11607 9007 11633
rect 9361 11607 9367 11633
rect 9393 11607 9399 11633
rect 12049 11607 12055 11633
rect 12081 11607 12087 11633
rect 7799 11601 7825 11607
rect 9591 11601 9617 11607
rect 7463 11577 7489 11583
rect 2137 11551 2143 11577
rect 2169 11551 2175 11577
rect 7177 11551 7183 11577
rect 7209 11551 7215 11577
rect 7463 11545 7489 11551
rect 7687 11577 7713 11583
rect 9417 11551 9423 11577
rect 9449 11551 9455 11577
rect 10313 11551 10319 11577
rect 10345 11551 10351 11577
rect 11937 11551 11943 11577
rect 11969 11551 11975 11577
rect 18825 11551 18831 11577
rect 18857 11551 18863 11577
rect 7687 11545 7713 11551
rect 7575 11521 7601 11527
rect 12279 11521 12305 11527
rect 5721 11495 5727 11521
rect 5753 11495 5759 11521
rect 6785 11495 6791 11521
rect 6817 11495 6823 11521
rect 10649 11495 10655 11521
rect 10681 11495 10687 11521
rect 11713 11495 11719 11521
rect 11745 11495 11751 11521
rect 7575 11489 7601 11495
rect 12279 11489 12305 11495
rect 967 11465 993 11471
rect 967 11433 993 11439
rect 9647 11465 9673 11471
rect 9647 11433 9673 11439
rect 20007 11465 20033 11471
rect 20007 11433 20033 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 8527 11297 8553 11303
rect 8527 11265 8553 11271
rect 8807 11297 8833 11303
rect 8807 11265 8833 11271
rect 9535 11297 9561 11303
rect 9535 11265 9561 11271
rect 7631 11241 7657 11247
rect 7631 11209 7657 11215
rect 10991 11241 11017 11247
rect 10991 11209 11017 11215
rect 11159 11241 11185 11247
rect 11159 11209 11185 11215
rect 11495 11241 11521 11247
rect 13959 11241 13985 11247
rect 13337 11215 13343 11241
rect 13369 11215 13375 11241
rect 11495 11209 11521 11215
rect 13959 11209 13985 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 7463 11185 7489 11191
rect 10935 11185 10961 11191
rect 8577 11159 8583 11185
rect 8609 11159 8615 11185
rect 8969 11159 8975 11185
rect 9001 11159 9007 11185
rect 9809 11159 9815 11185
rect 9841 11159 9847 11185
rect 10313 11159 10319 11185
rect 10345 11159 10351 11185
rect 7463 11153 7489 11159
rect 10935 11153 10961 11159
rect 11271 11185 11297 11191
rect 13455 11185 13481 11191
rect 11601 11159 11607 11185
rect 11633 11159 11639 11185
rect 11937 11159 11943 11185
rect 11969 11159 11975 11185
rect 11271 11153 11297 11159
rect 13455 11153 13481 11159
rect 13679 11185 13705 11191
rect 14625 11159 14631 11185
rect 14657 11159 14663 11185
rect 14961 11159 14967 11185
rect 14993 11159 14999 11185
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 13679 11153 13705 11159
rect 7295 11129 7321 11135
rect 7295 11097 7321 11103
rect 7351 11129 7377 11135
rect 7351 11097 7377 11103
rect 8471 11129 8497 11135
rect 8471 11097 8497 11103
rect 9087 11129 9113 11135
rect 9087 11097 9113 11103
rect 11439 11129 11465 11135
rect 13791 11129 13817 11135
rect 12273 11103 12279 11129
rect 12305 11103 12311 11129
rect 11439 11097 11465 11103
rect 13791 11097 13817 11103
rect 14015 11129 14041 11135
rect 14015 11097 14041 11103
rect 8695 11073 8721 11079
rect 8695 11041 8721 11047
rect 8863 11073 8889 11079
rect 8863 11041 8889 11047
rect 9591 11073 9617 11079
rect 9591 11041 9617 11047
rect 9703 11073 9729 11079
rect 11047 11073 11073 11079
rect 10201 11047 10207 11073
rect 10233 11047 10239 11073
rect 9703 11041 9729 11047
rect 11047 11041 11073 11047
rect 13623 11073 13649 11079
rect 14737 11047 14743 11073
rect 14769 11047 14775 11073
rect 15073 11047 15079 11073
rect 15105 11047 15111 11073
rect 13623 11041 13649 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 8191 10905 8217 10911
rect 8191 10873 8217 10879
rect 9087 10905 9113 10911
rect 9087 10873 9113 10879
rect 10039 10905 10065 10911
rect 10039 10873 10065 10879
rect 10151 10905 10177 10911
rect 10151 10873 10177 10879
rect 11327 10905 11353 10911
rect 11327 10873 11353 10879
rect 11551 10905 11577 10911
rect 11551 10873 11577 10879
rect 12783 10905 12809 10911
rect 12783 10873 12809 10879
rect 7911 10849 7937 10855
rect 12055 10849 12081 10855
rect 6505 10823 6511 10849
rect 6537 10823 6543 10849
rect 8857 10823 8863 10849
rect 8889 10823 8895 10849
rect 7911 10817 7937 10823
rect 12055 10817 12081 10823
rect 12111 10849 12137 10855
rect 12111 10817 12137 10823
rect 12839 10849 12865 10855
rect 13617 10823 13623 10849
rect 13649 10823 13655 10849
rect 12839 10817 12865 10823
rect 7967 10793 7993 10799
rect 6169 10767 6175 10793
rect 6201 10767 6207 10793
rect 7967 10761 7993 10767
rect 8695 10793 8721 10799
rect 8695 10761 8721 10767
rect 9031 10793 9057 10799
rect 9031 10761 9057 10767
rect 9983 10793 10009 10799
rect 9983 10761 10009 10767
rect 11495 10793 11521 10799
rect 11495 10761 11521 10767
rect 11607 10793 11633 10799
rect 11607 10761 11633 10767
rect 11831 10793 11857 10799
rect 11831 10761 11857 10767
rect 11943 10793 11969 10799
rect 12671 10793 12697 10799
rect 12329 10767 12335 10793
rect 12361 10767 12367 10793
rect 11943 10761 11969 10767
rect 12671 10761 12697 10767
rect 13063 10793 13089 10799
rect 13225 10767 13231 10793
rect 13257 10767 13263 10793
rect 18825 10767 18831 10793
rect 18857 10767 18863 10793
rect 13063 10761 13089 10767
rect 20007 10737 20033 10743
rect 7569 10711 7575 10737
rect 7601 10711 7607 10737
rect 12105 10711 12111 10737
rect 12137 10711 12143 10737
rect 14681 10711 14687 10737
rect 14713 10711 14719 10737
rect 20007 10705 20033 10711
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 20007 10457 20033 10463
rect 20007 10425 20033 10431
rect 18825 10375 18831 10401
rect 18857 10375 18863 10401
rect 10817 10319 10823 10345
rect 10849 10319 10855 10345
rect 11153 10319 11159 10345
rect 11185 10319 11191 10345
rect 7127 10289 7153 10295
rect 7127 10257 7153 10263
rect 10655 10289 10681 10295
rect 10655 10257 10681 10263
rect 11327 10289 11353 10295
rect 11327 10257 11353 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 12559 10065 12585 10071
rect 8185 10039 8191 10065
rect 8217 10039 8223 10065
rect 9529 10039 9535 10065
rect 9561 10039 9567 10065
rect 10705 10039 10711 10065
rect 10737 10039 10743 10065
rect 12559 10033 12585 10039
rect 12671 10065 12697 10071
rect 12671 10033 12697 10039
rect 8359 10009 8385 10015
rect 2137 9983 2143 10009
rect 2169 9983 2175 10009
rect 6953 9983 6959 10009
rect 6985 9983 6991 10009
rect 7569 9983 7575 10009
rect 7601 9983 7607 10009
rect 8359 9977 8385 9983
rect 8695 10009 8721 10015
rect 9367 10009 9393 10015
rect 12727 10009 12753 10015
rect 8969 9983 8975 10009
rect 9001 9983 9007 10009
rect 9697 9983 9703 10009
rect 9729 9983 9735 10009
rect 8695 9977 8721 9983
rect 9367 9977 9393 9983
rect 12727 9977 12753 9983
rect 7799 9953 7825 9959
rect 5497 9927 5503 9953
rect 5529 9927 5535 9953
rect 6561 9927 6567 9953
rect 6593 9927 6599 9953
rect 7401 9927 7407 9953
rect 7433 9927 7439 9953
rect 7799 9921 7825 9927
rect 9199 9953 9225 9959
rect 9199 9921 9225 9927
rect 12951 9953 12977 9959
rect 12951 9921 12977 9927
rect 967 9897 993 9903
rect 967 9865 993 9871
rect 8807 9897 8833 9903
rect 8807 9865 8833 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 6343 9729 6369 9735
rect 6343 9697 6369 9703
rect 8807 9729 8833 9735
rect 8807 9697 8833 9703
rect 9087 9729 9113 9735
rect 9087 9697 9113 9703
rect 9311 9729 9337 9735
rect 9311 9697 9337 9703
rect 10207 9729 10233 9735
rect 10207 9697 10233 9703
rect 13007 9729 13033 9735
rect 13007 9697 13033 9703
rect 20007 9673 20033 9679
rect 12329 9647 12335 9673
rect 12361 9647 12367 9673
rect 20007 9641 20033 9647
rect 7911 9617 7937 9623
rect 7457 9591 7463 9617
rect 7489 9591 7495 9617
rect 7911 9585 7937 9591
rect 8527 9617 8553 9623
rect 8527 9585 8553 9591
rect 9143 9617 9169 9623
rect 9871 9617 9897 9623
rect 13119 9617 13145 9623
rect 13343 9617 13369 9623
rect 9473 9591 9479 9617
rect 9505 9591 9511 9617
rect 10929 9591 10935 9617
rect 10961 9591 10967 9617
rect 13281 9591 13287 9617
rect 13313 9591 13319 9617
rect 9143 9585 9169 9591
rect 9871 9585 9897 9591
rect 13119 9585 13145 9591
rect 13343 9585 13369 9591
rect 14239 9617 14265 9623
rect 18825 9591 18831 9617
rect 18857 9591 18863 9617
rect 14239 9585 14265 9591
rect 6287 9561 6313 9567
rect 6287 9529 6313 9535
rect 7127 9561 7153 9567
rect 7127 9529 7153 9535
rect 7183 9561 7209 9567
rect 7183 9529 7209 9535
rect 7239 9561 7265 9567
rect 8359 9561 8385 9567
rect 7737 9535 7743 9561
rect 7769 9535 7775 9561
rect 7239 9529 7265 9535
rect 8359 9529 8385 9535
rect 9927 9561 9953 9567
rect 9927 9529 9953 9535
rect 10151 9561 10177 9567
rect 11265 9535 11271 9561
rect 11297 9535 11303 9561
rect 10151 9529 10177 9535
rect 7071 9505 7097 9511
rect 7071 9473 7097 9479
rect 8415 9505 8441 9511
rect 8415 9473 8441 9479
rect 8695 9505 8721 9511
rect 8695 9473 8721 9479
rect 8751 9505 8777 9511
rect 8751 9473 8777 9479
rect 9087 9505 9113 9511
rect 9087 9473 9113 9479
rect 9367 9505 9393 9511
rect 9367 9473 9393 9479
rect 10039 9505 10065 9511
rect 10039 9473 10065 9479
rect 10207 9505 10233 9511
rect 10207 9473 10233 9479
rect 12671 9505 12697 9511
rect 13399 9505 13425 9511
rect 12833 9479 12839 9505
rect 12865 9479 12871 9505
rect 12671 9473 12697 9479
rect 13399 9473 13425 9479
rect 13455 9505 13481 9511
rect 13455 9473 13481 9479
rect 14183 9505 14209 9511
rect 14183 9473 14209 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 11159 9337 11185 9343
rect 11159 9305 11185 9311
rect 11383 9337 11409 9343
rect 11383 9305 11409 9311
rect 7407 9281 7433 9287
rect 7407 9249 7433 9255
rect 7575 9281 7601 9287
rect 7575 9249 7601 9255
rect 8415 9281 8441 9287
rect 9591 9281 9617 9287
rect 11215 9281 11241 9287
rect 9137 9255 9143 9281
rect 9169 9255 9175 9281
rect 10593 9255 10599 9281
rect 10625 9255 10631 9281
rect 8415 9249 8441 9255
rect 9591 9249 9617 9255
rect 11215 9249 11241 9255
rect 12615 9281 12641 9287
rect 12615 9249 12641 9255
rect 8247 9225 8273 9231
rect 8247 9193 8273 9199
rect 8975 9225 9001 9231
rect 8975 9193 9001 9199
rect 9255 9225 9281 9231
rect 9255 9193 9281 9199
rect 9479 9225 9505 9231
rect 9479 9193 9505 9199
rect 9983 9225 10009 9231
rect 9983 9193 10009 9199
rect 10095 9225 10121 9231
rect 10095 9193 10121 9199
rect 10767 9225 10793 9231
rect 10767 9193 10793 9199
rect 10935 9225 10961 9231
rect 10935 9193 10961 9199
rect 11103 9225 11129 9231
rect 11103 9193 11129 9199
rect 11551 9225 11577 9231
rect 11551 9193 11577 9199
rect 11887 9225 11913 9231
rect 13063 9225 13089 9231
rect 11993 9199 11999 9225
rect 12025 9199 12031 9225
rect 12721 9199 12727 9225
rect 12753 9199 12759 9225
rect 13225 9199 13231 9225
rect 13257 9199 13263 9225
rect 13617 9199 13623 9225
rect 13649 9199 13655 9225
rect 11887 9193 11913 9199
rect 13063 9193 13089 9199
rect 9535 9169 9561 9175
rect 9535 9137 9561 9143
rect 12279 9169 12305 9175
rect 14681 9143 14687 9169
rect 14713 9143 14719 9169
rect 12279 9137 12305 9143
rect 10257 9087 10263 9113
rect 10289 9087 10295 9113
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 11887 8945 11913 8951
rect 11887 8913 11913 8919
rect 12223 8945 12249 8951
rect 12223 8913 12249 8919
rect 967 8889 993 8895
rect 11943 8889 11969 8895
rect 14631 8889 14657 8895
rect 7681 8863 7687 8889
rect 7713 8863 7719 8889
rect 14289 8863 14295 8889
rect 14321 8863 14327 8889
rect 967 8857 993 8863
rect 11943 8857 11969 8863
rect 14631 8857 14657 8863
rect 20007 8889 20033 8895
rect 20007 8857 20033 8863
rect 7351 8833 7377 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 7351 8801 7377 8807
rect 7575 8833 7601 8839
rect 10095 8833 10121 8839
rect 12559 8833 12585 8839
rect 7737 8807 7743 8833
rect 7769 8807 7775 8833
rect 7849 8807 7855 8833
rect 7881 8807 7887 8833
rect 8913 8807 8919 8833
rect 8945 8807 8951 8833
rect 11545 8807 11551 8833
rect 11577 8807 11583 8833
rect 12889 8807 12895 8833
rect 12921 8807 12927 8833
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 7575 8801 7601 8807
rect 10095 8801 10121 8807
rect 12559 8801 12585 8807
rect 10151 8777 10177 8783
rect 10823 8777 10849 8783
rect 12111 8777 12137 8783
rect 10649 8751 10655 8777
rect 10681 8751 10687 8777
rect 11433 8751 11439 8777
rect 11465 8751 11471 8777
rect 10151 8745 10177 8751
rect 10823 8745 10849 8751
rect 12111 8745 12137 8751
rect 12727 8777 12753 8783
rect 13225 8751 13231 8777
rect 13257 8751 13263 8777
rect 12727 8745 12753 8751
rect 7239 8721 7265 8727
rect 7239 8689 7265 8695
rect 7295 8721 7321 8727
rect 7295 8689 7321 8695
rect 7967 8721 7993 8727
rect 7967 8689 7993 8695
rect 8079 8721 8105 8727
rect 9535 8721 9561 8727
rect 10263 8721 10289 8727
rect 12615 8721 12641 8727
rect 9025 8695 9031 8721
rect 9057 8695 9063 8721
rect 9697 8695 9703 8721
rect 9729 8695 9735 8721
rect 12385 8695 12391 8721
rect 12417 8695 12423 8721
rect 8079 8689 8105 8695
rect 9535 8689 9561 8695
rect 10263 8689 10289 8695
rect 12615 8689 12641 8695
rect 14575 8721 14601 8727
rect 14575 8689 14601 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 7631 8553 7657 8559
rect 7631 8521 7657 8527
rect 7855 8553 7881 8559
rect 7855 8521 7881 8527
rect 13343 8553 13369 8559
rect 13343 8521 13369 8527
rect 13399 8553 13425 8559
rect 13399 8521 13425 8527
rect 13455 8553 13481 8559
rect 13455 8521 13481 8527
rect 6337 8471 6343 8497
rect 6369 8471 6375 8497
rect 7799 8441 7825 8447
rect 6001 8415 6007 8441
rect 6033 8415 6039 8441
rect 7799 8409 7825 8415
rect 7911 8441 7937 8447
rect 7911 8409 7937 8415
rect 8023 8441 8049 8447
rect 12671 8441 12697 8447
rect 9809 8415 9815 8441
rect 9841 8415 9847 8441
rect 8023 8409 8049 8415
rect 12671 8409 12697 8415
rect 13007 8441 13033 8447
rect 13007 8409 13033 8415
rect 13119 8385 13145 8391
rect 7401 8359 7407 8385
rect 7433 8359 7439 8385
rect 12105 8359 12111 8385
rect 12137 8359 12143 8385
rect 13119 8353 13145 8359
rect 13231 8385 13257 8391
rect 13231 8353 13257 8359
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 8415 8105 8441 8111
rect 7121 8079 7127 8105
rect 7153 8079 7159 8105
rect 8185 8079 8191 8105
rect 8217 8079 8223 8105
rect 8415 8073 8441 8079
rect 12111 8105 12137 8111
rect 12111 8073 12137 8079
rect 10823 8049 10849 8055
rect 6785 8023 6791 8049
rect 6817 8023 6823 8049
rect 10823 8017 10849 8023
rect 11551 8049 11577 8055
rect 11551 8017 11577 8023
rect 11775 8049 11801 8055
rect 11775 8017 11801 8023
rect 11887 8049 11913 8055
rect 11887 8017 11913 8023
rect 9647 7993 9673 7999
rect 9647 7961 9673 7967
rect 9703 7993 9729 7999
rect 9703 7961 9729 7967
rect 12055 7993 12081 7999
rect 12055 7961 12081 7967
rect 9535 7937 9561 7943
rect 11831 7937 11857 7943
rect 10649 7911 10655 7937
rect 10681 7911 10687 7937
rect 9535 7905 9561 7911
rect 11831 7905 11857 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 9087 7769 9113 7775
rect 9087 7737 9113 7743
rect 9815 7769 9841 7775
rect 9815 7737 9841 7743
rect 10375 7769 10401 7775
rect 11999 7769 12025 7775
rect 11825 7743 11831 7769
rect 11857 7743 11863 7769
rect 10375 7737 10401 7743
rect 11999 7737 12025 7743
rect 12615 7769 12641 7775
rect 12615 7737 12641 7743
rect 12727 7769 12753 7775
rect 12727 7737 12753 7743
rect 8975 7713 9001 7719
rect 8975 7681 9001 7687
rect 9143 7713 9169 7719
rect 9143 7681 9169 7687
rect 10431 7713 10457 7719
rect 10431 7681 10457 7687
rect 10487 7713 10513 7719
rect 10487 7681 10513 7687
rect 10879 7713 10905 7719
rect 10879 7681 10905 7687
rect 11047 7713 11073 7719
rect 11047 7681 11073 7687
rect 13007 7713 13033 7719
rect 13007 7681 13033 7687
rect 13119 7713 13145 7719
rect 13119 7681 13145 7687
rect 13175 7713 13201 7719
rect 13175 7681 13201 7687
rect 9255 7657 9281 7663
rect 9255 7625 9281 7631
rect 9927 7657 9953 7663
rect 9927 7625 9953 7631
rect 10151 7657 10177 7663
rect 10151 7625 10177 7631
rect 10319 7657 10345 7663
rect 12951 7657 12977 7663
rect 10705 7631 10711 7657
rect 10737 7631 10743 7657
rect 10319 7625 10345 7631
rect 12951 7625 12977 7631
rect 9871 7601 9897 7607
rect 9871 7569 9897 7575
rect 12223 7601 12249 7607
rect 12223 7569 12249 7575
rect 12671 7601 12697 7607
rect 12671 7569 12697 7575
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 8969 7295 8975 7321
rect 9001 7295 9007 7321
rect 9249 7295 9255 7321
rect 9281 7295 9287 7321
rect 11041 7295 11047 7321
rect 11073 7295 11079 7321
rect 12105 7295 12111 7321
rect 12137 7295 12143 7321
rect 12665 7295 12671 7321
rect 12697 7295 12703 7321
rect 13729 7295 13735 7321
rect 13761 7295 13767 7321
rect 9367 7265 9393 7271
rect 9647 7265 9673 7271
rect 7569 7239 7575 7265
rect 7601 7239 7607 7265
rect 7905 7239 7911 7265
rect 7937 7239 7943 7265
rect 9137 7239 9143 7265
rect 9169 7239 9175 7265
rect 9473 7239 9479 7265
rect 9505 7239 9511 7265
rect 9921 7239 9927 7265
rect 9953 7239 9959 7265
rect 10649 7239 10655 7265
rect 10681 7239 10687 7265
rect 12273 7239 12279 7265
rect 12305 7239 12311 7265
rect 9367 7233 9393 7239
rect 9647 7233 9673 7239
rect 9255 7153 9281 7159
rect 9255 7121 9281 7127
rect 9703 7153 9729 7159
rect 9703 7121 9729 7127
rect 9759 7153 9785 7159
rect 9759 7121 9785 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 9255 6985 9281 6991
rect 9255 6953 9281 6959
rect 11159 6985 11185 6991
rect 11159 6953 11185 6959
rect 12111 6985 12137 6991
rect 12111 6953 12137 6959
rect 8919 6929 8945 6935
rect 8919 6897 8945 6903
rect 9031 6929 9057 6935
rect 9865 6903 9871 6929
rect 9897 6903 9903 6929
rect 9031 6897 9057 6903
rect 9473 6847 9479 6873
rect 9505 6847 9511 6873
rect 10929 6791 10935 6817
rect 10961 6791 10967 6817
rect 8863 6761 8889 6767
rect 8863 6729 8889 6735
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 9479 6537 9505 6543
rect 8129 6511 8135 6537
rect 8161 6511 8167 6537
rect 9193 6511 9199 6537
rect 9225 6511 9231 6537
rect 9479 6505 9505 6511
rect 7737 6455 7743 6481
rect 7769 6455 7775 6481
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 9529 2143 9535 2169
rect 9561 2143 9567 2169
rect 13225 2143 13231 2169
rect 13257 2143 13263 2169
rect 10039 2057 10065 2063
rect 10039 2025 10065 2031
rect 13735 2057 13761 2063
rect 13735 2025 13761 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 9311 1833 9337 1839
rect 9311 1801 9337 1807
rect 11047 1833 11073 1839
rect 11047 1801 11073 1807
rect 8801 1751 8807 1777
rect 8833 1751 8839 1777
rect 10537 1751 10543 1777
rect 10569 1751 10575 1777
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 12783 19111 12809 19137
rect 9423 19055 9449 19081
rect 11103 19055 11129 19081
rect 9871 18999 9897 19025
rect 11999 18999 12025 19025
rect 12279 18999 12305 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 10375 18719 10401 18745
rect 9871 18607 9897 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9591 18327 9617 18353
rect 9199 18215 9225 18241
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 9927 13903 9953 13929
rect 18943 13903 18969 13929
rect 10263 13847 10289 13873
rect 11327 13847 11353 13873
rect 11607 13847 11633 13873
rect 19951 13847 19977 13873
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 9871 13567 9897 13593
rect 10711 13567 10737 13593
rect 20007 13567 20033 13593
rect 8471 13511 8497 13537
rect 10935 13511 10961 13537
rect 11047 13511 11073 13537
rect 18831 13511 18857 13537
rect 8807 13455 8833 13481
rect 10767 13455 10793 13481
rect 11159 13455 11185 13481
rect 11215 13455 11241 13481
rect 13175 13455 13201 13481
rect 13231 13455 13257 13481
rect 10095 13399 10121 13425
rect 10655 13399 10681 13425
rect 12559 13399 12585 13425
rect 13343 13399 13369 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 7519 13231 7545 13257
rect 9087 13231 9113 13257
rect 9759 13231 9785 13257
rect 9143 13175 9169 13201
rect 9815 13175 9841 13201
rect 14519 13175 14545 13201
rect 7295 13119 7321 13145
rect 8639 13119 8665 13145
rect 8863 13119 8889 13145
rect 8975 13119 9001 13145
rect 9255 13119 9281 13145
rect 9423 13119 9449 13145
rect 10487 13119 10513 13145
rect 12727 13119 12753 13145
rect 14407 13119 14433 13145
rect 18831 13119 18857 13145
rect 5839 13063 5865 13089
rect 6903 13063 6929 13089
rect 8919 13063 8945 13089
rect 10823 13063 10849 13089
rect 11887 13063 11913 13089
rect 12111 13063 12137 13089
rect 12335 13063 12361 13089
rect 13119 13063 13145 13089
rect 14183 13063 14209 13089
rect 19951 13063 19977 13089
rect 9759 13007 9785 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 967 12783 993 12809
rect 8247 12783 8273 12809
rect 9311 12783 9337 12809
rect 9871 12783 9897 12809
rect 13735 12783 13761 12809
rect 20007 12783 20033 12809
rect 2143 12727 2169 12753
rect 7463 12727 7489 12753
rect 7911 12727 7937 12753
rect 9479 12727 9505 12753
rect 11047 12727 11073 12753
rect 11327 12727 11353 12753
rect 11439 12727 11465 12753
rect 11607 12727 11633 12753
rect 12279 12727 12305 12753
rect 13959 12727 13985 12753
rect 18831 12727 18857 12753
rect 9647 12671 9673 12697
rect 11943 12671 11969 12697
rect 12671 12671 12697 12697
rect 7519 12615 7545 12641
rect 7631 12615 7657 12641
rect 10991 12615 11017 12641
rect 11103 12615 11129 12641
rect 11551 12615 11577 12641
rect 12111 12615 12137 12641
rect 14071 12615 14097 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 7687 12447 7713 12473
rect 8135 12447 8161 12473
rect 8975 12447 9001 12473
rect 9199 12447 9225 12473
rect 12671 12447 12697 12473
rect 13063 12447 13089 12473
rect 13119 12447 13145 12473
rect 13567 12447 13593 12473
rect 7799 12391 7825 12417
rect 13511 12391 13537 12417
rect 13679 12391 13705 12417
rect 2143 12335 2169 12361
rect 7407 12335 7433 12361
rect 7575 12335 7601 12361
rect 7911 12335 7937 12361
rect 8695 12335 8721 12361
rect 8807 12335 8833 12361
rect 9087 12335 9113 12361
rect 9255 12335 9281 12361
rect 9759 12335 9785 12361
rect 12615 12335 12641 12361
rect 12727 12335 12753 12361
rect 12951 12335 12977 12361
rect 13175 12335 13201 12361
rect 13343 12335 13369 12361
rect 18943 12335 18969 12361
rect 6007 12279 6033 12305
rect 7071 12279 7097 12305
rect 12223 12279 12249 12305
rect 967 12223 993 12249
rect 20007 12223 20033 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 20007 11999 20033 12025
rect 7463 11943 7489 11969
rect 7575 11943 7601 11969
rect 7687 11943 7713 11969
rect 7911 11943 7937 11969
rect 8807 11943 8833 11969
rect 18831 11943 18857 11969
rect 7295 11887 7321 11913
rect 7351 11887 7377 11913
rect 7743 11831 7769 11857
rect 8695 11831 8721 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 9143 11663 9169 11689
rect 9647 11663 9673 11689
rect 7799 11607 7825 11633
rect 8975 11607 9001 11633
rect 9367 11607 9393 11633
rect 9591 11607 9617 11633
rect 12055 11607 12081 11633
rect 2143 11551 2169 11577
rect 7183 11551 7209 11577
rect 7463 11551 7489 11577
rect 7687 11551 7713 11577
rect 9423 11551 9449 11577
rect 10319 11551 10345 11577
rect 11943 11551 11969 11577
rect 18831 11551 18857 11577
rect 5727 11495 5753 11521
rect 6791 11495 6817 11521
rect 7575 11495 7601 11521
rect 10655 11495 10681 11521
rect 11719 11495 11745 11521
rect 12279 11495 12305 11521
rect 967 11439 993 11465
rect 9647 11439 9673 11465
rect 20007 11439 20033 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 8527 11271 8553 11297
rect 8807 11271 8833 11297
rect 9535 11271 9561 11297
rect 7631 11215 7657 11241
rect 10991 11215 11017 11241
rect 11159 11215 11185 11241
rect 11495 11215 11521 11241
rect 13343 11215 13369 11241
rect 13959 11215 13985 11241
rect 20007 11215 20033 11241
rect 7463 11159 7489 11185
rect 8583 11159 8609 11185
rect 8975 11159 9001 11185
rect 9815 11159 9841 11185
rect 10319 11159 10345 11185
rect 10935 11159 10961 11185
rect 11271 11159 11297 11185
rect 11607 11159 11633 11185
rect 11943 11159 11969 11185
rect 13455 11159 13481 11185
rect 13679 11159 13705 11185
rect 14631 11159 14657 11185
rect 14967 11159 14993 11185
rect 18831 11159 18857 11185
rect 7295 11103 7321 11129
rect 7351 11103 7377 11129
rect 8471 11103 8497 11129
rect 9087 11103 9113 11129
rect 11439 11103 11465 11129
rect 12279 11103 12305 11129
rect 13791 11103 13817 11129
rect 14015 11103 14041 11129
rect 8695 11047 8721 11073
rect 8863 11047 8889 11073
rect 9591 11047 9617 11073
rect 9703 11047 9729 11073
rect 10207 11047 10233 11073
rect 11047 11047 11073 11073
rect 13623 11047 13649 11073
rect 14743 11047 14769 11073
rect 15079 11047 15105 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 8191 10879 8217 10905
rect 9087 10879 9113 10905
rect 10039 10879 10065 10905
rect 10151 10879 10177 10905
rect 11327 10879 11353 10905
rect 11551 10879 11577 10905
rect 12783 10879 12809 10905
rect 6511 10823 6537 10849
rect 7911 10823 7937 10849
rect 8863 10823 8889 10849
rect 12055 10823 12081 10849
rect 12111 10823 12137 10849
rect 12839 10823 12865 10849
rect 13623 10823 13649 10849
rect 6175 10767 6201 10793
rect 7967 10767 7993 10793
rect 8695 10767 8721 10793
rect 9031 10767 9057 10793
rect 9983 10767 10009 10793
rect 11495 10767 11521 10793
rect 11607 10767 11633 10793
rect 11831 10767 11857 10793
rect 11943 10767 11969 10793
rect 12335 10767 12361 10793
rect 12671 10767 12697 10793
rect 13063 10767 13089 10793
rect 13231 10767 13257 10793
rect 18831 10767 18857 10793
rect 7575 10711 7601 10737
rect 12111 10711 12137 10737
rect 14687 10711 14713 10737
rect 20007 10711 20033 10737
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 20007 10431 20033 10457
rect 18831 10375 18857 10401
rect 10823 10319 10849 10345
rect 11159 10319 11185 10345
rect 7127 10263 7153 10289
rect 10655 10263 10681 10289
rect 11327 10263 11353 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 8191 10039 8217 10065
rect 9535 10039 9561 10065
rect 10711 10039 10737 10065
rect 12559 10039 12585 10065
rect 12671 10039 12697 10065
rect 2143 9983 2169 10009
rect 6959 9983 6985 10009
rect 7575 9983 7601 10009
rect 8359 9983 8385 10009
rect 8695 9983 8721 10009
rect 8975 9983 9001 10009
rect 9367 9983 9393 10009
rect 9703 9983 9729 10009
rect 12727 9983 12753 10009
rect 5503 9927 5529 9953
rect 6567 9927 6593 9953
rect 7407 9927 7433 9953
rect 7799 9927 7825 9953
rect 9199 9927 9225 9953
rect 12951 9927 12977 9953
rect 967 9871 993 9897
rect 8807 9871 8833 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 6343 9703 6369 9729
rect 8807 9703 8833 9729
rect 9087 9703 9113 9729
rect 9311 9703 9337 9729
rect 10207 9703 10233 9729
rect 13007 9703 13033 9729
rect 12335 9647 12361 9673
rect 20007 9647 20033 9673
rect 7463 9591 7489 9617
rect 7911 9591 7937 9617
rect 8527 9591 8553 9617
rect 9143 9591 9169 9617
rect 9479 9591 9505 9617
rect 9871 9591 9897 9617
rect 10935 9591 10961 9617
rect 13119 9591 13145 9617
rect 13287 9591 13313 9617
rect 13343 9591 13369 9617
rect 14239 9591 14265 9617
rect 18831 9591 18857 9617
rect 6287 9535 6313 9561
rect 7127 9535 7153 9561
rect 7183 9535 7209 9561
rect 7239 9535 7265 9561
rect 7743 9535 7769 9561
rect 8359 9535 8385 9561
rect 9927 9535 9953 9561
rect 10151 9535 10177 9561
rect 11271 9535 11297 9561
rect 7071 9479 7097 9505
rect 8415 9479 8441 9505
rect 8695 9479 8721 9505
rect 8751 9479 8777 9505
rect 9087 9479 9113 9505
rect 9367 9479 9393 9505
rect 10039 9479 10065 9505
rect 10207 9479 10233 9505
rect 12671 9479 12697 9505
rect 12839 9479 12865 9505
rect 13399 9479 13425 9505
rect 13455 9479 13481 9505
rect 14183 9479 14209 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 11159 9311 11185 9337
rect 11383 9311 11409 9337
rect 7407 9255 7433 9281
rect 7575 9255 7601 9281
rect 8415 9255 8441 9281
rect 9143 9255 9169 9281
rect 9591 9255 9617 9281
rect 10599 9255 10625 9281
rect 11215 9255 11241 9281
rect 12615 9255 12641 9281
rect 8247 9199 8273 9225
rect 8975 9199 9001 9225
rect 9255 9199 9281 9225
rect 9479 9199 9505 9225
rect 9983 9199 10009 9225
rect 10095 9199 10121 9225
rect 10767 9199 10793 9225
rect 10935 9199 10961 9225
rect 11103 9199 11129 9225
rect 11551 9199 11577 9225
rect 11887 9199 11913 9225
rect 11999 9199 12025 9225
rect 12727 9199 12753 9225
rect 13063 9199 13089 9225
rect 13231 9199 13257 9225
rect 13623 9199 13649 9225
rect 9535 9143 9561 9169
rect 12279 9143 12305 9169
rect 14687 9143 14713 9169
rect 10263 9087 10289 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 11887 8919 11913 8945
rect 12223 8919 12249 8945
rect 967 8863 993 8889
rect 7687 8863 7713 8889
rect 11943 8863 11969 8889
rect 14295 8863 14321 8889
rect 14631 8863 14657 8889
rect 20007 8863 20033 8889
rect 2143 8807 2169 8833
rect 7351 8807 7377 8833
rect 7575 8807 7601 8833
rect 7743 8807 7769 8833
rect 7855 8807 7881 8833
rect 8919 8807 8945 8833
rect 10095 8807 10121 8833
rect 11551 8807 11577 8833
rect 12559 8807 12585 8833
rect 12895 8807 12921 8833
rect 18831 8807 18857 8833
rect 10151 8751 10177 8777
rect 10655 8751 10681 8777
rect 10823 8751 10849 8777
rect 11439 8751 11465 8777
rect 12111 8751 12137 8777
rect 12727 8751 12753 8777
rect 13231 8751 13257 8777
rect 7239 8695 7265 8721
rect 7295 8695 7321 8721
rect 7967 8695 7993 8721
rect 8079 8695 8105 8721
rect 9031 8695 9057 8721
rect 9535 8695 9561 8721
rect 9703 8695 9729 8721
rect 10263 8695 10289 8721
rect 12391 8695 12417 8721
rect 12615 8695 12641 8721
rect 14575 8695 14601 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7631 8527 7657 8553
rect 7855 8527 7881 8553
rect 13343 8527 13369 8553
rect 13399 8527 13425 8553
rect 13455 8527 13481 8553
rect 6343 8471 6369 8497
rect 6007 8415 6033 8441
rect 7799 8415 7825 8441
rect 7911 8415 7937 8441
rect 8023 8415 8049 8441
rect 9815 8415 9841 8441
rect 12671 8415 12697 8441
rect 13007 8415 13033 8441
rect 7407 8359 7433 8385
rect 12111 8359 12137 8385
rect 13119 8359 13145 8385
rect 13231 8359 13257 8385
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 7127 8079 7153 8105
rect 8191 8079 8217 8105
rect 8415 8079 8441 8105
rect 12111 8079 12137 8105
rect 6791 8023 6817 8049
rect 10823 8023 10849 8049
rect 11551 8023 11577 8049
rect 11775 8023 11801 8049
rect 11887 8023 11913 8049
rect 9647 7967 9673 7993
rect 9703 7967 9729 7993
rect 12055 7967 12081 7993
rect 9535 7911 9561 7937
rect 10655 7911 10681 7937
rect 11831 7911 11857 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 9087 7743 9113 7769
rect 9815 7743 9841 7769
rect 10375 7743 10401 7769
rect 11831 7743 11857 7769
rect 11999 7743 12025 7769
rect 12615 7743 12641 7769
rect 12727 7743 12753 7769
rect 8975 7687 9001 7713
rect 9143 7687 9169 7713
rect 10431 7687 10457 7713
rect 10487 7687 10513 7713
rect 10879 7687 10905 7713
rect 11047 7687 11073 7713
rect 13007 7687 13033 7713
rect 13119 7687 13145 7713
rect 13175 7687 13201 7713
rect 9255 7631 9281 7657
rect 9927 7631 9953 7657
rect 10151 7631 10177 7657
rect 10319 7631 10345 7657
rect 10711 7631 10737 7657
rect 12951 7631 12977 7657
rect 9871 7575 9897 7601
rect 12223 7575 12249 7601
rect 12671 7575 12697 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 8975 7295 9001 7321
rect 9255 7295 9281 7321
rect 11047 7295 11073 7321
rect 12111 7295 12137 7321
rect 12671 7295 12697 7321
rect 13735 7295 13761 7321
rect 7575 7239 7601 7265
rect 7911 7239 7937 7265
rect 9143 7239 9169 7265
rect 9367 7239 9393 7265
rect 9479 7239 9505 7265
rect 9647 7239 9673 7265
rect 9927 7239 9953 7265
rect 10655 7239 10681 7265
rect 12279 7239 12305 7265
rect 9255 7127 9281 7153
rect 9703 7127 9729 7153
rect 9759 7127 9785 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 9255 6959 9281 6985
rect 11159 6959 11185 6985
rect 12111 6959 12137 6985
rect 8919 6903 8945 6929
rect 9031 6903 9057 6929
rect 9871 6903 9897 6929
rect 9479 6847 9505 6873
rect 10935 6791 10961 6817
rect 8863 6735 8889 6761
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 8135 6511 8161 6537
rect 9199 6511 9225 6537
rect 9479 6511 9505 6537
rect 7743 6455 7769 6481
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 9535 2143 9561 2169
rect 13231 2143 13257 2169
rect 10039 2031 10065 2057
rect 13735 2031 13761 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 9311 1807 9337 1833
rect 11047 1807 11073 1833
rect 8807 1751 8833 1777
rect 10543 1751 10569 1777
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 9072 20600 9128 21000
rect 9408 20600 9464 21000
rect 9744 20600 9800 21000
rect 11088 20600 11144 21000
rect 11760 20600 11816 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 9086 18354 9114 20600
rect 9422 19081 9450 20600
rect 9758 19306 9786 20600
rect 9758 19273 9786 19278
rect 10374 19306 10402 19311
rect 9422 19055 9423 19081
rect 9449 19055 9450 19081
rect 9422 19049 9450 19055
rect 9870 19026 9898 19031
rect 9646 19025 9898 19026
rect 9646 18999 9871 19025
rect 9897 18999 9898 19025
rect 9646 18998 9898 18999
rect 9086 18321 9114 18326
rect 9590 18354 9618 18359
rect 9590 18307 9618 18326
rect 9198 18241 9226 18247
rect 9198 18215 9199 18241
rect 9225 18215 9226 18241
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 8470 13538 8498 13543
rect 8470 13491 8498 13510
rect 2086 13482 2114 13487
rect 966 12809 994 12815
rect 966 12783 967 12809
rect 993 12783 994 12809
rect 966 12474 994 12783
rect 966 12441 994 12446
rect 966 12250 994 12255
rect 966 12203 994 12222
rect 966 11466 994 11471
rect 966 11419 994 11438
rect 2086 9954 2114 13454
rect 8806 13481 8834 13487
rect 8806 13455 8807 13481
rect 8833 13455 8834 13481
rect 7518 13426 7546 13431
rect 7518 13258 7546 13398
rect 7294 13257 7546 13258
rect 7294 13231 7519 13257
rect 7545 13231 7546 13257
rect 7294 13230 7546 13231
rect 7294 13145 7322 13230
rect 7518 13225 7546 13230
rect 7910 13426 7938 13431
rect 7294 13119 7295 13145
rect 7321 13119 7322 13145
rect 7294 13113 7322 13119
rect 2142 13090 2170 13095
rect 2142 12753 2170 13062
rect 5838 13090 5866 13095
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 2142 12727 2143 12753
rect 2169 12727 2170 12753
rect 2142 12721 2170 12727
rect 5838 12698 5866 13062
rect 5838 12665 5866 12670
rect 6902 13089 6930 13095
rect 6902 13063 6903 13089
rect 6929 13063 6930 13089
rect 6902 12586 6930 13063
rect 6902 12553 6930 12558
rect 7294 12782 7490 12810
rect 2142 12362 2170 12367
rect 2142 12315 2170 12334
rect 6006 12362 6034 12367
rect 6006 12305 6034 12334
rect 6006 12279 6007 12305
rect 6033 12279 6034 12305
rect 6006 12273 6034 12279
rect 7070 12306 7098 12311
rect 7070 12259 7098 12278
rect 7182 12250 7210 12255
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 2142 11578 2170 11583
rect 2142 11531 2170 11550
rect 6174 11578 6202 11583
rect 5726 11522 5754 11527
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 5726 11130 5754 11494
rect 5726 11097 5754 11102
rect 6174 10793 6202 11550
rect 7182 11578 7210 12222
rect 7182 11531 7210 11550
rect 7294 11913 7322 12782
rect 7462 12753 7490 12782
rect 7462 12727 7463 12753
rect 7489 12727 7490 12753
rect 7462 12721 7490 12727
rect 7910 12754 7938 13398
rect 8806 13258 8834 13455
rect 9198 13426 9226 18215
rect 9646 15974 9674 18998
rect 9870 18993 9898 18998
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 10374 18745 10402 19278
rect 11102 19081 11130 20600
rect 11774 19138 11802 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 12782 19138 12810 19143
rect 11774 19105 11802 19110
rect 11830 19110 12082 19138
rect 11102 19055 11103 19081
rect 11129 19055 11130 19081
rect 11102 19049 11130 19055
rect 10374 18719 10375 18745
rect 10401 18719 10402 18745
rect 10374 18713 10402 18719
rect 9870 18634 9898 18639
rect 9590 15946 9674 15974
rect 9814 18633 9898 18634
rect 9814 18607 9871 18633
rect 9897 18607 9898 18633
rect 9814 18606 9898 18607
rect 9198 13398 9338 13426
rect 9086 13258 9114 13263
rect 8806 13257 9114 13258
rect 8806 13231 9087 13257
rect 9113 13231 9114 13257
rect 8806 13230 9114 13231
rect 9086 13225 9114 13230
rect 9142 13201 9170 13207
rect 9142 13175 9143 13201
rect 9169 13175 9170 13201
rect 8638 13146 8666 13151
rect 8862 13146 8890 13151
rect 8246 13090 8274 13095
rect 8246 12809 8274 13062
rect 8246 12783 8247 12809
rect 8273 12783 8274 12809
rect 8246 12777 8274 12783
rect 7910 12753 8162 12754
rect 7910 12727 7911 12753
rect 7937 12727 8162 12753
rect 7910 12726 8162 12727
rect 7910 12721 7938 12726
rect 7294 11887 7295 11913
rect 7321 11887 7322 11913
rect 6790 11522 6818 11527
rect 6790 11475 6818 11494
rect 7294 11129 7322 11887
rect 7350 12698 7378 12703
rect 7350 11913 7378 12670
rect 7518 12641 7546 12647
rect 7518 12615 7519 12641
rect 7545 12615 7546 12641
rect 7518 12474 7546 12615
rect 7518 12441 7546 12446
rect 7630 12641 7658 12647
rect 7630 12615 7631 12641
rect 7657 12615 7658 12641
rect 7406 12361 7434 12367
rect 7406 12335 7407 12361
rect 7433 12335 7434 12361
rect 7406 12250 7434 12335
rect 7574 12361 7602 12367
rect 7574 12335 7575 12361
rect 7601 12335 7602 12361
rect 7574 12306 7602 12335
rect 7406 12217 7434 12222
rect 7462 12278 7602 12306
rect 7462 11969 7490 12278
rect 7462 11943 7463 11969
rect 7489 11943 7490 11969
rect 7462 11937 7490 11943
rect 7574 12138 7602 12143
rect 7574 11969 7602 12110
rect 7574 11943 7575 11969
rect 7601 11943 7602 11969
rect 7574 11937 7602 11943
rect 7630 11970 7658 12615
rect 7686 12586 7714 12591
rect 7686 12473 7714 12558
rect 7686 12447 7687 12473
rect 7713 12447 7714 12473
rect 7686 12441 7714 12447
rect 8134 12473 8162 12726
rect 8638 12474 8666 13118
rect 8134 12447 8135 12473
rect 8161 12447 8162 12473
rect 7798 12418 7826 12423
rect 7798 12371 7826 12390
rect 7910 12362 7938 12367
rect 7742 12306 7770 12311
rect 7686 11970 7714 11975
rect 7630 11969 7714 11970
rect 7630 11943 7687 11969
rect 7713 11943 7714 11969
rect 7630 11942 7714 11943
rect 7686 11937 7714 11942
rect 7350 11887 7351 11913
rect 7377 11887 7378 11913
rect 7350 11881 7378 11887
rect 7742 11857 7770 12278
rect 7910 12138 7938 12334
rect 7742 11831 7743 11857
rect 7769 11831 7770 11857
rect 7742 11825 7770 11831
rect 7798 12110 7910 12138
rect 7798 11633 7826 12110
rect 7910 12105 7938 12110
rect 8134 12250 8162 12447
rect 7798 11607 7799 11633
rect 7825 11607 7826 11633
rect 7798 11601 7826 11607
rect 7910 11969 7938 11975
rect 7910 11943 7911 11969
rect 7937 11943 7938 11969
rect 7462 11577 7490 11583
rect 7462 11551 7463 11577
rect 7489 11551 7490 11577
rect 7462 11185 7490 11551
rect 7518 11578 7546 11583
rect 7518 11410 7546 11550
rect 7686 11577 7714 11583
rect 7686 11551 7687 11577
rect 7713 11551 7714 11577
rect 7574 11522 7602 11527
rect 7574 11475 7602 11494
rect 7518 11382 7658 11410
rect 7630 11241 7658 11382
rect 7686 11354 7714 11551
rect 7686 11321 7714 11326
rect 7910 11298 7938 11943
rect 7910 11265 7938 11270
rect 7630 11215 7631 11241
rect 7657 11215 7658 11241
rect 7630 11209 7658 11215
rect 7462 11159 7463 11185
rect 7489 11159 7490 11185
rect 7462 11153 7490 11159
rect 7294 11103 7295 11129
rect 7321 11103 7322 11129
rect 6510 10850 6538 10855
rect 6510 10803 6538 10822
rect 6174 10767 6175 10793
rect 6201 10767 6202 10793
rect 6174 10761 6202 10767
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 7126 10289 7154 10295
rect 7126 10263 7127 10289
rect 7153 10263 7154 10289
rect 7126 10094 7154 10263
rect 7294 10094 7322 11103
rect 7350 11130 7378 11135
rect 7350 11083 7378 11102
rect 8134 10906 8162 12222
rect 8526 12446 8666 12474
rect 8750 13145 8890 13146
rect 8750 13119 8863 13145
rect 8889 13119 8890 13145
rect 8750 13118 8890 13119
rect 8526 11297 8554 12446
rect 8694 12418 8722 12423
rect 8694 12361 8722 12390
rect 8694 12335 8695 12361
rect 8721 12335 8722 12361
rect 8694 12329 8722 12335
rect 8750 12362 8778 13118
rect 8862 13113 8890 13118
rect 8974 13145 9002 13151
rect 8974 13119 8975 13145
rect 9001 13119 9002 13145
rect 8918 13090 8946 13095
rect 8918 13043 8946 13062
rect 8974 12473 9002 13119
rect 8974 12447 8975 12473
rect 9001 12447 9002 12473
rect 8974 12441 9002 12447
rect 9142 12418 9170 13175
rect 9254 13146 9282 13151
rect 9254 13099 9282 13118
rect 9310 12810 9338 13398
rect 9422 13146 9450 13151
rect 9422 13099 9450 13118
rect 9198 12809 9506 12810
rect 9198 12783 9311 12809
rect 9337 12783 9506 12809
rect 9198 12782 9506 12783
rect 9198 12473 9226 12782
rect 9310 12777 9338 12782
rect 9478 12753 9506 12782
rect 9478 12727 9479 12753
rect 9505 12727 9506 12753
rect 9478 12721 9506 12727
rect 9590 12698 9618 15946
rect 9814 13594 9842 18606
rect 9870 18601 9898 18606
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 11326 14266 11354 14271
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9926 13929 9954 13935
rect 9926 13903 9927 13929
rect 9953 13903 9954 13929
rect 9870 13594 9898 13599
rect 9758 13593 9898 13594
rect 9758 13567 9871 13593
rect 9897 13567 9898 13593
rect 9758 13566 9898 13567
rect 9758 13257 9786 13566
rect 9870 13561 9898 13566
rect 9926 13538 9954 13903
rect 10262 13874 10290 13879
rect 11326 13874 11354 14238
rect 10262 13873 10738 13874
rect 10262 13847 10263 13873
rect 10289 13847 10738 13873
rect 10262 13846 10738 13847
rect 10262 13841 10290 13846
rect 10710 13593 10738 13846
rect 10710 13567 10711 13593
rect 10737 13567 10738 13593
rect 10710 13561 10738 13567
rect 11158 13873 11354 13874
rect 11158 13847 11327 13873
rect 11353 13847 11354 13873
rect 11158 13846 11354 13847
rect 9926 13426 9954 13510
rect 10934 13538 10962 13543
rect 11046 13538 11074 13543
rect 10934 13537 11074 13538
rect 10934 13511 10935 13537
rect 10961 13511 11047 13537
rect 11073 13511 11074 13537
rect 10934 13510 11074 13511
rect 10934 13505 10962 13510
rect 11046 13505 11074 13510
rect 10766 13481 10794 13487
rect 10766 13455 10767 13481
rect 10793 13455 10794 13481
rect 10094 13426 10122 13431
rect 9926 13398 10094 13426
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9758 13231 9759 13257
rect 9785 13231 9786 13257
rect 9758 13225 9786 13231
rect 9814 13202 9842 13207
rect 9814 13155 9842 13174
rect 9702 13146 9730 13151
rect 10094 13146 10122 13398
rect 10486 13426 10514 13431
rect 10486 13146 10514 13398
rect 10654 13426 10682 13431
rect 10654 13425 10738 13426
rect 10654 13399 10655 13425
rect 10681 13399 10738 13425
rect 10654 13398 10738 13399
rect 10654 13393 10682 13398
rect 9730 13118 9786 13146
rect 9702 13113 9730 13118
rect 9758 13033 9786 13118
rect 9758 13007 9759 13033
rect 9785 13007 9786 13033
rect 9758 13001 9786 13007
rect 9870 13118 10122 13146
rect 10318 13145 10514 13146
rect 10318 13119 10487 13145
rect 10513 13119 10514 13145
rect 10318 13118 10514 13119
rect 9870 12809 9898 13118
rect 9870 12783 9871 12809
rect 9897 12783 9898 12809
rect 9870 12777 9898 12783
rect 9646 12698 9674 12703
rect 9590 12697 9674 12698
rect 9590 12671 9647 12697
rect 9673 12671 9674 12697
rect 9590 12670 9674 12671
rect 9646 12665 9674 12670
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9198 12447 9199 12473
rect 9225 12447 9226 12473
rect 9198 12441 9226 12447
rect 8750 12138 8778 12334
rect 8806 12362 8834 12367
rect 9086 12362 9114 12367
rect 8806 12361 9114 12362
rect 8806 12335 8807 12361
rect 8833 12335 9087 12361
rect 9113 12335 9114 12361
rect 8806 12334 9114 12335
rect 8806 12329 8834 12334
rect 9086 12329 9114 12334
rect 8750 12110 8890 12138
rect 8806 11970 8834 11975
rect 8526 11271 8527 11297
rect 8553 11271 8554 11297
rect 8526 11265 8554 11271
rect 8582 11969 8834 11970
rect 8582 11943 8807 11969
rect 8833 11943 8834 11969
rect 8582 11942 8834 11943
rect 8582 11185 8610 11942
rect 8806 11937 8834 11942
rect 8694 11858 8722 11863
rect 8862 11858 8890 12110
rect 8694 11857 8890 11858
rect 8694 11831 8695 11857
rect 8721 11831 8890 11857
rect 8694 11830 8890 11831
rect 8694 11825 8722 11830
rect 8974 11690 9002 11695
rect 8974 11634 9002 11662
rect 9142 11689 9170 12390
rect 9254 12362 9282 12367
rect 9702 12362 9730 12367
rect 9254 12361 9506 12362
rect 9254 12335 9255 12361
rect 9281 12335 9506 12361
rect 9254 12334 9506 12335
rect 9254 12329 9282 12334
rect 9142 11663 9143 11689
rect 9169 11663 9170 11689
rect 9142 11657 9170 11663
rect 9086 11634 9114 11639
rect 8918 11633 9002 11634
rect 8918 11607 8975 11633
rect 9001 11607 9002 11633
rect 8918 11606 9002 11607
rect 8806 11298 8834 11303
rect 8806 11251 8834 11270
rect 8582 11159 8583 11185
rect 8609 11159 8610 11185
rect 8470 11129 8498 11135
rect 8470 11103 8471 11129
rect 8497 11103 8498 11129
rect 8190 10906 8218 10911
rect 8134 10905 8218 10906
rect 8134 10879 8191 10905
rect 8217 10879 8218 10905
rect 8134 10878 8218 10879
rect 8190 10873 8218 10878
rect 7910 10850 7938 10855
rect 7910 10803 7938 10822
rect 6958 10066 7154 10094
rect 7238 10066 7322 10094
rect 7574 10794 7602 10799
rect 7574 10737 7602 10766
rect 7966 10794 7994 10799
rect 7966 10747 7994 10766
rect 7574 10711 7575 10737
rect 7601 10711 7602 10737
rect 2142 10010 2170 10015
rect 2142 9963 2170 9982
rect 5502 10010 5530 10015
rect 2086 9921 2114 9926
rect 5502 9953 5530 9982
rect 6958 10009 6986 10066
rect 6958 9983 6959 10009
rect 6985 9983 6986 10009
rect 6566 9954 6594 9959
rect 5502 9927 5503 9953
rect 5529 9927 5530 9953
rect 966 9898 994 9903
rect 966 9851 994 9870
rect 5502 9842 5530 9927
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 5502 9809 5530 9814
rect 6342 9953 6594 9954
rect 6342 9927 6567 9953
rect 6593 9927 6594 9953
rect 6342 9926 6594 9927
rect 2238 9781 2370 9786
rect 6342 9729 6370 9926
rect 6566 9921 6594 9926
rect 6342 9703 6343 9729
rect 6369 9703 6370 9729
rect 6342 9697 6370 9703
rect 6286 9562 6314 9567
rect 6286 9515 6314 9534
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 966 8889 994 8895
rect 966 8863 967 8889
rect 993 8863 994 8889
rect 966 8442 994 8863
rect 2142 8834 2170 8839
rect 2142 8787 2170 8806
rect 6958 8554 6986 9983
rect 7182 9842 7210 9847
rect 7126 9562 7154 9567
rect 7126 9515 7154 9534
rect 7182 9561 7210 9814
rect 7182 9535 7183 9561
rect 7209 9535 7210 9561
rect 7182 9529 7210 9535
rect 7238 9562 7266 10066
rect 7574 10009 7602 10711
rect 8470 10094 8498 11103
rect 7574 9983 7575 10009
rect 7601 9983 7602 10009
rect 7574 9977 7602 9983
rect 8190 10066 8498 10094
rect 8190 10065 8218 10066
rect 8190 10039 8191 10065
rect 8217 10039 8218 10065
rect 7238 9515 7266 9534
rect 7406 9953 7434 9959
rect 7798 9954 7826 9959
rect 7406 9927 7407 9953
rect 7433 9927 7434 9953
rect 7070 9505 7098 9511
rect 7070 9479 7071 9505
rect 7097 9479 7098 9505
rect 7070 9114 7098 9479
rect 7406 9506 7434 9927
rect 7630 9953 7826 9954
rect 7630 9927 7799 9953
rect 7825 9927 7826 9953
rect 7630 9926 7826 9927
rect 7462 9730 7490 9735
rect 7462 9617 7490 9702
rect 7462 9591 7463 9617
rect 7489 9591 7490 9617
rect 7462 9585 7490 9591
rect 7406 9478 7490 9506
rect 7406 9281 7434 9287
rect 7406 9255 7407 9281
rect 7433 9255 7434 9281
rect 7070 9081 7098 9086
rect 7350 9114 7378 9119
rect 7350 8833 7378 9086
rect 7350 8807 7351 8833
rect 7377 8807 7378 8833
rect 7350 8801 7378 8807
rect 7406 8834 7434 9255
rect 7238 8722 7266 8727
rect 7238 8675 7266 8694
rect 7294 8721 7322 8727
rect 7294 8695 7295 8721
rect 7321 8695 7322 8721
rect 6790 8526 6958 8554
rect 6342 8498 6370 8503
rect 6342 8451 6370 8470
rect 966 8409 994 8414
rect 6006 8442 6034 8447
rect 6006 8395 6034 8414
rect 6790 8442 6818 8526
rect 6958 8521 6986 8526
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 6790 8049 6818 8414
rect 7126 8106 7154 8111
rect 7294 8106 7322 8695
rect 7406 8498 7434 8806
rect 7406 8465 7434 8470
rect 7462 9226 7490 9478
rect 7574 9282 7602 9287
rect 7630 9282 7658 9926
rect 7798 9921 7826 9926
rect 7910 9674 7938 9679
rect 7910 9617 7938 9646
rect 7910 9591 7911 9617
rect 7937 9591 7938 9617
rect 7910 9585 7938 9591
rect 7742 9562 7770 9567
rect 7742 9515 7770 9534
rect 8078 9506 8106 9511
rect 7574 9281 7658 9282
rect 7574 9255 7575 9281
rect 7601 9255 7658 9281
rect 7574 9254 7658 9255
rect 8022 9478 8078 9506
rect 7574 9249 7602 9254
rect 7406 8386 7434 8391
rect 7462 8386 7490 9198
rect 7742 9114 7770 9119
rect 7686 8890 7714 8895
rect 7574 8889 7714 8890
rect 7574 8863 7687 8889
rect 7713 8863 7714 8889
rect 7574 8862 7714 8863
rect 7574 8833 7602 8862
rect 7686 8857 7714 8862
rect 7574 8807 7575 8833
rect 7601 8807 7602 8833
rect 7574 8801 7602 8807
rect 7742 8833 7770 9086
rect 7742 8807 7743 8833
rect 7769 8807 7770 8833
rect 7742 8801 7770 8807
rect 7854 8834 7882 8839
rect 7854 8787 7882 8806
rect 7910 8778 7938 8783
rect 7854 8722 7882 8727
rect 7518 8554 7546 8559
rect 7630 8554 7658 8559
rect 7546 8553 7658 8554
rect 7546 8527 7631 8553
rect 7657 8527 7658 8553
rect 7546 8526 7658 8527
rect 7518 8521 7546 8526
rect 7406 8385 7490 8386
rect 7406 8359 7407 8385
rect 7433 8359 7490 8385
rect 7406 8358 7490 8359
rect 7406 8353 7434 8358
rect 7126 8105 7322 8106
rect 7126 8079 7127 8105
rect 7153 8079 7322 8105
rect 7126 8078 7322 8079
rect 7574 8106 7602 8526
rect 7630 8521 7658 8526
rect 7854 8553 7882 8694
rect 7854 8527 7855 8553
rect 7881 8527 7882 8553
rect 7854 8521 7882 8527
rect 7126 8073 7154 8078
rect 6790 8023 6791 8049
rect 6817 8023 6818 8049
rect 6790 8017 6818 8023
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 7574 7266 7602 8078
rect 7798 8441 7826 8447
rect 7798 8415 7799 8441
rect 7825 8415 7826 8441
rect 7798 8386 7826 8415
rect 7910 8442 7938 8750
rect 7966 8721 7994 8727
rect 7966 8695 7967 8721
rect 7993 8695 7994 8721
rect 7966 8554 7994 8695
rect 7966 8521 7994 8526
rect 7910 8441 7994 8442
rect 7910 8415 7911 8441
rect 7937 8415 7994 8441
rect 7910 8414 7994 8415
rect 7910 8409 7938 8414
rect 7798 7714 7826 8358
rect 7966 8330 7994 8414
rect 8022 8441 8050 9478
rect 8078 9473 8106 9478
rect 8022 8415 8023 8441
rect 8049 8415 8050 8441
rect 8022 8409 8050 8415
rect 8078 8722 8106 8727
rect 8190 8722 8218 10039
rect 8358 10009 8386 10015
rect 8358 9983 8359 10009
rect 8385 9983 8386 10009
rect 8358 9674 8386 9983
rect 8358 9641 8386 9646
rect 8526 9618 8554 9623
rect 8526 9571 8554 9590
rect 8358 9561 8386 9567
rect 8358 9535 8359 9561
rect 8385 9535 8386 9561
rect 8358 9282 8386 9535
rect 8582 9562 8610 11159
rect 8694 11074 8722 11079
rect 8694 11027 8722 11046
rect 8862 11073 8890 11079
rect 8862 11047 8863 11073
rect 8889 11047 8890 11073
rect 8862 10962 8890 11047
rect 8862 10929 8890 10934
rect 8862 10850 8890 10855
rect 8918 10850 8946 11606
rect 8974 11601 9002 11606
rect 9030 11606 9086 11634
rect 8974 11186 9002 11191
rect 9030 11186 9058 11606
rect 9086 11601 9114 11606
rect 9366 11634 9394 11639
rect 9366 11587 9394 11606
rect 9422 11578 9450 11583
rect 9422 11531 9450 11550
rect 8974 11185 9058 11186
rect 8974 11159 8975 11185
rect 9001 11159 9058 11185
rect 8974 11158 9058 11159
rect 8974 11153 9002 11158
rect 9030 11074 9058 11158
rect 9086 11130 9114 11135
rect 9086 11083 9114 11102
rect 9030 10906 9058 11046
rect 9478 10962 9506 12334
rect 9646 11690 9674 11695
rect 9646 11643 9674 11662
rect 9590 11634 9618 11639
rect 9590 11587 9618 11606
rect 9646 11466 9674 11471
rect 9702 11466 9730 12334
rect 9646 11465 9730 11466
rect 9646 11439 9647 11465
rect 9673 11439 9730 11465
rect 9646 11438 9730 11439
rect 9758 12361 9786 12367
rect 9758 12335 9759 12361
rect 9785 12335 9786 12361
rect 9646 11433 9674 11438
rect 9534 11354 9562 11359
rect 9534 11297 9562 11326
rect 9534 11271 9535 11297
rect 9561 11271 9562 11297
rect 9534 11265 9562 11271
rect 9590 11074 9618 11079
rect 9702 11074 9730 11079
rect 9590 11027 9618 11046
rect 9646 11073 9730 11074
rect 9646 11047 9703 11073
rect 9729 11047 9730 11073
rect 9646 11046 9730 11047
rect 9478 10934 9618 10962
rect 9086 10906 9114 10911
rect 9030 10905 9114 10906
rect 9030 10879 9087 10905
rect 9113 10879 9114 10905
rect 9030 10878 9114 10879
rect 9086 10873 9114 10878
rect 8750 10849 8946 10850
rect 8750 10823 8863 10849
rect 8889 10823 8946 10849
rect 8750 10822 8946 10823
rect 8694 10794 8722 10799
rect 8694 10009 8722 10766
rect 8694 9983 8695 10009
rect 8721 9983 8722 10009
rect 8694 9977 8722 9983
rect 8750 9618 8778 10822
rect 8862 10817 8890 10822
rect 9030 10793 9058 10799
rect 9030 10767 9031 10793
rect 9057 10767 9058 10793
rect 8974 10010 9002 10015
rect 8974 9963 9002 9982
rect 8806 9898 8834 9903
rect 9030 9898 9058 10767
rect 9534 10122 9562 10127
rect 9534 10065 9562 10094
rect 9534 10039 9535 10065
rect 9561 10039 9562 10065
rect 9534 10033 9562 10039
rect 9366 10010 9394 10015
rect 9198 9954 9226 9959
rect 9198 9907 9226 9926
rect 8806 9897 9058 9898
rect 8806 9871 8807 9897
rect 8833 9871 9058 9897
rect 8806 9870 9058 9871
rect 8806 9865 8834 9870
rect 8806 9786 8834 9791
rect 8806 9729 8834 9758
rect 8806 9703 8807 9729
rect 8833 9703 8834 9729
rect 8806 9697 8834 9703
rect 8582 9529 8610 9534
rect 8638 9590 8778 9618
rect 8414 9506 8442 9511
rect 8414 9505 8498 9506
rect 8414 9479 8415 9505
rect 8441 9479 8498 9505
rect 8414 9478 8498 9479
rect 8414 9473 8442 9478
rect 8470 9450 8498 9478
rect 8638 9450 8666 9590
rect 8470 9422 8666 9450
rect 8694 9505 8722 9511
rect 8694 9479 8695 9505
rect 8721 9479 8722 9505
rect 8414 9282 8442 9287
rect 8358 9254 8414 9282
rect 8414 9235 8442 9254
rect 8246 9226 8274 9231
rect 8246 9179 8274 9198
rect 8078 8721 8218 8722
rect 8078 8695 8079 8721
rect 8105 8695 8218 8721
rect 8078 8694 8218 8695
rect 8470 8722 8498 9422
rect 8694 9282 8722 9479
rect 8750 9506 8778 9511
rect 8750 9459 8778 9478
rect 8806 9338 8834 9343
rect 8862 9338 8890 9870
rect 9086 9730 9114 9735
rect 8834 9310 8890 9338
rect 9030 9702 9086 9730
rect 8806 9305 8834 9310
rect 8694 9226 8722 9254
rect 9030 9282 9058 9702
rect 9086 9683 9114 9702
rect 9310 9730 9338 9735
rect 9366 9730 9394 9982
rect 9310 9729 9394 9730
rect 9310 9703 9311 9729
rect 9337 9703 9394 9729
rect 9310 9702 9394 9703
rect 9590 9786 9618 10934
rect 9310 9697 9338 9702
rect 9478 9674 9506 9679
rect 9142 9618 9170 9623
rect 9170 9590 9226 9618
rect 9142 9571 9170 9590
rect 9086 9506 9114 9511
rect 9086 9459 9114 9478
rect 9030 9249 9058 9254
rect 9142 9281 9170 9287
rect 9142 9255 9143 9281
rect 9169 9255 9170 9281
rect 8974 9226 9002 9231
rect 8694 9225 9002 9226
rect 8694 9199 8975 9225
rect 9001 9199 9002 9225
rect 8694 9198 9002 9199
rect 8918 8833 8946 9198
rect 8974 9193 9002 9198
rect 9142 9226 9170 9255
rect 9198 9226 9226 9590
rect 9478 9617 9506 9646
rect 9478 9591 9479 9617
rect 9505 9591 9506 9617
rect 9366 9505 9394 9511
rect 9366 9479 9367 9505
rect 9393 9479 9394 9505
rect 9254 9226 9282 9231
rect 9198 9225 9282 9226
rect 9198 9199 9255 9225
rect 9281 9199 9282 9225
rect 9198 9198 9282 9199
rect 9142 9193 9170 9198
rect 9254 9193 9282 9198
rect 8918 8807 8919 8833
rect 8945 8807 8946 8833
rect 8918 8801 8946 8807
rect 9366 9058 9394 9479
rect 9478 9338 9506 9591
rect 9478 9305 9506 9310
rect 9590 9281 9618 9758
rect 9590 9255 9591 9281
rect 9617 9255 9618 9281
rect 8078 8442 8106 8694
rect 8470 8689 8498 8694
rect 9030 8721 9058 8727
rect 9030 8695 9031 8721
rect 9057 8695 9058 8721
rect 9030 8554 9058 8695
rect 9030 8521 9058 8526
rect 8078 8409 8106 8414
rect 9366 8330 9394 9030
rect 9478 9226 9506 9231
rect 9478 8778 9506 9198
rect 9534 9169 9562 9175
rect 9534 9143 9535 9169
rect 9561 9143 9562 9169
rect 9534 8834 9562 9143
rect 9590 9170 9618 9255
rect 9646 10794 9674 11046
rect 9702 11041 9730 11046
rect 9758 10850 9786 12335
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9814 11578 9842 11583
rect 9814 11242 9842 11550
rect 10318 11577 10346 13118
rect 10486 13113 10514 13118
rect 10318 11551 10319 11577
rect 10345 11551 10346 11577
rect 10318 11545 10346 11551
rect 10654 11521 10682 11527
rect 10654 11495 10655 11521
rect 10681 11495 10682 11521
rect 9814 11185 9842 11214
rect 9814 11159 9815 11185
rect 9841 11159 9842 11185
rect 9814 11153 9842 11159
rect 10318 11242 10346 11247
rect 10318 11185 10346 11214
rect 10654 11242 10682 11495
rect 10710 11242 10738 13398
rect 10766 12642 10794 13455
rect 11158 13481 11186 13846
rect 11326 13841 11354 13846
rect 11606 13874 11634 13879
rect 11158 13455 11159 13481
rect 11185 13455 11186 13481
rect 11158 13449 11186 13455
rect 11214 13481 11242 13487
rect 11214 13455 11215 13481
rect 11241 13455 11242 13481
rect 11214 13426 11242 13455
rect 11606 13482 11634 13846
rect 11606 13449 11634 13454
rect 11214 13393 11242 13398
rect 11550 13426 11578 13431
rect 10822 13090 10850 13095
rect 10822 13089 11074 13090
rect 10822 13063 10823 13089
rect 10849 13063 11074 13089
rect 10822 13062 11074 13063
rect 10822 13057 10850 13062
rect 11046 12753 11074 13062
rect 11046 12727 11047 12753
rect 11073 12727 11074 12753
rect 11046 12721 11074 12727
rect 11326 12754 11354 12759
rect 11438 12754 11466 12759
rect 11326 12753 11466 12754
rect 11326 12727 11327 12753
rect 11353 12727 11439 12753
rect 11465 12727 11466 12753
rect 11326 12726 11466 12727
rect 11550 12754 11578 13398
rect 11830 13090 11858 19110
rect 11998 19025 12026 19031
rect 11998 18999 11999 19025
rect 12025 18999 12026 19025
rect 11998 14266 12026 18999
rect 12054 19026 12082 19110
rect 12782 19091 12810 19110
rect 12278 19026 12306 19031
rect 12054 19025 12306 19026
rect 12054 18999 12279 19025
rect 12305 18999 12306 19025
rect 12054 18998 12306 18999
rect 12278 18993 12306 18998
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 11998 14233 12026 14238
rect 18942 13929 18970 13935
rect 18942 13903 18943 13929
rect 18969 13903 18970 13929
rect 12110 13874 12138 13879
rect 11886 13090 11914 13095
rect 11830 13089 11914 13090
rect 11830 13063 11887 13089
rect 11913 13063 11914 13089
rect 11830 13062 11914 13063
rect 11606 12754 11634 12759
rect 11550 12726 11606 12754
rect 11326 12721 11354 12726
rect 11438 12721 11466 12726
rect 11606 12707 11634 12726
rect 10766 12609 10794 12614
rect 10990 12641 11018 12647
rect 10990 12615 10991 12641
rect 11017 12615 11018 12641
rect 10990 12474 11018 12615
rect 10990 12441 11018 12446
rect 11046 12642 11074 12647
rect 11102 12642 11130 12647
rect 11074 12641 11130 12642
rect 11074 12615 11103 12641
rect 11129 12615 11130 12641
rect 11074 12614 11130 12615
rect 10990 11242 11018 11247
rect 10710 11214 10962 11242
rect 10654 11209 10682 11214
rect 10318 11159 10319 11185
rect 10345 11159 10346 11185
rect 10206 11074 10234 11079
rect 10206 11027 10234 11046
rect 10150 11018 10178 11023
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 10038 10906 10066 10911
rect 10038 10859 10066 10878
rect 10150 10905 10178 10990
rect 10150 10879 10151 10905
rect 10177 10879 10178 10905
rect 10150 10873 10178 10879
rect 9758 10822 9842 10850
rect 9646 9226 9674 10766
rect 9814 10066 9842 10822
rect 9982 10794 10010 10799
rect 9982 10747 10010 10766
rect 10318 10346 10346 11159
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9702 10009 9730 10015
rect 9702 9983 9703 10009
rect 9729 9983 9730 10009
rect 9702 9954 9730 9983
rect 9702 9921 9730 9926
rect 9646 9193 9674 9198
rect 9590 9137 9618 9142
rect 9534 8806 9786 8834
rect 9478 8745 9506 8750
rect 9534 8722 9562 8727
rect 9702 8722 9730 8727
rect 9534 8675 9562 8694
rect 9646 8721 9730 8722
rect 9646 8695 9703 8721
rect 9729 8695 9730 8721
rect 9646 8694 9730 8695
rect 7966 8302 8218 8330
rect 8190 8105 8218 8302
rect 9254 8302 9394 8330
rect 8190 8079 8191 8105
rect 8217 8079 8218 8105
rect 8190 8073 8218 8079
rect 8414 8106 8442 8111
rect 8414 8059 8442 8078
rect 9030 7854 9170 7882
rect 7798 7681 7826 7686
rect 8974 7714 9002 7719
rect 8974 7667 9002 7686
rect 8974 7322 9002 7327
rect 9030 7322 9058 7854
rect 8806 7321 9058 7322
rect 8806 7295 8975 7321
rect 9001 7295 9058 7321
rect 8806 7294 9058 7295
rect 9086 7769 9114 7775
rect 9086 7743 9087 7769
rect 9113 7743 9114 7769
rect 7910 7266 7938 7271
rect 7574 7265 7770 7266
rect 7574 7239 7575 7265
rect 7601 7239 7770 7265
rect 7574 7238 7770 7239
rect 7574 7233 7602 7238
rect 7742 6986 7770 7238
rect 7910 7219 7938 7238
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 7742 6481 7770 6958
rect 8134 6762 8162 6767
rect 8134 6537 8162 6734
rect 8134 6511 8135 6537
rect 8161 6511 8162 6537
rect 8134 6505 8162 6511
rect 7742 6455 7743 6481
rect 7769 6455 7770 6481
rect 7742 6449 7770 6455
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8806 1777 8834 7294
rect 8974 7289 9002 7294
rect 9086 7266 9114 7743
rect 9142 7713 9170 7854
rect 9142 7687 9143 7713
rect 9169 7687 9170 7713
rect 9142 7681 9170 7687
rect 9254 7658 9282 8302
rect 9646 7994 9674 8694
rect 9702 8689 9730 8694
rect 9646 7947 9674 7966
rect 9702 7993 9730 7999
rect 9702 7967 9703 7993
rect 9729 7967 9730 7993
rect 9534 7938 9562 7943
rect 9198 7657 9282 7658
rect 9198 7631 9255 7657
rect 9281 7631 9282 7657
rect 9198 7630 9282 7631
rect 9142 7266 9170 7271
rect 9086 7265 9170 7266
rect 9086 7239 9143 7265
rect 9169 7239 9170 7265
rect 9086 7238 9170 7239
rect 9142 7233 9170 7238
rect 9030 7154 9058 7159
rect 8918 6930 8946 6935
rect 8918 6929 9002 6930
rect 8918 6903 8919 6929
rect 8945 6903 9002 6929
rect 8918 6902 9002 6903
rect 8918 6897 8946 6902
rect 8974 6818 9002 6902
rect 9030 6929 9058 7126
rect 9030 6903 9031 6929
rect 9057 6903 9058 6929
rect 9030 6897 9058 6903
rect 9198 6818 9226 7630
rect 9254 7625 9282 7630
rect 9366 7937 9562 7938
rect 9366 7911 9535 7937
rect 9561 7911 9562 7937
rect 9366 7910 9562 7911
rect 9310 7602 9338 7607
rect 9254 7321 9282 7327
rect 9254 7295 9255 7321
rect 9281 7295 9282 7321
rect 9254 7266 9282 7295
rect 9254 7233 9282 7238
rect 9254 7154 9282 7159
rect 9310 7154 9338 7574
rect 9366 7265 9394 7910
rect 9534 7905 9562 7910
rect 9702 7882 9730 7967
rect 9702 7849 9730 7854
rect 9758 7770 9786 8806
rect 9814 8441 9842 10038
rect 9870 10122 9898 10127
rect 10318 10094 10346 10318
rect 9870 9617 9898 10094
rect 10262 10066 10346 10094
rect 10542 11074 10570 11079
rect 9870 9591 9871 9617
rect 9897 9591 9898 9617
rect 9870 9585 9898 9591
rect 9926 9730 9954 9735
rect 9926 9561 9954 9702
rect 10206 9730 10234 9735
rect 10206 9683 10234 9702
rect 9926 9535 9927 9561
rect 9953 9535 9954 9561
rect 9926 9529 9954 9535
rect 10150 9561 10178 9567
rect 10150 9535 10151 9561
rect 10177 9535 10178 9561
rect 10038 9506 10066 9511
rect 10038 9505 10122 9506
rect 10038 9479 10039 9505
rect 10065 9479 10122 9505
rect 10038 9478 10122 9479
rect 10038 9473 10066 9478
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9870 9282 9898 9287
rect 9898 9254 10010 9282
rect 9870 9249 9898 9254
rect 9982 9225 10010 9254
rect 9982 9199 9983 9225
rect 10009 9199 10010 9225
rect 9982 9193 10010 9199
rect 10094 9225 10122 9478
rect 10150 9338 10178 9535
rect 10206 9506 10234 9511
rect 10206 9459 10234 9478
rect 10262 9394 10290 10066
rect 10150 9305 10178 9310
rect 10206 9366 10290 9394
rect 10094 9199 10095 9225
rect 10121 9199 10122 9225
rect 10094 9193 10122 9199
rect 9870 9170 9898 9175
rect 9870 9058 9898 9142
rect 10206 9114 10234 9366
rect 9870 9025 9898 9030
rect 10094 9086 10234 9114
rect 10262 9113 10290 9119
rect 10262 9087 10263 9113
rect 10289 9087 10290 9113
rect 10094 8833 10122 9086
rect 10262 8834 10290 9087
rect 10094 8807 10095 8833
rect 10121 8807 10122 8833
rect 10094 8801 10122 8807
rect 10206 8806 10290 8834
rect 10150 8778 10178 8783
rect 10150 8731 10178 8750
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9814 8415 9815 8441
rect 9841 8415 9842 8441
rect 9814 8409 9842 8415
rect 10206 8386 10234 8806
rect 10262 8722 10290 8727
rect 10262 8721 10514 8722
rect 10262 8695 10263 8721
rect 10289 8695 10514 8721
rect 10262 8694 10514 8695
rect 10262 8689 10290 8694
rect 10206 8353 10234 8358
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9814 7770 9842 7775
rect 9366 7239 9367 7265
rect 9393 7239 9394 7265
rect 9366 7233 9394 7239
rect 9478 7769 9842 7770
rect 9478 7743 9815 7769
rect 9841 7743 9842 7769
rect 9478 7742 9842 7743
rect 9478 7265 9506 7742
rect 9814 7737 9842 7742
rect 9926 7770 9954 7775
rect 10374 7770 10402 7775
rect 9478 7239 9479 7265
rect 9505 7239 9506 7265
rect 9478 7233 9506 7239
rect 9646 7658 9674 7663
rect 9646 7265 9674 7630
rect 9926 7657 9954 7742
rect 9926 7631 9927 7657
rect 9953 7631 9954 7657
rect 9870 7601 9898 7607
rect 9870 7575 9871 7601
rect 9897 7575 9898 7601
rect 9870 7266 9898 7575
rect 9646 7239 9647 7265
rect 9673 7239 9674 7265
rect 9646 7233 9674 7239
rect 9814 7238 9898 7266
rect 9926 7602 9954 7631
rect 10150 7769 10402 7770
rect 10150 7743 10375 7769
rect 10401 7743 10402 7769
rect 10150 7742 10402 7743
rect 10150 7657 10178 7742
rect 10374 7737 10402 7742
rect 10430 7713 10458 7719
rect 10430 7687 10431 7713
rect 10457 7687 10458 7713
rect 10150 7631 10151 7657
rect 10177 7631 10178 7657
rect 10150 7625 10178 7631
rect 10318 7658 10346 7663
rect 10318 7611 10346 7630
rect 9926 7265 9954 7574
rect 9926 7239 9927 7265
rect 9953 7239 9954 7265
rect 9254 7153 9338 7154
rect 9254 7127 9255 7153
rect 9281 7127 9338 7153
rect 9254 7126 9338 7127
rect 9702 7154 9730 7159
rect 9254 7121 9282 7126
rect 9702 7107 9730 7126
rect 9758 7153 9786 7159
rect 9758 7127 9759 7153
rect 9785 7127 9786 7153
rect 9254 6986 9282 6991
rect 9254 6939 9282 6958
rect 9478 6986 9506 6991
rect 8974 6790 9226 6818
rect 9478 6873 9506 6958
rect 9478 6847 9479 6873
rect 9505 6847 9506 6873
rect 8862 6762 8890 6767
rect 8862 6715 8890 6734
rect 9198 6538 9226 6543
rect 9198 6491 9226 6510
rect 9478 6537 9506 6847
rect 9478 6511 9479 6537
rect 9505 6511 9506 6537
rect 9478 6505 9506 6511
rect 9534 6538 9562 6543
rect 9534 2169 9562 6510
rect 9758 6538 9786 7127
rect 9814 6930 9842 7238
rect 9926 7233 9954 7239
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9870 6930 9898 6935
rect 9814 6929 9898 6930
rect 9814 6903 9871 6929
rect 9897 6903 9898 6929
rect 9814 6902 9898 6903
rect 9870 6897 9898 6902
rect 10430 6762 10458 7687
rect 10486 7713 10514 8694
rect 10486 7687 10487 7713
rect 10513 7687 10514 7713
rect 10486 7681 10514 7687
rect 10542 7994 10570 11046
rect 10822 10345 10850 11214
rect 10934 11185 10962 11214
rect 10990 11195 11018 11214
rect 10934 11159 10935 11185
rect 10961 11159 10962 11185
rect 10934 11153 10962 11159
rect 11046 11073 11074 12614
rect 11102 12609 11130 12614
rect 11550 12642 11578 12647
rect 11550 12595 11578 12614
rect 11830 12642 11858 13062
rect 11886 13057 11914 13062
rect 12110 13090 12138 13846
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 18830 13537 18858 13543
rect 18830 13511 18831 13537
rect 18857 13511 18858 13537
rect 13174 13481 13202 13487
rect 13174 13455 13175 13481
rect 13201 13455 13202 13481
rect 12558 13425 12586 13431
rect 12558 13399 12559 13425
rect 12585 13399 12586 13425
rect 12334 13090 12362 13095
rect 12110 13089 12334 13090
rect 12110 13063 12111 13089
rect 12137 13063 12334 13089
rect 12110 13062 12334 13063
rect 12110 13057 12138 13062
rect 11942 12754 11970 12759
rect 11942 12697 11970 12726
rect 11942 12671 11943 12697
rect 11969 12671 11970 12697
rect 11942 12665 11970 12671
rect 12278 12754 12306 12759
rect 12334 12754 12362 13062
rect 12558 13090 12586 13399
rect 13174 13426 13202 13455
rect 13174 13393 13202 13398
rect 13230 13481 13258 13487
rect 13230 13455 13231 13481
rect 13257 13455 13258 13481
rect 12558 13057 12586 13062
rect 12726 13145 12754 13151
rect 12726 13119 12727 13145
rect 12753 13119 12754 13145
rect 12726 13090 12754 13119
rect 12726 13057 12754 13062
rect 13118 13089 13146 13095
rect 13118 13063 13119 13089
rect 13145 13063 13146 13089
rect 12278 12753 12362 12754
rect 12278 12727 12279 12753
rect 12305 12727 12362 12753
rect 12278 12726 12362 12727
rect 11830 12609 11858 12614
rect 12110 12642 12138 12647
rect 12110 12595 12138 12614
rect 12222 12306 12250 12311
rect 12278 12306 12306 12726
rect 12670 12697 12698 12703
rect 12670 12671 12671 12697
rect 12697 12671 12698 12697
rect 12670 12473 12698 12671
rect 12670 12447 12671 12473
rect 12697 12447 12698 12473
rect 12670 12441 12698 12447
rect 12838 12642 12866 12647
rect 12614 12362 12642 12367
rect 12726 12362 12754 12367
rect 12614 12315 12642 12334
rect 12670 12361 12754 12362
rect 12670 12335 12727 12361
rect 12753 12335 12754 12361
rect 12670 12334 12754 12335
rect 12222 12305 12306 12306
rect 12222 12279 12223 12305
rect 12249 12279 12306 12305
rect 12222 12278 12306 12279
rect 12054 11634 12082 11639
rect 12054 11587 12082 11606
rect 11942 11578 11970 11583
rect 11718 11550 11942 11578
rect 11718 11522 11746 11550
rect 11942 11531 11970 11550
rect 11606 11521 11746 11522
rect 11606 11495 11719 11521
rect 11745 11495 11746 11521
rect 11606 11494 11746 11495
rect 12222 11522 12250 12278
rect 12278 11522 12306 11527
rect 12222 11521 12362 11522
rect 12222 11495 12279 11521
rect 12305 11495 12362 11521
rect 12222 11494 12362 11495
rect 11158 11270 11354 11298
rect 11158 11241 11186 11270
rect 11158 11215 11159 11241
rect 11185 11215 11186 11241
rect 11158 11209 11186 11215
rect 11326 11242 11354 11270
rect 11494 11242 11522 11247
rect 11326 11241 11522 11242
rect 11326 11215 11495 11241
rect 11521 11215 11522 11241
rect 11326 11214 11522 11215
rect 11494 11209 11522 11214
rect 11270 11185 11298 11191
rect 11270 11159 11271 11185
rect 11297 11159 11298 11185
rect 11270 11130 11298 11159
rect 11606 11185 11634 11494
rect 11718 11489 11746 11494
rect 12278 11489 12306 11494
rect 12110 11298 12138 11303
rect 11606 11159 11607 11185
rect 11633 11159 11634 11185
rect 11606 11153 11634 11159
rect 11942 11185 11970 11191
rect 11942 11159 11943 11185
rect 11969 11159 11970 11185
rect 11438 11130 11466 11135
rect 11270 11097 11298 11102
rect 11326 11129 11466 11130
rect 11326 11103 11439 11129
rect 11465 11103 11466 11129
rect 11326 11102 11466 11103
rect 11046 11047 11047 11073
rect 11073 11047 11074 11073
rect 11046 11018 11074 11047
rect 11326 11018 11354 11102
rect 11438 11097 11466 11102
rect 11550 11130 11578 11135
rect 11046 10985 11074 10990
rect 11270 10990 11354 11018
rect 11270 10626 11298 10990
rect 11326 10906 11354 10911
rect 11494 10906 11522 10911
rect 11326 10905 11494 10906
rect 11326 10879 11327 10905
rect 11353 10879 11494 10905
rect 11326 10878 11494 10879
rect 11326 10873 11354 10878
rect 11494 10873 11522 10878
rect 11550 10905 11578 11102
rect 11550 10879 11551 10905
rect 11577 10879 11578 10905
rect 11550 10873 11578 10879
rect 11942 10906 11970 11159
rect 11942 10873 11970 10878
rect 12054 10849 12082 10855
rect 12054 10823 12055 10849
rect 12081 10823 12082 10849
rect 11494 10794 11522 10799
rect 11270 10598 11466 10626
rect 10822 10319 10823 10345
rect 10849 10319 10850 10345
rect 10654 10289 10682 10295
rect 10654 10263 10655 10289
rect 10681 10263 10682 10289
rect 10654 9730 10682 10263
rect 10710 10066 10738 10071
rect 10710 10019 10738 10038
rect 10822 10010 10850 10319
rect 11158 10346 11186 10351
rect 11158 10299 11186 10318
rect 11326 10289 11354 10295
rect 11326 10263 11327 10289
rect 11353 10263 11354 10289
rect 10822 9977 10850 9982
rect 11102 10122 11130 10127
rect 10654 9697 10682 9702
rect 10934 9618 10962 9623
rect 10934 9617 11018 9618
rect 10934 9591 10935 9617
rect 10961 9591 11018 9617
rect 10934 9590 11018 9591
rect 10934 9585 10962 9590
rect 10654 9506 10682 9511
rect 10598 9281 10626 9287
rect 10598 9255 10599 9281
rect 10625 9255 10626 9281
rect 10598 9170 10626 9255
rect 10598 9137 10626 9142
rect 10654 8777 10682 9478
rect 10654 8751 10655 8777
rect 10681 8751 10682 8777
rect 10654 8745 10682 8751
rect 10766 9225 10794 9231
rect 10766 9199 10767 9225
rect 10793 9199 10794 9225
rect 10766 8778 10794 9199
rect 10934 9226 10962 9231
rect 10934 9179 10962 9198
rect 10822 8778 10850 8783
rect 10766 8750 10822 8778
rect 10822 8731 10850 8750
rect 10990 8442 11018 9590
rect 11102 9225 11130 10094
rect 11270 9562 11298 9567
rect 11158 9561 11298 9562
rect 11158 9535 11271 9561
rect 11297 9535 11298 9561
rect 11158 9534 11298 9535
rect 11158 9337 11186 9534
rect 11270 9529 11298 9534
rect 11326 9394 11354 10263
rect 11326 9361 11354 9366
rect 11158 9311 11159 9337
rect 11185 9311 11186 9337
rect 11158 9305 11186 9311
rect 11382 9338 11410 9343
rect 11382 9291 11410 9310
rect 11214 9282 11242 9287
rect 11214 9235 11242 9254
rect 11102 9199 11103 9225
rect 11129 9199 11130 9225
rect 11102 9193 11130 9199
rect 11438 9170 11466 10598
rect 11494 10178 11522 10766
rect 11494 10145 11522 10150
rect 11606 10793 11634 10799
rect 11606 10767 11607 10793
rect 11633 10767 11634 10793
rect 11606 10094 11634 10767
rect 11830 10794 11858 10799
rect 11942 10794 11970 10799
rect 11830 10793 11970 10794
rect 11830 10767 11831 10793
rect 11857 10767 11943 10793
rect 11969 10767 11970 10793
rect 11830 10766 11970 10767
rect 11830 10761 11858 10766
rect 11438 9137 11466 9142
rect 11494 10066 11634 10094
rect 11942 10066 11970 10766
rect 12054 10794 12082 10823
rect 12110 10849 12138 11270
rect 12278 11130 12306 11135
rect 12110 10823 12111 10849
rect 12137 10823 12138 10849
rect 12110 10817 12138 10823
rect 12166 11129 12306 11130
rect 12166 11103 12279 11129
rect 12305 11103 12306 11129
rect 12166 11102 12306 11103
rect 12054 10761 12082 10766
rect 12110 10738 12138 10743
rect 12166 10738 12194 11102
rect 12278 11097 12306 11102
rect 12278 10906 12306 10911
rect 12334 10906 12362 11494
rect 12670 11242 12698 12334
rect 12726 12329 12754 12334
rect 12306 10878 12362 10906
rect 12614 11214 12698 11242
rect 12278 10873 12306 10878
rect 12334 10794 12362 10799
rect 12334 10747 12362 10766
rect 12110 10737 12194 10738
rect 12110 10711 12111 10737
rect 12137 10711 12194 10737
rect 12110 10710 12194 10711
rect 12110 10705 12138 10710
rect 11494 9226 11522 10066
rect 11942 10033 11970 10038
rect 12558 10066 12586 10071
rect 12558 10019 12586 10038
rect 12614 10010 12642 11214
rect 12782 10962 12810 10967
rect 12782 10905 12810 10934
rect 12782 10879 12783 10905
rect 12809 10879 12810 10905
rect 12782 10873 12810 10879
rect 12838 10850 12866 12614
rect 13062 12474 13090 12479
rect 13062 12427 13090 12446
rect 13118 12473 13146 13063
rect 13230 13090 13258 13455
rect 13230 13057 13258 13062
rect 13342 13425 13370 13431
rect 13342 13399 13343 13425
rect 13369 13399 13370 13425
rect 13118 12447 13119 12473
rect 13145 12447 13146 12473
rect 13118 12441 13146 12447
rect 12950 12418 12978 12423
rect 12950 12361 12978 12390
rect 12950 12335 12951 12361
rect 12977 12335 12978 12361
rect 12950 12329 12978 12335
rect 13174 12362 13202 12367
rect 13174 12315 13202 12334
rect 13342 12361 13370 13399
rect 18830 13258 18858 13511
rect 18830 13225 18858 13230
rect 14518 13202 14546 13207
rect 14518 13155 14546 13174
rect 14406 13146 14434 13151
rect 14182 13118 14406 13146
rect 13958 13090 13986 13095
rect 14182 13090 14210 13118
rect 14406 13099 14434 13118
rect 18830 13146 18858 13151
rect 18830 13099 18858 13118
rect 13986 13089 14210 13090
rect 13986 13063 14183 13089
rect 14209 13063 14210 13089
rect 13986 13062 14210 13063
rect 13734 12809 13762 12815
rect 13734 12783 13735 12809
rect 13761 12783 13762 12809
rect 13734 12754 13762 12783
rect 13566 12726 13734 12754
rect 13510 12642 13538 12647
rect 13342 12335 13343 12361
rect 13369 12335 13370 12361
rect 13342 12329 13370 12335
rect 13454 12474 13482 12479
rect 13342 11241 13370 11247
rect 13342 11215 13343 11241
rect 13369 11215 13370 11241
rect 13342 10962 13370 11215
rect 13454 11186 13482 12446
rect 13510 12417 13538 12614
rect 13566 12473 13594 12726
rect 13734 12721 13762 12726
rect 13958 12753 13986 13062
rect 14182 13057 14210 13062
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 13958 12727 13959 12753
rect 13985 12727 13986 12753
rect 13958 12721 13986 12727
rect 18830 12754 18858 12759
rect 18830 12707 18858 12726
rect 14070 12642 14098 12647
rect 14070 12595 14098 12614
rect 18942 12642 18970 13903
rect 19950 13873 19978 13879
rect 19950 13847 19951 13873
rect 19977 13847 19978 13873
rect 19950 13482 19978 13847
rect 19950 13449 19978 13454
rect 20006 13593 20034 13599
rect 20006 13567 20007 13593
rect 20033 13567 20034 13593
rect 20006 13146 20034 13567
rect 20006 13113 20034 13118
rect 19950 13089 19978 13095
rect 19950 13063 19951 13089
rect 19977 13063 19978 13089
rect 19950 12810 19978 13063
rect 19950 12777 19978 12782
rect 20006 12809 20034 12815
rect 20006 12783 20007 12809
rect 20033 12783 20034 12809
rect 18942 12609 18970 12614
rect 13566 12447 13567 12473
rect 13593 12447 13594 12473
rect 13566 12441 13594 12447
rect 20006 12474 20034 12783
rect 20006 12441 20034 12446
rect 13510 12391 13511 12417
rect 13537 12391 13538 12417
rect 13510 12385 13538 12391
rect 13678 12418 13706 12423
rect 13678 12371 13706 12390
rect 18942 12361 18970 12367
rect 18942 12335 18943 12361
rect 18969 12335 18970 12361
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 18830 11970 18858 11975
rect 18774 11969 18858 11970
rect 18774 11943 18831 11969
rect 18857 11943 18858 11969
rect 18774 11942 18858 11943
rect 18774 11578 18802 11942
rect 18830 11937 18858 11942
rect 18942 11634 18970 12335
rect 20006 12249 20034 12255
rect 20006 12223 20007 12249
rect 20033 12223 20034 12249
rect 20006 12138 20034 12223
rect 20006 12105 20034 12110
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 20006 11802 20034 11999
rect 20006 11769 20034 11774
rect 18942 11601 18970 11606
rect 18774 11545 18802 11550
rect 18830 11577 18858 11583
rect 18830 11551 18831 11577
rect 18857 11551 18858 11577
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 18830 11354 18858 11551
rect 20006 11466 20034 11471
rect 20006 11419 20034 11438
rect 17598 11349 17730 11354
rect 18774 11326 18858 11354
rect 13958 11242 13986 11247
rect 13342 10929 13370 10934
rect 13398 11185 13482 11186
rect 13398 11159 13455 11185
rect 13481 11159 13482 11185
rect 13398 11158 13482 11159
rect 13062 10906 13090 10911
rect 12838 10849 12922 10850
rect 12838 10823 12839 10849
rect 12865 10823 12922 10849
rect 12838 10822 12922 10823
rect 12838 10817 12866 10822
rect 12670 10794 12698 10799
rect 12670 10747 12698 10766
rect 12614 9977 12642 9982
rect 12670 10065 12698 10071
rect 12670 10039 12671 10065
rect 12697 10039 12698 10065
rect 12670 9786 12698 10039
rect 12670 9753 12698 9758
rect 12726 10009 12754 10015
rect 12726 9983 12727 10009
rect 12753 9983 12754 10009
rect 12334 9673 12362 9679
rect 12334 9647 12335 9673
rect 12361 9647 12362 9673
rect 11886 9394 11914 9399
rect 11438 8778 11466 8783
rect 11494 8778 11522 9198
rect 11550 9225 11578 9231
rect 11550 9199 11551 9225
rect 11577 9199 11578 9225
rect 11550 8946 11578 9199
rect 11550 8833 11578 8918
rect 11886 9225 11914 9366
rect 11886 9199 11887 9225
rect 11913 9199 11914 9225
rect 11886 8945 11914 9199
rect 11886 8919 11887 8945
rect 11913 8919 11914 8945
rect 11886 8913 11914 8919
rect 11998 9225 12026 9231
rect 11998 9199 11999 9225
rect 12025 9199 12026 9225
rect 11942 8890 11970 8895
rect 11942 8843 11970 8862
rect 11550 8807 11551 8833
rect 11577 8807 11578 8833
rect 11550 8801 11578 8807
rect 11438 8777 11522 8778
rect 11438 8751 11439 8777
rect 11465 8751 11522 8777
rect 11438 8750 11522 8751
rect 11942 8778 11970 8783
rect 11998 8778 12026 9199
rect 12278 9169 12306 9175
rect 12278 9143 12279 9169
rect 12305 9143 12306 9169
rect 12278 9002 12306 9143
rect 12278 8969 12306 8974
rect 12222 8946 12250 8951
rect 12222 8899 12250 8918
rect 12334 8890 12362 9647
rect 12670 9506 12698 9511
rect 12726 9506 12754 9983
rect 12838 9898 12866 9903
rect 12670 9505 12754 9506
rect 12670 9479 12671 9505
rect 12697 9479 12754 9505
rect 12670 9478 12754 9479
rect 12782 9786 12810 9791
rect 12614 9281 12642 9287
rect 12614 9255 12615 9281
rect 12641 9255 12642 9281
rect 12334 8857 12362 8862
rect 12558 8946 12586 8951
rect 12614 8946 12642 9255
rect 12586 8918 12642 8946
rect 12558 8833 12586 8918
rect 12558 8807 12559 8833
rect 12585 8807 12586 8833
rect 12558 8801 12586 8807
rect 12110 8778 12138 8783
rect 11970 8750 12026 8778
rect 12054 8777 12138 8778
rect 12054 8751 12111 8777
rect 12137 8751 12138 8777
rect 12054 8750 12138 8751
rect 11438 8745 11466 8750
rect 10990 8409 11018 8414
rect 11774 8554 11802 8559
rect 10878 8386 10906 8391
rect 10822 8050 10850 8055
rect 10542 7658 10570 7966
rect 10710 8022 10822 8050
rect 10654 7937 10682 7943
rect 10654 7911 10655 7937
rect 10681 7911 10682 7937
rect 10654 7770 10682 7911
rect 10654 7737 10682 7742
rect 10542 7625 10570 7630
rect 10710 7657 10738 8022
rect 10822 8003 10850 8022
rect 10878 7713 10906 8358
rect 11774 8386 11802 8526
rect 11550 8049 11578 8055
rect 11550 8023 11551 8049
rect 11577 8023 11578 8049
rect 11550 7994 11578 8023
rect 11774 8049 11802 8358
rect 11774 8023 11775 8049
rect 11801 8023 11802 8049
rect 11774 8017 11802 8023
rect 11886 8050 11914 8055
rect 11550 7961 11578 7966
rect 11830 7938 11858 7943
rect 11830 7891 11858 7910
rect 11830 7770 11858 7775
rect 11886 7770 11914 8022
rect 11942 7994 11970 8750
rect 12054 8106 12082 8750
rect 12110 8745 12138 8750
rect 12390 8722 12418 8727
rect 12390 8675 12418 8694
rect 12614 8721 12642 8727
rect 12614 8695 12615 8721
rect 12641 8695 12642 8721
rect 12166 8442 12194 8447
rect 12110 8386 12138 8391
rect 12166 8386 12194 8414
rect 12110 8385 12194 8386
rect 12110 8359 12111 8385
rect 12137 8359 12194 8385
rect 12110 8358 12194 8359
rect 12110 8353 12138 8358
rect 12110 8106 12138 8111
rect 12054 8105 12138 8106
rect 12054 8079 12111 8105
rect 12137 8079 12138 8105
rect 12054 8078 12138 8079
rect 12054 7994 12082 7999
rect 11942 7993 12082 7994
rect 11942 7967 12055 7993
rect 12081 7967 12082 7993
rect 11942 7966 12082 7967
rect 12054 7961 12082 7966
rect 12110 7882 12138 8078
rect 11830 7769 11914 7770
rect 11830 7743 11831 7769
rect 11857 7743 11914 7769
rect 11830 7742 11914 7743
rect 11998 7854 12138 7882
rect 11998 7769 12026 7854
rect 11998 7743 11999 7769
rect 12025 7743 12026 7769
rect 11830 7737 11858 7742
rect 11998 7737 12026 7743
rect 10878 7687 10879 7713
rect 10905 7687 10906 7713
rect 10878 7681 10906 7687
rect 11046 7713 11074 7719
rect 11046 7687 11047 7713
rect 11073 7687 11074 7713
rect 10710 7631 10711 7657
rect 10737 7631 10738 7657
rect 10710 7625 10738 7631
rect 11046 7321 11074 7687
rect 11046 7295 11047 7321
rect 11073 7295 11074 7321
rect 11046 7289 11074 7295
rect 12110 7321 12138 7854
rect 12166 7602 12194 8358
rect 12614 8050 12642 8695
rect 12670 8722 12698 9478
rect 12726 9225 12754 9231
rect 12726 9199 12727 9225
rect 12753 9199 12754 9225
rect 12726 8890 12754 9199
rect 12726 8857 12754 8862
rect 12726 8778 12754 8783
rect 12782 8778 12810 9758
rect 12838 9505 12866 9870
rect 12838 9479 12839 9505
rect 12865 9479 12866 9505
rect 12838 9282 12866 9479
rect 12838 9249 12866 9254
rect 12894 9002 12922 10822
rect 13062 10794 13090 10878
rect 13398 10850 13426 11158
rect 13454 11153 13482 11158
rect 13678 11241 13986 11242
rect 13678 11215 13959 11241
rect 13985 11215 13986 11241
rect 13678 11214 13986 11215
rect 13678 11185 13706 11214
rect 13958 11209 13986 11214
rect 13678 11159 13679 11185
rect 13705 11159 13706 11185
rect 13678 11153 13706 11159
rect 14630 11185 14658 11191
rect 14630 11159 14631 11185
rect 14657 11159 14658 11185
rect 13790 11130 13818 11135
rect 13790 11083 13818 11102
rect 14014 11129 14042 11135
rect 14014 11103 14015 11129
rect 14041 11103 14042 11129
rect 13286 10822 13426 10850
rect 13622 11073 13650 11079
rect 13622 11047 13623 11073
rect 13649 11047 13650 11073
rect 13622 10849 13650 11047
rect 14014 11074 14042 11103
rect 14014 11041 14042 11046
rect 14630 11074 14658 11159
rect 14966 11185 14994 11191
rect 14966 11159 14967 11185
rect 14993 11159 14994 11185
rect 13622 10823 13623 10849
rect 13649 10823 13650 10849
rect 13230 10794 13258 10799
rect 13062 10793 13258 10794
rect 13062 10767 13063 10793
rect 13089 10767 13231 10793
rect 13257 10767 13258 10793
rect 13062 10766 13258 10767
rect 13062 10761 13090 10766
rect 13230 10761 13258 10766
rect 13006 10010 13034 10015
rect 12950 9953 12978 9959
rect 12950 9927 12951 9953
rect 12977 9927 12978 9953
rect 12950 9226 12978 9927
rect 13006 9729 13034 9982
rect 13286 9898 13314 10822
rect 13622 10817 13650 10823
rect 14630 10738 14658 11046
rect 14742 11073 14770 11079
rect 14742 11047 14743 11073
rect 14769 11047 14770 11073
rect 14686 10738 14714 10743
rect 14630 10737 14714 10738
rect 14630 10711 14687 10737
rect 14713 10711 14714 10737
rect 14630 10710 14714 10711
rect 14686 10705 14714 10710
rect 14742 10402 14770 11047
rect 14966 11074 14994 11159
rect 14966 11041 14994 11046
rect 15078 11073 15106 11079
rect 15078 11047 15079 11073
rect 15105 11047 15106 11073
rect 15078 10794 15106 11047
rect 18774 11074 18802 11326
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 18774 11041 18802 11046
rect 18830 11185 18858 11191
rect 18830 11159 18831 11185
rect 18857 11159 18858 11185
rect 18830 10962 18858 11159
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 18830 10929 18858 10934
rect 15078 10761 15106 10766
rect 18830 10794 18858 10799
rect 18830 10747 18858 10766
rect 20006 10794 20034 10799
rect 20006 10737 20034 10766
rect 20006 10711 20007 10737
rect 20033 10711 20034 10737
rect 20006 10705 20034 10711
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 20006 10458 20034 10463
rect 20006 10411 20034 10430
rect 14742 10369 14770 10374
rect 18830 10402 18858 10407
rect 18830 10355 18858 10374
rect 13286 9865 13314 9870
rect 17598 9814 17730 9819
rect 13286 9786 13314 9791
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 13314 9758 13370 9786
rect 17598 9781 17730 9786
rect 13286 9753 13314 9758
rect 13006 9703 13007 9729
rect 13033 9703 13034 9729
rect 13006 9697 13034 9703
rect 13118 9617 13146 9623
rect 13118 9591 13119 9617
rect 13145 9591 13146 9617
rect 13062 9226 13090 9245
rect 12950 9198 13062 9226
rect 12894 8969 12922 8974
rect 12726 8777 12810 8778
rect 12726 8751 12727 8777
rect 12753 8751 12810 8777
rect 12726 8750 12810 8751
rect 12894 8834 12922 8839
rect 13006 8834 13034 9198
rect 13062 9193 13090 9198
rect 12894 8833 13034 8834
rect 12894 8807 12895 8833
rect 12921 8807 13034 8833
rect 12894 8806 13034 8807
rect 12726 8745 12754 8750
rect 12670 8689 12698 8694
rect 12670 8442 12698 8447
rect 12670 8395 12698 8414
rect 12894 8442 12922 8806
rect 12894 8409 12922 8414
rect 13006 8722 13034 8727
rect 13006 8441 13034 8694
rect 13006 8415 13007 8441
rect 13033 8415 13034 8441
rect 13006 8409 13034 8415
rect 13118 8386 13146 9591
rect 13286 9617 13314 9623
rect 13286 9591 13287 9617
rect 13313 9591 13314 9617
rect 13230 9226 13258 9231
rect 13230 9179 13258 9198
rect 13118 8339 13146 8358
rect 13174 9002 13202 9007
rect 12614 8017 12642 8022
rect 12614 7938 12642 7943
rect 12614 7769 12642 7910
rect 12614 7743 12615 7769
rect 12641 7743 12642 7769
rect 12614 7737 12642 7743
rect 12726 7882 12754 7887
rect 12726 7769 12754 7854
rect 12726 7743 12727 7769
rect 12753 7743 12754 7769
rect 12726 7737 12754 7743
rect 13006 7714 13034 7719
rect 12950 7713 13034 7714
rect 12950 7687 13007 7713
rect 13033 7687 13034 7713
rect 12950 7686 13034 7687
rect 12950 7657 12978 7686
rect 13006 7681 13034 7686
rect 13118 7713 13146 7719
rect 13118 7687 13119 7713
rect 13145 7687 13146 7713
rect 12950 7631 12951 7657
rect 12977 7631 12978 7657
rect 12950 7625 12978 7631
rect 12222 7602 12250 7607
rect 12166 7601 12250 7602
rect 12166 7575 12223 7601
rect 12249 7575 12250 7601
rect 12166 7574 12250 7575
rect 12110 7295 12111 7321
rect 12137 7295 12138 7321
rect 12110 7289 12138 7295
rect 10654 7265 10682 7271
rect 10654 7239 10655 7265
rect 10681 7239 10682 7265
rect 10654 6986 10682 7239
rect 12222 7266 12250 7574
rect 12670 7601 12698 7607
rect 12670 7575 12671 7601
rect 12697 7575 12698 7601
rect 12670 7321 12698 7575
rect 12670 7295 12671 7321
rect 12697 7295 12698 7321
rect 12670 7289 12698 7295
rect 13118 7322 13146 7687
rect 13174 7713 13202 8974
rect 13230 8778 13258 8783
rect 13230 8731 13258 8750
rect 13230 8386 13258 8391
rect 13286 8386 13314 9591
rect 13342 9617 13370 9758
rect 20006 9673 20034 9679
rect 20006 9647 20007 9673
rect 20033 9647 20034 9673
rect 13342 9591 13343 9617
rect 13369 9591 13370 9617
rect 13342 8553 13370 9591
rect 14238 9618 14266 9623
rect 14238 9571 14266 9590
rect 14686 9618 14714 9623
rect 13398 9505 13426 9511
rect 13398 9479 13399 9505
rect 13425 9479 13426 9505
rect 13398 9226 13426 9479
rect 13454 9506 13482 9511
rect 14182 9506 14210 9511
rect 13454 9505 14210 9506
rect 13454 9479 13455 9505
rect 13481 9479 14183 9505
rect 14209 9479 14210 9505
rect 13454 9478 14210 9479
rect 13454 9473 13482 9478
rect 14182 9473 14210 9478
rect 13622 9226 13650 9231
rect 13398 9225 13650 9226
rect 13398 9199 13623 9225
rect 13649 9199 13650 9225
rect 13398 9198 13650 9199
rect 13622 9193 13650 9198
rect 14686 9169 14714 9590
rect 18830 9618 18858 9623
rect 18830 9571 18858 9590
rect 20006 9450 20034 9647
rect 20006 9417 20034 9422
rect 14686 9143 14687 9169
rect 14713 9143 14714 9169
rect 14686 9137 14714 9143
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 14294 8890 14322 8895
rect 14294 8843 14322 8862
rect 14630 8890 14658 8895
rect 14630 8843 14658 8862
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 13342 8527 13343 8553
rect 13369 8527 13370 8553
rect 13342 8521 13370 8527
rect 13398 8778 13426 8783
rect 13398 8553 13426 8750
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 13398 8527 13399 8553
rect 13425 8527 13426 8553
rect 13398 8521 13426 8527
rect 13454 8722 13482 8727
rect 13454 8553 13482 8694
rect 14574 8722 14602 8727
rect 14574 8675 14602 8694
rect 13454 8527 13455 8553
rect 13481 8527 13482 8553
rect 13454 8521 13482 8527
rect 13230 8385 13314 8386
rect 13230 8359 13231 8385
rect 13257 8359 13314 8385
rect 13230 8358 13314 8359
rect 13230 7882 13258 8358
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 13230 7849 13258 7854
rect 13174 7687 13175 7713
rect 13201 7687 13202 7713
rect 13174 7681 13202 7687
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 12278 7266 12306 7271
rect 12222 7265 12306 7266
rect 12222 7239 12279 7265
rect 12305 7239 12306 7265
rect 12222 7238 12306 7239
rect 10654 6953 10682 6958
rect 11158 6986 11186 6991
rect 11158 6939 11186 6958
rect 12110 6986 12138 6991
rect 12278 6986 12306 7238
rect 12138 6958 12306 6986
rect 12110 6939 12138 6958
rect 10934 6817 10962 6823
rect 10934 6791 10935 6817
rect 10961 6791 10962 6817
rect 10542 6762 10570 6767
rect 10430 6734 10542 6762
rect 9758 6505 9786 6510
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9534 2143 9535 2169
rect 9561 2143 9562 2169
rect 9534 2137 9562 2143
rect 9422 2058 9450 2063
rect 9310 1834 9338 1839
rect 8806 1751 8807 1777
rect 8833 1751 8834 1777
rect 8806 1745 8834 1751
rect 9086 1833 9338 1834
rect 9086 1807 9311 1833
rect 9337 1807 9338 1833
rect 9086 1806 9338 1807
rect 9086 400 9114 1806
rect 9310 1801 9338 1806
rect 9422 400 9450 2030
rect 10038 2058 10066 2063
rect 10038 2011 10066 2030
rect 10430 1834 10458 1839
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10430 400 10458 1806
rect 10542 1777 10570 6734
rect 10934 6762 10962 6791
rect 10934 6729 10962 6734
rect 13118 4214 13146 7294
rect 13734 7322 13762 7327
rect 13734 7275 13762 7294
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 13118 4186 13258 4214
rect 13230 2169 13258 4186
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 13230 2143 13231 2169
rect 13257 2143 13258 2169
rect 13230 2137 13258 2143
rect 13118 2058 13146 2063
rect 11046 1834 11074 1839
rect 11046 1787 11074 1806
rect 10542 1751 10543 1777
rect 10569 1751 10570 1777
rect 10542 1745 10570 1751
rect 13118 400 13146 2030
rect 13734 2058 13762 2063
rect 13734 2011 13762 2030
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 9072 0 9128 400
rect 9408 0 9464 400
rect 10416 0 10472 400
rect 13104 0 13160 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 9758 19278 9786 19306
rect 10374 19278 10402 19306
rect 9086 18326 9114 18354
rect 9590 18353 9618 18354
rect 9590 18327 9591 18353
rect 9591 18327 9617 18353
rect 9617 18327 9618 18353
rect 9590 18326 9618 18327
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 8470 13537 8498 13538
rect 8470 13511 8471 13537
rect 8471 13511 8497 13537
rect 8497 13511 8498 13537
rect 8470 13510 8498 13511
rect 2086 13454 2114 13482
rect 966 12446 994 12474
rect 966 12249 994 12250
rect 966 12223 967 12249
rect 967 12223 993 12249
rect 993 12223 994 12249
rect 966 12222 994 12223
rect 966 11465 994 11466
rect 966 11439 967 11465
rect 967 11439 993 11465
rect 993 11439 994 11465
rect 966 11438 994 11439
rect 7518 13398 7546 13426
rect 7910 13398 7938 13426
rect 2142 13062 2170 13090
rect 5838 13089 5866 13090
rect 5838 13063 5839 13089
rect 5839 13063 5865 13089
rect 5865 13063 5866 13089
rect 5838 13062 5866 13063
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 5838 12670 5866 12698
rect 6902 12558 6930 12586
rect 2142 12361 2170 12362
rect 2142 12335 2143 12361
rect 2143 12335 2169 12361
rect 2169 12335 2170 12361
rect 2142 12334 2170 12335
rect 6006 12334 6034 12362
rect 7070 12305 7098 12306
rect 7070 12279 7071 12305
rect 7071 12279 7097 12305
rect 7097 12279 7098 12305
rect 7070 12278 7098 12279
rect 7182 12222 7210 12250
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 2142 11577 2170 11578
rect 2142 11551 2143 11577
rect 2143 11551 2169 11577
rect 2169 11551 2170 11577
rect 2142 11550 2170 11551
rect 6174 11550 6202 11578
rect 5726 11521 5754 11522
rect 5726 11495 5727 11521
rect 5727 11495 5753 11521
rect 5753 11495 5754 11521
rect 5726 11494 5754 11495
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 5726 11102 5754 11130
rect 7182 11577 7210 11578
rect 7182 11551 7183 11577
rect 7183 11551 7209 11577
rect 7209 11551 7210 11577
rect 7182 11550 7210 11551
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 11774 19110 11802 19138
rect 8638 13145 8666 13146
rect 8638 13119 8639 13145
rect 8639 13119 8665 13145
rect 8665 13119 8666 13145
rect 8638 13118 8666 13119
rect 8246 13062 8274 13090
rect 6790 11521 6818 11522
rect 6790 11495 6791 11521
rect 6791 11495 6817 11521
rect 6817 11495 6818 11521
rect 6790 11494 6818 11495
rect 7350 12670 7378 12698
rect 7518 12446 7546 12474
rect 7406 12222 7434 12250
rect 7574 12110 7602 12138
rect 7686 12558 7714 12586
rect 7798 12417 7826 12418
rect 7798 12391 7799 12417
rect 7799 12391 7825 12417
rect 7825 12391 7826 12417
rect 7798 12390 7826 12391
rect 7910 12361 7938 12362
rect 7910 12335 7911 12361
rect 7911 12335 7937 12361
rect 7937 12335 7938 12361
rect 7910 12334 7938 12335
rect 7742 12278 7770 12306
rect 7910 12110 7938 12138
rect 8134 12222 8162 12250
rect 7518 11550 7546 11578
rect 7574 11521 7602 11522
rect 7574 11495 7575 11521
rect 7575 11495 7601 11521
rect 7601 11495 7602 11521
rect 7574 11494 7602 11495
rect 7686 11326 7714 11354
rect 7910 11270 7938 11298
rect 6510 10849 6538 10850
rect 6510 10823 6511 10849
rect 6511 10823 6537 10849
rect 6537 10823 6538 10849
rect 6510 10822 6538 10823
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 7350 11129 7378 11130
rect 7350 11103 7351 11129
rect 7351 11103 7377 11129
rect 7377 11103 7378 11129
rect 7350 11102 7378 11103
rect 8694 12390 8722 12418
rect 8918 13089 8946 13090
rect 8918 13063 8919 13089
rect 8919 13063 8945 13089
rect 8945 13063 8946 13089
rect 8918 13062 8946 13063
rect 9254 13145 9282 13146
rect 9254 13119 9255 13145
rect 9255 13119 9281 13145
rect 9281 13119 9282 13145
rect 9254 13118 9282 13119
rect 9422 13145 9450 13146
rect 9422 13119 9423 13145
rect 9423 13119 9449 13145
rect 9449 13119 9450 13145
rect 9422 13118 9450 13119
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 11326 14238 11354 14266
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 9926 13510 9954 13538
rect 10094 13425 10122 13426
rect 10094 13399 10095 13425
rect 10095 13399 10121 13425
rect 10121 13399 10122 13425
rect 10094 13398 10122 13399
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9814 13201 9842 13202
rect 9814 13175 9815 13201
rect 9815 13175 9841 13201
rect 9841 13175 9842 13201
rect 9814 13174 9842 13175
rect 10486 13398 10514 13426
rect 9702 13118 9730 13146
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9142 12390 9170 12418
rect 8750 12334 8778 12362
rect 8974 11662 9002 11690
rect 8806 11297 8834 11298
rect 8806 11271 8807 11297
rect 8807 11271 8833 11297
rect 8833 11271 8834 11297
rect 8806 11270 8834 11271
rect 7910 10849 7938 10850
rect 7910 10823 7911 10849
rect 7911 10823 7937 10849
rect 7937 10823 7938 10849
rect 7910 10822 7938 10823
rect 7574 10766 7602 10794
rect 7966 10793 7994 10794
rect 7966 10767 7967 10793
rect 7967 10767 7993 10793
rect 7993 10767 7994 10793
rect 7966 10766 7994 10767
rect 2142 10009 2170 10010
rect 2142 9983 2143 10009
rect 2143 9983 2169 10009
rect 2169 9983 2170 10009
rect 2142 9982 2170 9983
rect 5502 9982 5530 10010
rect 2086 9926 2114 9954
rect 966 9897 994 9898
rect 966 9871 967 9897
rect 967 9871 993 9897
rect 993 9871 994 9897
rect 966 9870 994 9871
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 5502 9814 5530 9842
rect 2342 9786 2370 9787
rect 6286 9561 6314 9562
rect 6286 9535 6287 9561
rect 6287 9535 6313 9561
rect 6313 9535 6314 9561
rect 6286 9534 6314 9535
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 2142 8833 2170 8834
rect 2142 8807 2143 8833
rect 2143 8807 2169 8833
rect 2169 8807 2170 8833
rect 2142 8806 2170 8807
rect 7182 9814 7210 9842
rect 7126 9561 7154 9562
rect 7126 9535 7127 9561
rect 7127 9535 7153 9561
rect 7153 9535 7154 9561
rect 7126 9534 7154 9535
rect 7238 9561 7266 9562
rect 7238 9535 7239 9561
rect 7239 9535 7265 9561
rect 7265 9535 7266 9561
rect 7238 9534 7266 9535
rect 7462 9702 7490 9730
rect 7070 9086 7098 9114
rect 7350 9086 7378 9114
rect 7406 8806 7434 8834
rect 7238 8721 7266 8722
rect 7238 8695 7239 8721
rect 7239 8695 7265 8721
rect 7265 8695 7266 8721
rect 7238 8694 7266 8695
rect 6958 8526 6986 8554
rect 6342 8497 6370 8498
rect 6342 8471 6343 8497
rect 6343 8471 6369 8497
rect 6369 8471 6370 8497
rect 6342 8470 6370 8471
rect 966 8414 994 8442
rect 6006 8441 6034 8442
rect 6006 8415 6007 8441
rect 6007 8415 6033 8441
rect 6033 8415 6034 8441
rect 6006 8414 6034 8415
rect 6790 8414 6818 8442
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 7406 8470 7434 8498
rect 7910 9646 7938 9674
rect 7742 9561 7770 9562
rect 7742 9535 7743 9561
rect 7743 9535 7769 9561
rect 7769 9535 7770 9561
rect 7742 9534 7770 9535
rect 8078 9478 8106 9506
rect 7462 9198 7490 9226
rect 7742 9086 7770 9114
rect 7854 8833 7882 8834
rect 7854 8807 7855 8833
rect 7855 8807 7881 8833
rect 7881 8807 7882 8833
rect 7854 8806 7882 8807
rect 7910 8750 7938 8778
rect 7854 8694 7882 8722
rect 7518 8526 7546 8554
rect 7574 8078 7602 8106
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 7966 8526 7994 8554
rect 7798 8358 7826 8386
rect 8358 9646 8386 9674
rect 8526 9617 8554 9618
rect 8526 9591 8527 9617
rect 8527 9591 8553 9617
rect 8553 9591 8554 9617
rect 8526 9590 8554 9591
rect 8694 11073 8722 11074
rect 8694 11047 8695 11073
rect 8695 11047 8721 11073
rect 8721 11047 8722 11073
rect 8694 11046 8722 11047
rect 8862 10934 8890 10962
rect 9086 11606 9114 11634
rect 9366 11633 9394 11634
rect 9366 11607 9367 11633
rect 9367 11607 9393 11633
rect 9393 11607 9394 11633
rect 9366 11606 9394 11607
rect 9422 11577 9450 11578
rect 9422 11551 9423 11577
rect 9423 11551 9449 11577
rect 9449 11551 9450 11577
rect 9422 11550 9450 11551
rect 9086 11129 9114 11130
rect 9086 11103 9087 11129
rect 9087 11103 9113 11129
rect 9113 11103 9114 11129
rect 9086 11102 9114 11103
rect 9030 11046 9058 11074
rect 9702 12334 9730 12362
rect 9646 11689 9674 11690
rect 9646 11663 9647 11689
rect 9647 11663 9673 11689
rect 9673 11663 9674 11689
rect 9646 11662 9674 11663
rect 9590 11633 9618 11634
rect 9590 11607 9591 11633
rect 9591 11607 9617 11633
rect 9617 11607 9618 11633
rect 9590 11606 9618 11607
rect 9534 11326 9562 11354
rect 9590 11073 9618 11074
rect 9590 11047 9591 11073
rect 9591 11047 9617 11073
rect 9617 11047 9618 11073
rect 9590 11046 9618 11047
rect 8694 10793 8722 10794
rect 8694 10767 8695 10793
rect 8695 10767 8721 10793
rect 8721 10767 8722 10793
rect 8694 10766 8722 10767
rect 8974 10009 9002 10010
rect 8974 9983 8975 10009
rect 8975 9983 9001 10009
rect 9001 9983 9002 10009
rect 8974 9982 9002 9983
rect 9534 10094 9562 10122
rect 9366 10009 9394 10010
rect 9366 9983 9367 10009
rect 9367 9983 9393 10009
rect 9393 9983 9394 10009
rect 9366 9982 9394 9983
rect 9198 9953 9226 9954
rect 9198 9927 9199 9953
rect 9199 9927 9225 9953
rect 9225 9927 9226 9953
rect 9198 9926 9226 9927
rect 8806 9758 8834 9786
rect 8582 9534 8610 9562
rect 8414 9281 8442 9282
rect 8414 9255 8415 9281
rect 8415 9255 8441 9281
rect 8441 9255 8442 9281
rect 8414 9254 8442 9255
rect 8246 9225 8274 9226
rect 8246 9199 8247 9225
rect 8247 9199 8273 9225
rect 8273 9199 8274 9225
rect 8246 9198 8274 9199
rect 8750 9505 8778 9506
rect 8750 9479 8751 9505
rect 8751 9479 8777 9505
rect 8777 9479 8778 9505
rect 8750 9478 8778 9479
rect 8806 9310 8834 9338
rect 9086 9729 9114 9730
rect 9086 9703 9087 9729
rect 9087 9703 9113 9729
rect 9113 9703 9114 9729
rect 9086 9702 9114 9703
rect 8694 9254 8722 9282
rect 9590 9758 9618 9786
rect 9478 9646 9506 9674
rect 9142 9617 9170 9618
rect 9142 9591 9143 9617
rect 9143 9591 9169 9617
rect 9169 9591 9170 9617
rect 9142 9590 9170 9591
rect 9086 9505 9114 9506
rect 9086 9479 9087 9505
rect 9087 9479 9113 9505
rect 9113 9479 9114 9505
rect 9086 9478 9114 9479
rect 9030 9254 9058 9282
rect 9142 9198 9170 9226
rect 9478 9310 9506 9338
rect 9366 9030 9394 9058
rect 8470 8694 8498 8722
rect 9030 8526 9058 8554
rect 8078 8414 8106 8442
rect 9478 9225 9506 9226
rect 9478 9199 9479 9225
rect 9479 9199 9505 9225
rect 9505 9199 9506 9225
rect 9478 9198 9506 9199
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 9814 11550 9842 11578
rect 9814 11214 9842 11242
rect 10318 11214 10346 11242
rect 10654 11214 10682 11242
rect 11606 13873 11634 13874
rect 11606 13847 11607 13873
rect 11607 13847 11633 13873
rect 11633 13847 11634 13873
rect 11606 13846 11634 13847
rect 11606 13454 11634 13482
rect 11214 13398 11242 13426
rect 11550 13398 11578 13426
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 11998 14238 12026 14266
rect 12110 13846 12138 13874
rect 11606 12753 11634 12754
rect 11606 12727 11607 12753
rect 11607 12727 11633 12753
rect 11633 12727 11634 12753
rect 11606 12726 11634 12727
rect 10766 12614 10794 12642
rect 10990 12446 11018 12474
rect 11046 12614 11074 12642
rect 10206 11073 10234 11074
rect 10206 11047 10207 11073
rect 10207 11047 10233 11073
rect 10233 11047 10234 11073
rect 10206 11046 10234 11047
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 10150 10990 10178 11018
rect 10038 10905 10066 10906
rect 10038 10879 10039 10905
rect 10039 10879 10065 10905
rect 10065 10879 10066 10905
rect 10038 10878 10066 10879
rect 9646 10766 9674 10794
rect 9982 10793 10010 10794
rect 9982 10767 9983 10793
rect 9983 10767 10009 10793
rect 10009 10767 10010 10793
rect 9982 10766 10010 10767
rect 10318 10318 10346 10346
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9814 10038 9842 10066
rect 9702 9926 9730 9954
rect 9646 9198 9674 9226
rect 9590 9142 9618 9170
rect 9478 8750 9506 8778
rect 9534 8721 9562 8722
rect 9534 8695 9535 8721
rect 9535 8695 9561 8721
rect 9561 8695 9562 8721
rect 9534 8694 9562 8695
rect 8414 8105 8442 8106
rect 8414 8079 8415 8105
rect 8415 8079 8441 8105
rect 8441 8079 8442 8105
rect 8414 8078 8442 8079
rect 7798 7686 7826 7714
rect 8974 7713 9002 7714
rect 8974 7687 8975 7713
rect 8975 7687 9001 7713
rect 9001 7687 9002 7713
rect 8974 7686 9002 7687
rect 7910 7265 7938 7266
rect 7910 7239 7911 7265
rect 7911 7239 7937 7265
rect 7937 7239 7938 7265
rect 7910 7238 7938 7239
rect 7742 6958 7770 6986
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 8134 6734 8162 6762
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9646 7993 9674 7994
rect 9646 7967 9647 7993
rect 9647 7967 9673 7993
rect 9673 7967 9674 7993
rect 9646 7966 9674 7967
rect 9030 7126 9058 7154
rect 9310 7574 9338 7602
rect 9254 7238 9282 7266
rect 9702 7854 9730 7882
rect 9870 10094 9898 10122
rect 10542 11046 10570 11074
rect 9926 9702 9954 9730
rect 10206 9729 10234 9730
rect 10206 9703 10207 9729
rect 10207 9703 10233 9729
rect 10233 9703 10234 9729
rect 10206 9702 10234 9703
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9870 9254 9898 9282
rect 10206 9505 10234 9506
rect 10206 9479 10207 9505
rect 10207 9479 10233 9505
rect 10233 9479 10234 9505
rect 10206 9478 10234 9479
rect 10150 9310 10178 9338
rect 9870 9142 9898 9170
rect 9870 9030 9898 9058
rect 10150 8777 10178 8778
rect 10150 8751 10151 8777
rect 10151 8751 10177 8777
rect 10177 8751 10178 8777
rect 10150 8750 10178 8751
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 10206 8358 10234 8386
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 9926 7742 9954 7770
rect 9646 7630 9674 7658
rect 10318 7657 10346 7658
rect 10318 7631 10319 7657
rect 10319 7631 10345 7657
rect 10345 7631 10346 7657
rect 10318 7630 10346 7631
rect 9926 7574 9954 7602
rect 9702 7153 9730 7154
rect 9702 7127 9703 7153
rect 9703 7127 9729 7153
rect 9729 7127 9730 7153
rect 9702 7126 9730 7127
rect 9254 6985 9282 6986
rect 9254 6959 9255 6985
rect 9255 6959 9281 6985
rect 9281 6959 9282 6985
rect 9254 6958 9282 6959
rect 9478 6958 9506 6986
rect 8862 6761 8890 6762
rect 8862 6735 8863 6761
rect 8863 6735 8889 6761
rect 8889 6735 8890 6761
rect 8862 6734 8890 6735
rect 9198 6537 9226 6538
rect 9198 6511 9199 6537
rect 9199 6511 9225 6537
rect 9225 6511 9226 6537
rect 9198 6510 9226 6511
rect 9534 6510 9562 6538
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 10990 11241 11018 11242
rect 10990 11215 10991 11241
rect 10991 11215 11017 11241
rect 11017 11215 11018 11241
rect 10990 11214 11018 11215
rect 11550 12641 11578 12642
rect 11550 12615 11551 12641
rect 11551 12615 11577 12641
rect 11577 12615 11578 12641
rect 11550 12614 11578 12615
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 12334 13089 12362 13090
rect 12334 13063 12335 13089
rect 12335 13063 12361 13089
rect 12361 13063 12362 13089
rect 12334 13062 12362 13063
rect 11942 12726 11970 12754
rect 13174 13398 13202 13426
rect 12558 13062 12586 13090
rect 12726 13062 12754 13090
rect 11830 12614 11858 12642
rect 12110 12641 12138 12642
rect 12110 12615 12111 12641
rect 12111 12615 12137 12641
rect 12137 12615 12138 12641
rect 12110 12614 12138 12615
rect 12838 12614 12866 12642
rect 12614 12361 12642 12362
rect 12614 12335 12615 12361
rect 12615 12335 12641 12361
rect 12641 12335 12642 12361
rect 12614 12334 12642 12335
rect 12054 11633 12082 11634
rect 12054 11607 12055 11633
rect 12055 11607 12081 11633
rect 12081 11607 12082 11633
rect 12054 11606 12082 11607
rect 11942 11577 11970 11578
rect 11942 11551 11943 11577
rect 11943 11551 11969 11577
rect 11969 11551 11970 11577
rect 11942 11550 11970 11551
rect 12110 11270 12138 11298
rect 11270 11102 11298 11130
rect 11550 11102 11578 11130
rect 11046 10990 11074 11018
rect 11494 10878 11522 10906
rect 11942 10878 11970 10906
rect 11494 10793 11522 10794
rect 11494 10767 11495 10793
rect 11495 10767 11521 10793
rect 11521 10767 11522 10793
rect 11494 10766 11522 10767
rect 10710 10065 10738 10066
rect 10710 10039 10711 10065
rect 10711 10039 10737 10065
rect 10737 10039 10738 10065
rect 10710 10038 10738 10039
rect 11158 10345 11186 10346
rect 11158 10319 11159 10345
rect 11159 10319 11185 10345
rect 11185 10319 11186 10345
rect 11158 10318 11186 10319
rect 10822 9982 10850 10010
rect 11102 10094 11130 10122
rect 10654 9702 10682 9730
rect 10654 9478 10682 9506
rect 10598 9142 10626 9170
rect 10934 9225 10962 9226
rect 10934 9199 10935 9225
rect 10935 9199 10961 9225
rect 10961 9199 10962 9225
rect 10934 9198 10962 9199
rect 10822 8777 10850 8778
rect 10822 8751 10823 8777
rect 10823 8751 10849 8777
rect 10849 8751 10850 8777
rect 10822 8750 10850 8751
rect 11326 9366 11354 9394
rect 11382 9337 11410 9338
rect 11382 9311 11383 9337
rect 11383 9311 11409 9337
rect 11409 9311 11410 9337
rect 11382 9310 11410 9311
rect 11214 9281 11242 9282
rect 11214 9255 11215 9281
rect 11215 9255 11241 9281
rect 11241 9255 11242 9281
rect 11214 9254 11242 9255
rect 11494 10150 11522 10178
rect 11438 9142 11466 9170
rect 12054 10766 12082 10794
rect 12278 10878 12306 10906
rect 12334 10793 12362 10794
rect 12334 10767 12335 10793
rect 12335 10767 12361 10793
rect 12361 10767 12362 10793
rect 12334 10766 12362 10767
rect 11942 10038 11970 10066
rect 12558 10065 12586 10066
rect 12558 10039 12559 10065
rect 12559 10039 12585 10065
rect 12585 10039 12586 10065
rect 12558 10038 12586 10039
rect 12782 10934 12810 10962
rect 13062 12473 13090 12474
rect 13062 12447 13063 12473
rect 13063 12447 13089 12473
rect 13089 12447 13090 12473
rect 13062 12446 13090 12447
rect 13230 13062 13258 13090
rect 12950 12390 12978 12418
rect 13174 12361 13202 12362
rect 13174 12335 13175 12361
rect 13175 12335 13201 12361
rect 13201 12335 13202 12361
rect 13174 12334 13202 12335
rect 18830 13230 18858 13258
rect 14518 13201 14546 13202
rect 14518 13175 14519 13201
rect 14519 13175 14545 13201
rect 14545 13175 14546 13201
rect 14518 13174 14546 13175
rect 14406 13145 14434 13146
rect 14406 13119 14407 13145
rect 14407 13119 14433 13145
rect 14433 13119 14434 13145
rect 14406 13118 14434 13119
rect 18830 13145 18858 13146
rect 18830 13119 18831 13145
rect 18831 13119 18857 13145
rect 18857 13119 18858 13145
rect 18830 13118 18858 13119
rect 13958 13062 13986 13090
rect 13734 12726 13762 12754
rect 13510 12614 13538 12642
rect 13454 12446 13482 12474
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 18830 12753 18858 12754
rect 18830 12727 18831 12753
rect 18831 12727 18857 12753
rect 18857 12727 18858 12753
rect 18830 12726 18858 12727
rect 14070 12641 14098 12642
rect 14070 12615 14071 12641
rect 14071 12615 14097 12641
rect 14097 12615 14098 12641
rect 14070 12614 14098 12615
rect 19950 13454 19978 13482
rect 20006 13118 20034 13146
rect 19950 12782 19978 12810
rect 18942 12614 18970 12642
rect 20006 12446 20034 12474
rect 13678 12417 13706 12418
rect 13678 12391 13679 12417
rect 13679 12391 13705 12417
rect 13705 12391 13706 12417
rect 13678 12390 13706 12391
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 20006 12110 20034 12138
rect 20006 11774 20034 11802
rect 18942 11606 18970 11634
rect 18774 11550 18802 11578
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 20006 11465 20034 11466
rect 20006 11439 20007 11465
rect 20007 11439 20033 11465
rect 20033 11439 20034 11465
rect 20006 11438 20034 11439
rect 13342 10934 13370 10962
rect 13062 10878 13090 10906
rect 12670 10793 12698 10794
rect 12670 10767 12671 10793
rect 12671 10767 12697 10793
rect 12697 10767 12698 10793
rect 12670 10766 12698 10767
rect 12614 9982 12642 10010
rect 12670 9758 12698 9786
rect 11886 9366 11914 9394
rect 11494 9198 11522 9226
rect 11550 8918 11578 8946
rect 11942 8889 11970 8890
rect 11942 8863 11943 8889
rect 11943 8863 11969 8889
rect 11969 8863 11970 8889
rect 11942 8862 11970 8863
rect 12278 8974 12306 9002
rect 12222 8945 12250 8946
rect 12222 8919 12223 8945
rect 12223 8919 12249 8945
rect 12249 8919 12250 8945
rect 12222 8918 12250 8919
rect 12838 9870 12866 9898
rect 12782 9758 12810 9786
rect 12334 8862 12362 8890
rect 12558 8918 12586 8946
rect 11942 8750 11970 8778
rect 10990 8414 11018 8442
rect 11774 8526 11802 8554
rect 10878 8358 10906 8386
rect 10542 7966 10570 7994
rect 10822 8049 10850 8050
rect 10822 8023 10823 8049
rect 10823 8023 10849 8049
rect 10849 8023 10850 8049
rect 10822 8022 10850 8023
rect 10654 7742 10682 7770
rect 10542 7630 10570 7658
rect 11774 8358 11802 8386
rect 11886 8049 11914 8050
rect 11886 8023 11887 8049
rect 11887 8023 11913 8049
rect 11913 8023 11914 8049
rect 11886 8022 11914 8023
rect 11550 7966 11578 7994
rect 11830 7937 11858 7938
rect 11830 7911 11831 7937
rect 11831 7911 11857 7937
rect 11857 7911 11858 7937
rect 11830 7910 11858 7911
rect 12390 8721 12418 8722
rect 12390 8695 12391 8721
rect 12391 8695 12417 8721
rect 12417 8695 12418 8721
rect 12390 8694 12418 8695
rect 12166 8414 12194 8442
rect 12726 8862 12754 8890
rect 12838 9254 12866 9282
rect 13790 11129 13818 11130
rect 13790 11103 13791 11129
rect 13791 11103 13817 11129
rect 13817 11103 13818 11129
rect 13790 11102 13818 11103
rect 14014 11046 14042 11074
rect 14630 11046 14658 11074
rect 13006 9982 13034 10010
rect 14966 11046 14994 11074
rect 18774 11046 18802 11074
rect 20006 11102 20034 11130
rect 18830 10934 18858 10962
rect 15078 10766 15106 10794
rect 18830 10793 18858 10794
rect 18830 10767 18831 10793
rect 18831 10767 18857 10793
rect 18857 10767 18858 10793
rect 18830 10766 18858 10767
rect 20006 10766 20034 10794
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 20006 10457 20034 10458
rect 20006 10431 20007 10457
rect 20007 10431 20033 10457
rect 20033 10431 20034 10457
rect 20006 10430 20034 10431
rect 14742 10374 14770 10402
rect 18830 10401 18858 10402
rect 18830 10375 18831 10401
rect 18831 10375 18857 10401
rect 18857 10375 18858 10401
rect 18830 10374 18858 10375
rect 13286 9870 13314 9898
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 13286 9758 13314 9786
rect 13062 9225 13090 9226
rect 13062 9199 13063 9225
rect 13063 9199 13089 9225
rect 13089 9199 13090 9225
rect 13062 9198 13090 9199
rect 12894 8974 12922 9002
rect 12670 8694 12698 8722
rect 12670 8441 12698 8442
rect 12670 8415 12671 8441
rect 12671 8415 12697 8441
rect 12697 8415 12698 8441
rect 12670 8414 12698 8415
rect 12894 8414 12922 8442
rect 13006 8694 13034 8722
rect 13230 9225 13258 9226
rect 13230 9199 13231 9225
rect 13231 9199 13257 9225
rect 13257 9199 13258 9225
rect 13230 9198 13258 9199
rect 13118 8385 13146 8386
rect 13118 8359 13119 8385
rect 13119 8359 13145 8385
rect 13145 8359 13146 8385
rect 13118 8358 13146 8359
rect 13174 8974 13202 9002
rect 12614 8022 12642 8050
rect 12614 7910 12642 7938
rect 12726 7854 12754 7882
rect 13230 8777 13258 8778
rect 13230 8751 13231 8777
rect 13231 8751 13257 8777
rect 13257 8751 13258 8777
rect 13230 8750 13258 8751
rect 14238 9617 14266 9618
rect 14238 9591 14239 9617
rect 14239 9591 14265 9617
rect 14265 9591 14266 9617
rect 14238 9590 14266 9591
rect 14686 9590 14714 9618
rect 18830 9617 18858 9618
rect 18830 9591 18831 9617
rect 18831 9591 18857 9617
rect 18857 9591 18858 9617
rect 18830 9590 18858 9591
rect 20006 9422 20034 9450
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 14294 8889 14322 8890
rect 14294 8863 14295 8889
rect 14295 8863 14321 8889
rect 14321 8863 14322 8889
rect 14294 8862 14322 8863
rect 14630 8889 14658 8890
rect 14630 8863 14631 8889
rect 14631 8863 14657 8889
rect 14657 8863 14658 8889
rect 14630 8862 14658 8863
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 13398 8750 13426 8778
rect 20006 8750 20034 8778
rect 13454 8694 13482 8722
rect 14574 8721 14602 8722
rect 14574 8695 14575 8721
rect 14575 8695 14601 8721
rect 14601 8695 14602 8721
rect 14574 8694 14602 8695
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 13230 7854 13258 7882
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 13118 7294 13146 7322
rect 10654 6958 10682 6986
rect 11158 6985 11186 6986
rect 11158 6959 11159 6985
rect 11159 6959 11185 6985
rect 11185 6959 11186 6985
rect 11158 6958 11186 6959
rect 12110 6985 12138 6986
rect 12110 6959 12111 6985
rect 12111 6959 12137 6985
rect 12137 6959 12138 6985
rect 12110 6958 12138 6959
rect 10542 6734 10570 6762
rect 9758 6510 9786 6538
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9422 2030 9450 2058
rect 10038 2057 10066 2058
rect 10038 2031 10039 2057
rect 10039 2031 10065 2057
rect 10065 2031 10066 2057
rect 10038 2030 10066 2031
rect 10430 1806 10458 1834
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 10934 6734 10962 6762
rect 13734 7321 13762 7322
rect 13734 7295 13735 7321
rect 13735 7295 13761 7321
rect 13761 7295 13762 7321
rect 13734 7294 13762 7295
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 13118 2030 13146 2058
rect 11046 1833 11074 1834
rect 11046 1807 11047 1833
rect 11047 1807 11073 1833
rect 11073 1807 11074 1833
rect 11046 1806 11074 1807
rect 13734 2057 13762 2058
rect 13734 2031 13735 2057
rect 13735 2031 13761 2057
rect 13761 2031 13762 2057
rect 13734 2030 13762 2031
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
<< metal3 >>
rect 9753 19278 9758 19306
rect 9786 19278 10374 19306
rect 10402 19278 10407 19306
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 11769 19110 11774 19138
rect 11802 19110 12782 19138
rect 12810 19110 12815 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9081 18326 9086 18354
rect 9114 18326 9590 18354
rect 9618 18326 9623 18354
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 11321 14238 11326 14266
rect 11354 14238 11998 14266
rect 12026 14238 12031 14266
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 11601 13846 11606 13874
rect 11634 13846 12110 13874
rect 12138 13846 12143 13874
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 8465 13510 8470 13538
rect 8498 13510 9926 13538
rect 9954 13510 9959 13538
rect 0 13482 400 13496
rect 0 13454 2086 13482
rect 2114 13454 2119 13482
rect 0 13440 400 13454
rect 8470 13426 8498 13510
rect 20600 13482 21000 13496
rect 10934 13454 11606 13482
rect 11634 13454 11639 13482
rect 19945 13454 19950 13482
rect 19978 13454 21000 13482
rect 10934 13426 10962 13454
rect 20600 13440 21000 13454
rect 7513 13398 7518 13426
rect 7546 13398 7910 13426
rect 7938 13398 8498 13426
rect 10089 13398 10094 13426
rect 10122 13398 10486 13426
rect 10514 13398 10962 13426
rect 11209 13398 11214 13426
rect 11242 13398 11550 13426
rect 11578 13398 13174 13426
rect 13202 13398 13207 13426
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 11214 13202 11242 13398
rect 15946 13230 18830 13258
rect 18858 13230 18863 13258
rect 15946 13202 15974 13230
rect 9809 13174 9814 13202
rect 9842 13174 11242 13202
rect 14513 13174 14518 13202
rect 14546 13174 15974 13202
rect 20600 13146 21000 13160
rect 8633 13118 8638 13146
rect 8666 13118 9254 13146
rect 9282 13118 9287 13146
rect 9417 13118 9422 13146
rect 9450 13118 9702 13146
rect 9730 13118 9735 13146
rect 14401 13118 14406 13146
rect 14434 13118 18830 13146
rect 18858 13118 18863 13146
rect 20001 13118 20006 13146
rect 20034 13118 21000 13146
rect 20600 13104 21000 13118
rect 2137 13062 2142 13090
rect 2170 13062 5838 13090
rect 5866 13062 5871 13090
rect 8241 13062 8246 13090
rect 8274 13062 8918 13090
rect 8946 13062 8951 13090
rect 12329 13062 12334 13090
rect 12362 13062 12558 13090
rect 12586 13062 12726 13090
rect 12754 13062 12759 13090
rect 13225 13062 13230 13090
rect 13258 13062 13958 13090
rect 13986 13062 13991 13090
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 20600 12810 21000 12824
rect 19945 12782 19950 12810
rect 19978 12782 21000 12810
rect 20600 12768 21000 12782
rect 11601 12726 11606 12754
rect 11634 12726 11942 12754
rect 11970 12726 11975 12754
rect 13729 12726 13734 12754
rect 13762 12726 18830 12754
rect 18858 12726 18863 12754
rect 5833 12670 5838 12698
rect 5866 12670 7350 12698
rect 7378 12670 7383 12698
rect 10761 12614 10766 12642
rect 10794 12614 11046 12642
rect 11074 12614 11079 12642
rect 11545 12614 11550 12642
rect 11578 12614 11830 12642
rect 11858 12614 11863 12642
rect 12105 12614 12110 12642
rect 12138 12614 12838 12642
rect 12866 12614 13510 12642
rect 13538 12614 13543 12642
rect 14065 12614 14070 12642
rect 14098 12614 18942 12642
rect 18970 12614 18975 12642
rect 6897 12558 6902 12586
rect 6930 12558 7686 12586
rect 7714 12558 7719 12586
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 0 12474 400 12488
rect 20600 12474 21000 12488
rect 0 12446 966 12474
rect 994 12446 999 12474
rect 7513 12446 7518 12474
rect 7546 12446 7551 12474
rect 10985 12446 10990 12474
rect 11018 12446 13062 12474
rect 13090 12446 13454 12474
rect 13482 12446 13487 12474
rect 20001 12446 20006 12474
rect 20034 12446 21000 12474
rect 0 12432 400 12446
rect 7518 12362 7546 12446
rect 20600 12432 21000 12446
rect 7793 12390 7798 12418
rect 7826 12390 8694 12418
rect 8722 12390 9142 12418
rect 9170 12390 9175 12418
rect 12945 12390 12950 12418
rect 12978 12390 13678 12418
rect 13706 12390 13711 12418
rect 2137 12334 2142 12362
rect 2170 12334 6006 12362
rect 6034 12334 7546 12362
rect 7905 12334 7910 12362
rect 7938 12334 8750 12362
rect 8778 12334 8783 12362
rect 9697 12334 9702 12362
rect 9730 12334 12614 12362
rect 12642 12334 13174 12362
rect 13202 12334 13207 12362
rect 7065 12278 7070 12306
rect 7098 12278 7742 12306
rect 7770 12278 7775 12306
rect 961 12222 966 12250
rect 994 12222 999 12250
rect 7177 12222 7182 12250
rect 7210 12222 7406 12250
rect 7434 12222 8134 12250
rect 8162 12222 8167 12250
rect 0 12138 400 12152
rect 966 12138 994 12222
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 20600 12138 21000 12152
rect 0 12110 994 12138
rect 7569 12110 7574 12138
rect 7602 12110 7910 12138
rect 7938 12110 7943 12138
rect 20001 12110 20006 12138
rect 20034 12110 21000 12138
rect 0 12096 400 12110
rect 20600 12096 21000 12110
rect 20600 11802 21000 11816
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 20600 11760 21000 11774
rect 8969 11662 8974 11690
rect 9002 11662 9646 11690
rect 9674 11662 9679 11690
rect 9081 11606 9086 11634
rect 9114 11606 9366 11634
rect 9394 11606 9590 11634
rect 9618 11606 9623 11634
rect 12049 11606 12054 11634
rect 12082 11606 18942 11634
rect 18970 11606 18975 11634
rect 2137 11550 2142 11578
rect 2170 11550 4214 11578
rect 6169 11550 6174 11578
rect 6202 11550 7182 11578
rect 7210 11550 7518 11578
rect 7546 11550 7551 11578
rect 9417 11550 9422 11578
rect 9450 11550 9814 11578
rect 9842 11550 9847 11578
rect 11937 11550 11942 11578
rect 11970 11550 18774 11578
rect 18802 11550 18807 11578
rect 4186 11522 4214 11550
rect 4186 11494 5726 11522
rect 5754 11494 5759 11522
rect 6785 11494 6790 11522
rect 6818 11494 7574 11522
rect 7602 11494 7607 11522
rect 0 11466 400 11480
rect 20600 11466 21000 11480
rect 0 11438 966 11466
rect 994 11438 999 11466
rect 20001 11438 20006 11466
rect 20034 11438 21000 11466
rect 0 11424 400 11438
rect 20600 11424 21000 11438
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 7681 11326 7686 11354
rect 7714 11326 9534 11354
rect 9562 11326 10094 11354
rect 10066 11298 10094 11326
rect 7905 11270 7910 11298
rect 7938 11270 8806 11298
rect 8834 11270 8839 11298
rect 10066 11270 12110 11298
rect 12138 11270 12143 11298
rect 9809 11214 9814 11242
rect 9842 11214 10318 11242
rect 10346 11214 10351 11242
rect 10649 11214 10654 11242
rect 10682 11214 10990 11242
rect 11018 11214 11023 11242
rect 20600 11130 21000 11144
rect 5721 11102 5726 11130
rect 5754 11102 7350 11130
rect 7378 11102 7383 11130
rect 9081 11102 9086 11130
rect 9114 11102 10094 11130
rect 11265 11102 11270 11130
rect 11298 11102 11550 11130
rect 11578 11102 13790 11130
rect 13818 11102 13823 11130
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 10066 11074 10094 11102
rect 20600 11088 21000 11102
rect 8689 11046 8694 11074
rect 8722 11046 9030 11074
rect 9058 11046 9063 11074
rect 9585 11046 9590 11074
rect 9618 11046 9623 11074
rect 10066 11046 10206 11074
rect 10234 11046 10542 11074
rect 10570 11046 10575 11074
rect 14009 11046 14014 11074
rect 14042 11046 14630 11074
rect 14658 11046 14966 11074
rect 14994 11046 18774 11074
rect 18802 11046 18807 11074
rect 9590 10962 9618 11046
rect 10145 10990 10150 11018
rect 10178 10990 11046 11018
rect 11074 10990 11079 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 8857 10934 8862 10962
rect 8890 10934 9618 10962
rect 12777 10934 12782 10962
rect 12810 10934 13342 10962
rect 13370 10934 18830 10962
rect 18858 10934 18863 10962
rect 8862 10850 8890 10934
rect 9590 10906 9618 10934
rect 9590 10878 10038 10906
rect 10066 10878 10071 10906
rect 11489 10878 11494 10906
rect 11522 10878 11942 10906
rect 11970 10878 12278 10906
rect 12306 10878 13062 10906
rect 13090 10878 13095 10906
rect 6505 10822 6510 10850
rect 6538 10822 7910 10850
rect 7938 10822 8890 10850
rect 20600 10794 21000 10808
rect 7569 10766 7574 10794
rect 7602 10766 7966 10794
rect 7994 10766 8694 10794
rect 8722 10766 8727 10794
rect 9641 10766 9646 10794
rect 9674 10766 9982 10794
rect 10010 10766 10015 10794
rect 11489 10766 11494 10794
rect 11522 10766 12054 10794
rect 12082 10766 12087 10794
rect 12329 10766 12334 10794
rect 12362 10766 12670 10794
rect 12698 10766 12703 10794
rect 15073 10766 15078 10794
rect 15106 10766 18830 10794
rect 18858 10766 18863 10794
rect 20001 10766 20006 10794
rect 20034 10766 21000 10794
rect 20600 10752 21000 10766
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 20600 10458 21000 10472
rect 20001 10430 20006 10458
rect 20034 10430 21000 10458
rect 20600 10416 21000 10430
rect 14737 10374 14742 10402
rect 14770 10374 18830 10402
rect 18858 10374 18863 10402
rect 10313 10318 10318 10346
rect 10346 10318 11158 10346
rect 11186 10318 11191 10346
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 11489 10150 11494 10178
rect 11522 10150 11527 10178
rect 11494 10122 11522 10150
rect 9529 10094 9534 10122
rect 9562 10094 9870 10122
rect 9898 10094 11102 10122
rect 11130 10094 11522 10122
rect 9809 10038 9814 10066
rect 9842 10038 10710 10066
rect 10738 10038 10743 10066
rect 11937 10038 11942 10066
rect 11970 10038 12558 10066
rect 12586 10038 12591 10066
rect 2137 9982 2142 10010
rect 2170 9982 5502 10010
rect 5530 9982 5535 10010
rect 8969 9982 8974 10010
rect 9002 9982 9366 10010
rect 9394 9982 9399 10010
rect 10817 9982 10822 10010
rect 10850 9982 12614 10010
rect 12642 9982 13006 10010
rect 13034 9982 13039 10010
rect 2081 9926 2086 9954
rect 2114 9926 9198 9954
rect 9226 9926 9702 9954
rect 9730 9926 9735 9954
rect 961 9870 966 9898
rect 994 9870 999 9898
rect 12833 9870 12838 9898
rect 12866 9870 13286 9898
rect 13314 9870 13319 9898
rect 0 9786 400 9800
rect 966 9786 994 9870
rect 5497 9814 5502 9842
rect 5530 9814 7182 9842
rect 7210 9814 7215 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 0 9758 994 9786
rect 8801 9758 8806 9786
rect 8834 9758 9590 9786
rect 9618 9758 9623 9786
rect 12665 9758 12670 9786
rect 12698 9758 12782 9786
rect 12810 9758 13286 9786
rect 13314 9758 13319 9786
rect 0 9744 400 9758
rect 7457 9702 7462 9730
rect 7490 9702 9086 9730
rect 9114 9702 9119 9730
rect 9921 9702 9926 9730
rect 9954 9702 10206 9730
rect 10234 9702 10654 9730
rect 10682 9702 10687 9730
rect 7905 9646 7910 9674
rect 7938 9646 8358 9674
rect 8386 9646 9478 9674
rect 9506 9646 9511 9674
rect 8521 9590 8526 9618
rect 8554 9590 9142 9618
rect 9170 9590 9175 9618
rect 14233 9590 14238 9618
rect 14266 9590 14686 9618
rect 14714 9590 18830 9618
rect 18858 9590 18863 9618
rect 6281 9534 6286 9562
rect 6314 9534 7126 9562
rect 7154 9534 7159 9562
rect 7233 9534 7238 9562
rect 7266 9534 7742 9562
rect 7770 9534 7775 9562
rect 8577 9534 8582 9562
rect 8610 9534 9114 9562
rect 9086 9506 9114 9534
rect 8073 9478 8078 9506
rect 8106 9478 8750 9506
rect 8778 9478 8783 9506
rect 9081 9478 9086 9506
rect 9114 9478 10206 9506
rect 10234 9478 10654 9506
rect 10682 9478 10687 9506
rect 20600 9450 21000 9464
rect 20001 9422 20006 9450
rect 20034 9422 21000 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 20600 9408 21000 9422
rect 11321 9366 11326 9394
rect 11354 9366 11886 9394
rect 11914 9366 11919 9394
rect 8801 9310 8806 9338
rect 8834 9310 8839 9338
rect 9473 9310 9478 9338
rect 9506 9310 10150 9338
rect 10178 9310 11382 9338
rect 11410 9310 11415 9338
rect 8409 9254 8414 9282
rect 8442 9254 8694 9282
rect 8722 9254 8727 9282
rect 8806 9226 8834 9310
rect 9025 9254 9030 9282
rect 9058 9254 9870 9282
rect 9898 9254 9903 9282
rect 9982 9254 11130 9282
rect 11209 9254 11214 9282
rect 11242 9254 12838 9282
rect 12866 9254 12871 9282
rect 9982 9226 10010 9254
rect 11102 9226 11130 9254
rect 7457 9198 7462 9226
rect 7490 9198 8246 9226
rect 8274 9198 8834 9226
rect 9137 9198 9142 9226
rect 9170 9198 9478 9226
rect 9506 9198 9646 9226
rect 9674 9198 9679 9226
rect 9758 9198 10010 9226
rect 10066 9198 10934 9226
rect 10962 9198 10967 9226
rect 11102 9198 11494 9226
rect 11522 9198 11527 9226
rect 13057 9198 13062 9226
rect 13090 9198 13230 9226
rect 13258 9198 13263 9226
rect 9758 9170 9786 9198
rect 10066 9170 10094 9198
rect 9585 9142 9590 9170
rect 9618 9142 9786 9170
rect 9865 9142 9870 9170
rect 9898 9142 10094 9170
rect 10593 9142 10598 9170
rect 10626 9142 11438 9170
rect 11466 9142 11471 9170
rect 10598 9114 10626 9142
rect 7065 9086 7070 9114
rect 7098 9086 7350 9114
rect 7378 9086 7742 9114
rect 7770 9086 10626 9114
rect 9361 9030 9366 9058
rect 9394 9030 9870 9058
rect 9898 9030 9903 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 12273 8974 12278 9002
rect 12306 8974 12894 9002
rect 12922 8974 13174 9002
rect 13202 8974 13207 9002
rect 11545 8918 11550 8946
rect 11578 8918 12222 8946
rect 12250 8918 12558 8946
rect 12586 8918 12591 8946
rect 11937 8862 11942 8890
rect 11970 8862 12334 8890
rect 12362 8862 12726 8890
rect 12754 8862 12759 8890
rect 14289 8862 14294 8890
rect 14322 8862 14630 8890
rect 14658 8862 15974 8890
rect 15946 8834 15974 8862
rect 2137 8806 2142 8834
rect 2170 8806 4214 8834
rect 7401 8806 7406 8834
rect 7434 8806 7854 8834
rect 7882 8806 7887 8834
rect 15946 8806 18830 8834
rect 18858 8806 18863 8834
rect 4186 8778 4214 8806
rect 20600 8778 21000 8792
rect 4186 8750 7910 8778
rect 7938 8750 7943 8778
rect 9473 8750 9478 8778
rect 9506 8750 10150 8778
rect 10178 8750 10183 8778
rect 10817 8750 10822 8778
rect 10850 8750 11942 8778
rect 11970 8750 11975 8778
rect 13225 8750 13230 8778
rect 13258 8750 13398 8778
rect 13426 8750 13431 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 20600 8736 21000 8750
rect 7233 8694 7238 8722
rect 7266 8694 7854 8722
rect 7882 8694 7887 8722
rect 8465 8694 8470 8722
rect 8498 8694 9534 8722
rect 9562 8694 9567 8722
rect 12385 8694 12390 8722
rect 12418 8694 12670 8722
rect 12698 8694 13006 8722
rect 13034 8694 13039 8722
rect 13449 8694 13454 8722
rect 13482 8694 14574 8722
rect 14602 8694 14607 8722
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 6953 8526 6958 8554
rect 6986 8526 7518 8554
rect 7546 8526 7551 8554
rect 7961 8526 7966 8554
rect 7994 8526 9030 8554
rect 9058 8526 11774 8554
rect 11802 8526 11807 8554
rect 6337 8470 6342 8498
rect 6370 8470 7406 8498
rect 7434 8470 7439 8498
rect 0 8442 400 8456
rect 0 8414 966 8442
rect 994 8414 999 8442
rect 6001 8414 6006 8442
rect 6034 8414 6790 8442
rect 6818 8414 6823 8442
rect 8073 8414 8078 8442
rect 8106 8414 8111 8442
rect 10985 8414 10990 8442
rect 11018 8414 12166 8442
rect 12194 8414 12670 8442
rect 12698 8414 12894 8442
rect 12922 8414 12927 8442
rect 0 8400 400 8414
rect 8078 8386 8106 8414
rect 7793 8358 7798 8386
rect 7826 8358 8106 8386
rect 10201 8358 10206 8386
rect 10234 8358 10878 8386
rect 10906 8358 10911 8386
rect 11769 8358 11774 8386
rect 11802 8358 13118 8386
rect 13146 8358 13151 8386
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 7569 8078 7574 8106
rect 7602 8078 8414 8106
rect 8442 8078 8447 8106
rect 10817 8022 10822 8050
rect 10850 8022 11886 8050
rect 11914 8022 12614 8050
rect 12642 8022 12647 8050
rect 9641 7966 9646 7994
rect 9674 7966 10094 7994
rect 10537 7966 10542 7994
rect 10570 7966 11550 7994
rect 11578 7966 11583 7994
rect 10066 7938 10094 7966
rect 10066 7910 11746 7938
rect 11825 7910 11830 7938
rect 11858 7910 12614 7938
rect 12642 7910 12647 7938
rect 11718 7882 11746 7910
rect 9697 7854 9702 7882
rect 9730 7854 9735 7882
rect 11718 7854 12726 7882
rect 12754 7854 13230 7882
rect 13258 7854 13263 7882
rect 9702 7770 9730 7854
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 9702 7742 9926 7770
rect 9954 7742 10654 7770
rect 10682 7742 10687 7770
rect 7793 7686 7798 7714
rect 7826 7686 8974 7714
rect 9002 7686 9007 7714
rect 9641 7630 9646 7658
rect 9674 7630 10318 7658
rect 10346 7630 10542 7658
rect 10570 7630 10575 7658
rect 9305 7574 9310 7602
rect 9338 7574 9926 7602
rect 9954 7574 9959 7602
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 13113 7294 13118 7322
rect 13146 7294 13734 7322
rect 13762 7294 13767 7322
rect 7905 7238 7910 7266
rect 7938 7238 9254 7266
rect 9282 7238 9287 7266
rect 9025 7126 9030 7154
rect 9058 7126 9702 7154
rect 9730 7126 9735 7154
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 7737 6958 7742 6986
rect 7770 6958 9254 6986
rect 9282 6958 9478 6986
rect 9506 6958 10654 6986
rect 10682 6958 11158 6986
rect 11186 6958 12110 6986
rect 12138 6958 12143 6986
rect 8129 6734 8134 6762
rect 8162 6734 8862 6762
rect 8890 6734 8895 6762
rect 10537 6734 10542 6762
rect 10570 6734 10934 6762
rect 10962 6734 10967 6762
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9193 6510 9198 6538
rect 9226 6510 9534 6538
rect 9562 6510 9758 6538
rect 9786 6510 9791 6538
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 9417 2030 9422 2058
rect 9450 2030 10038 2058
rect 10066 2030 10071 2058
rect 13113 2030 13118 2058
rect 13146 2030 13734 2058
rect 13762 2030 13767 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 10425 1806 10430 1834
rect 10458 1806 11046 1834
rect 11074 1806 11079 1834
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _094_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12880 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _095_
timestamp 1698175906
transform -1 0 11648 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _096_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8008 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _097_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7392 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _098_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8064 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _099_
timestamp 1698175906
transform 1 0 8960 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12040 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _101_
timestamp 1698175906
transform -1 0 11424 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _102_
timestamp 1698175906
transform -1 0 10472 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9184 0 1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _104_
timestamp 1698175906
transform -1 0 12208 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1698175906
transform -1 0 10920 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _106_
timestamp 1698175906
transform -1 0 8960 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7952 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _108_
timestamp 1698175906
transform 1 0 8176 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_
timestamp 1698175906
transform 1 0 8904 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _110_
timestamp 1698175906
transform 1 0 9912 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _111_
timestamp 1698175906
transform 1 0 10080 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11816 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1698175906
transform -1 0 12208 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _115_
timestamp 1698175906
transform -1 0 11312 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7224 0 -1 10192
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _118_
timestamp 1698175906
transform -1 0 7672 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _119_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698175906
transform 1 0 9296 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12040 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _122_
timestamp 1698175906
transform 1 0 12600 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9240 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _124_
timestamp 1698175906
transform -1 0 11312 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _126_
timestamp 1698175906
transform 1 0 8288 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _127_
timestamp 1698175906
transform -1 0 9240 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _128_
timestamp 1698175906
transform 1 0 9800 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _129_
timestamp 1698175906
transform 1 0 9912 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _130_
timestamp 1698175906
transform 1 0 10808 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform 1 0 9464 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform 1 0 8792 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _133_
timestamp 1698175906
transform -1 0 12096 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _134_
timestamp 1698175906
transform 1 0 12488 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _135_
timestamp 1698175906
transform -1 0 14336 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _136_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12936 0 1 9408
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8792 0 -1 11760
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform 1 0 7224 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _139_
timestamp 1698175906
transform 1 0 7560 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _140_
timestamp 1698175906
transform -1 0 11704 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _141_
timestamp 1698175906
transform 1 0 10920 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform 1 0 9520 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _143_
timestamp 1698175906
transform 1 0 13104 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _144_
timestamp 1698175906
transform 1 0 12992 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _145_
timestamp 1698175906
transform -1 0 14728 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _146_
timestamp 1698175906
transform 1 0 12936 0 -1 8624
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _147_
timestamp 1698175906
transform -1 0 11704 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_
timestamp 1698175906
transform -1 0 9352 0 -1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _149_
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _150_
timestamp 1698175906
transform -1 0 8456 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _151_
timestamp 1698175906
transform 1 0 8400 0 1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _152_
timestamp 1698175906
transform -1 0 9072 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _153_
timestamp 1698175906
transform -1 0 10864 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _154_
timestamp 1698175906
transform -1 0 8904 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _155_
timestamp 1698175906
transform 1 0 7728 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _156_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8176 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _157_
timestamp 1698175906
transform 1 0 7168 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _158_
timestamp 1698175906
transform -1 0 10920 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _159_
timestamp 1698175906
transform -1 0 9688 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform 1 0 10024 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _161_
timestamp 1698175906
transform 1 0 10248 0 -1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _162_
timestamp 1698175906
transform 1 0 9744 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _163_
timestamp 1698175906
transform -1 0 9912 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _164_
timestamp 1698175906
transform -1 0 9464 0 -1 13328
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _165_
timestamp 1698175906
transform 1 0 11368 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _166_
timestamp 1698175906
transform -1 0 12824 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _167_
timestamp 1698175906
transform 1 0 11424 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _168_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11368 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _169_
timestamp 1698175906
transform -1 0 14112 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _170_
timestamp 1698175906
transform 1 0 13440 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _171_
timestamp 1698175906
transform 1 0 13440 0 -1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _172_
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _173_
timestamp 1698175906
transform -1 0 9912 0 1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _174_
timestamp 1698175906
transform 1 0 7224 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _175_
timestamp 1698175906
transform 1 0 7448 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _176_
timestamp 1698175906
transform 1 0 9576 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _177_
timestamp 1698175906
transform -1 0 9128 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _178_
timestamp 1698175906
transform 1 0 8904 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _179_
timestamp 1698175906
transform -1 0 9800 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _180_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9576 0 1 7056
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _181_
timestamp 1698175906
transform -1 0 12936 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _182_
timestamp 1698175906
transform 1 0 11872 0 -1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _183_
timestamp 1698175906
transform -1 0 11984 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _184_
timestamp 1698175906
transform -1 0 13272 0 -1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _185_
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _186_
timestamp 1698175906
transform 1 0 7000 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _187_
timestamp 1698175906
transform 1 0 6216 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _188_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7560 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _189_
timestamp 1698175906
transform 1 0 9800 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _190_
timestamp 1698175906
transform 1 0 6048 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _191_
timestamp 1698175906
transform 1 0 5880 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _192_
timestamp 1698175906
transform 1 0 10808 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _193_
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_
timestamp 1698175906
transform 1 0 13160 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1698175906
transform -1 0 7392 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _196_
timestamp 1698175906
transform 1 0 10360 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _197_
timestamp 1698175906
transform 1 0 12656 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _198_
timestamp 1698175906
transform 1 0 12768 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _199_
timestamp 1698175906
transform 1 0 7784 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _200_
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1698175906
transform 1 0 9408 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_
timestamp 1698175906
transform 1 0 8344 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform 1 0 10192 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform 1 0 13160 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform 1 0 12208 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform -1 0 7280 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform 1 0 7672 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform 1 0 7448 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform 1 0 11816 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 12208 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform -1 0 7056 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _212_
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _213_
timestamp 1698175906
transform 1 0 13832 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _214_
timestamp 1698175906
transform 1 0 11816 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _215_
timestamp 1698175906
transform 1 0 9408 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _216_
timestamp 1698175906
transform 1 0 14280 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _217_
timestamp 1698175906
transform 1 0 14840 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8120 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__CLK
timestamp 1698175906
transform -1 0 11648 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__CLK
timestamp 1698175906
transform 1 0 8176 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__CLK
timestamp 1698175906
transform 1 0 7616 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__CLK
timestamp 1698175906
transform 1 0 12936 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__CLK
timestamp 1698175906
transform 1 0 12208 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__CLK
timestamp 1698175906
transform 1 0 13048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1698175906
transform 1 0 7504 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__CLK
timestamp 1698175906
transform 1 0 12320 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__CLK
timestamp 1698175906
transform 1 0 12544 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__CLK
timestamp 1698175906
transform 1 0 9856 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__CLK
timestamp 1698175906
transform 1 0 8400 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__CLK
timestamp 1698175906
transform 1 0 11144 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK
timestamp 1698175906
transform 1 0 10080 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1698175906
transform 1 0 12264 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform 1 0 13048 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 12096 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 7616 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform -1 0 9520 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 9240 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 11312 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 12096 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform -1 0 7168 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 9184 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9632 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform 1 0 9520 0 -1 8624
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 9632 0 -1 12544
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10416 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698175906
transform 1 0 11928 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698175906
transform 1 0 12040 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698175906
transform 1 0 9072 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_154
timestamp 1698175906
transform 1 0 9296 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_156
timestamp 1698175906
transform 1 0 9408 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_183 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10920 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_199
timestamp 1698175906
transform 1 0 11816 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 12264 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_220
timestamp 1698175906
transform 1 0 12992 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_222
timestamp 1698175906
transform 1 0 13104 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_249
timestamp 1698175906
transform 1 0 14616 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_265
timestamp 1698175906
transform 1 0 15512 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_273
timestamp 1698175906
transform 1 0 15960 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_277
timestamp 1698175906
transform 1 0 16184 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698175906
transform 1 0 16296 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_123
timestamp 1698175906
transform 1 0 7560 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_154
timestamp 1698175906
transform 1 0 9296 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_158
timestamp 1698175906
transform 1 0 9520 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 10416 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_144
timestamp 1698175906
transform 1 0 8736 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_151
timestamp 1698175906
transform 1 0 9128 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_155
timestamp 1698175906
transform 1 0 9352 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_185
timestamp 1698175906
transform 1 0 11032 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_189
timestamp 1698175906
transform 1 0 11256 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_197
timestamp 1698175906
transform 1 0 11704 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_201
timestamp 1698175906
transform 1 0 11928 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_203
timestamp 1698175906
transform 1 0 12040 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698175906
transform 1 0 12208 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_115
timestamp 1698175906
transform 1 0 7112 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_119
timestamp 1698175906
transform 1 0 7336 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_167
timestamp 1698175906
transform 1 0 10024 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_235
timestamp 1698175906
transform 1 0 13832 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698175906
transform 1 0 14280 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 8288 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_146
timestamp 1698175906
transform 1 0 8848 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_155
timestamp 1698175906
transform 1 0 9352 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_159
timestamp 1698175906
transform 1 0 9576 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_161
timestamp 1698175906
transform 1 0 9688 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_170
timestamp 1698175906
transform 1 0 10192 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_187
timestamp 1698175906
transform 1 0 11144 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_195
timestamp 1698175906
transform 1 0 11592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_197
timestamp 1698175906
transform 1 0 11704 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_204
timestamp 1698175906
transform 1 0 12096 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698175906
transform 1 0 12320 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_225
timestamp 1698175906
transform 1 0 13272 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_257
timestamp 1698175906
transform 1 0 15064 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_273
timestamp 1698175906
transform 1 0 15960 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698175906
transform 1 0 16184 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 16296 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_136
timestamp 1698175906
transform 1 0 8288 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_140
timestamp 1698175906
transform 1 0 8512 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_156
timestamp 1698175906
transform 1 0 9408 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_163
timestamp 1698175906
transform 1 0 9800 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698175906
transform 1 0 10248 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_183
timestamp 1698175906
transform 1 0 10920 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_191
timestamp 1698175906
transform 1 0 11368 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_193
timestamp 1698175906
transform 1 0 11480 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_206
timestamp 1698175906
transform 1 0 12208 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_238
timestamp 1698175906
transform 1 0 14000 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698175906
transform 1 0 14224 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 14336 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_88
timestamp 1698175906
transform 1 0 5600 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_92
timestamp 1698175906
transform 1 0 5824 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_122
timestamp 1698175906
transform 1 0 7504 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_134
timestamp 1698175906
transform 1 0 8176 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698175906
transform 1 0 8400 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698175906
transform 1 0 12320 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_216
timestamp 1698175906
transform 1 0 12768 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_218
timestamp 1698175906
transform 1 0 12880 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_231
timestamp 1698175906
transform 1 0 13608 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_263
timestamp 1698175906
transform 1 0 15400 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 16296 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 20048 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 20160 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_115
timestamp 1698175906
transform 1 0 7112 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_134
timestamp 1698175906
transform 1 0 8176 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_142
timestamp 1698175906
transform 1 0 8624 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_144
timestamp 1698175906
transform 1 0 8736 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_151
timestamp 1698175906
transform 1 0 9128 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_155
timestamp 1698175906
transform 1 0 9352 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_163
timestamp 1698175906
transform 1 0 9800 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698175906
transform 1 0 10304 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 10416 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_183
timestamp 1698175906
transform 1 0 10920 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_197
timestamp 1698175906
transform 1 0 11704 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_251
timestamp 1698175906
transform 1 0 14728 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_104
timestamp 1698175906
transform 1 0 6496 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_112
timestamp 1698175906
transform 1 0 6944 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_116
timestamp 1698175906
transform 1 0 7168 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_118
timestamp 1698175906
transform 1 0 7280 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_125
timestamp 1698175906
transform 1 0 7672 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_133
timestamp 1698175906
transform 1 0 8120 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_146
timestamp 1698175906
transform 1 0 8848 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_161
timestamp 1698175906
transform 1 0 9688 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_173
timestamp 1698175906
transform 1 0 10360 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_175
timestamp 1698175906
transform 1 0 10472 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_196
timestamp 1698175906
transform 1 0 11648 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_198
timestamp 1698175906
transform 1 0 11760 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 12376 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_218
timestamp 1698175906
transform 1 0 12880 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_220
timestamp 1698175906
transform 1 0 12992 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_252
timestamp 1698175906
transform 1 0 14784 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_268
timestamp 1698175906
transform 1 0 15680 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698175906
transform 1 0 16128 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 20048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 20160 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_69
timestamp 1698175906
transform 1 0 4536 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_85
timestamp 1698175906
transform 1 0 5432 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_93
timestamp 1698175906
transform 1 0 5880 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_97
timestamp 1698175906
transform 1 0 6104 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_103
timestamp 1698175906
transform 1 0 6440 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_111
timestamp 1698175906
transform 1 0 6888 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_123
timestamp 1698175906
transform 1 0 7560 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_131
timestamp 1698175906
transform 1 0 8008 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_135
timestamp 1698175906
transform 1 0 8232 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_147
timestamp 1698175906
transform 1 0 8904 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_159
timestamp 1698175906
transform 1 0 9576 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698175906
transform 1 0 10360 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_177
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_210
timestamp 1698175906
transform 1 0 12432 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_212
timestamp 1698175906
transform 1 0 12544 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_231
timestamp 1698175906
transform 1 0 13608 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_239
timestamp 1698175906
transform 1 0 14056 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 14336 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 2240 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 4032 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 4480 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_80
timestamp 1698175906
transform 1 0 5152 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_84
timestamp 1698175906
transform 1 0 5376 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_114
timestamp 1698175906
transform 1 0 7056 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_116
timestamp 1698175906
transform 1 0 7168 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_129
timestamp 1698175906
transform 1 0 7896 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 8456 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_150
timestamp 1698175906
transform 1 0 9072 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_217
timestamp 1698175906
transform 1 0 12824 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_221
timestamp 1698175906
transform 1 0 13048 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_253
timestamp 1698175906
transform 1 0 14840 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_269
timestamp 1698175906
transform 1 0 15736 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698175906
transform 1 0 16184 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 16296 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 20048 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 20160 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_111
timestamp 1698175906
transform 1 0 6888 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_113
timestamp 1698175906
transform 1 0 7000 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_116
timestamp 1698175906
transform 1 0 7168 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_148
timestamp 1698175906
transform 1 0 8960 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_164
timestamp 1698175906
transform 1 0 9856 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_172
timestamp 1698175906
transform 1 0 10304 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698175906
transform 1 0 10416 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_183
timestamp 1698175906
transform 1 0 10920 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_185
timestamp 1698175906
transform 1 0 11032 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_192
timestamp 1698175906
transform 1 0 11424 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_224
timestamp 1698175906
transform 1 0 13216 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_240
timestamp 1698175906
transform 1 0 14112 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 14336 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 18648 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_88
timestamp 1698175906
transform 1 0 5600 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_125
timestamp 1698175906
transform 1 0 7672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_127
timestamp 1698175906
transform 1 0 7784 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_132
timestamp 1698175906
transform 1 0 8064 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698175906
transform 1 0 8288 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_152
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_160
timestamp 1698175906
transform 1 0 9632 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_164
timestamp 1698175906
transform 1 0 9856 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_170
timestamp 1698175906
transform 1 0 10192 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_186
timestamp 1698175906
transform 1 0 11088 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_219
timestamp 1698175906
transform 1 0 12936 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_252
timestamp 1698175906
transform 1 0 14784 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_268
timestamp 1698175906
transform 1 0 15680 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698175906
transform 1 0 16128 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_115
timestamp 1698175906
transform 1 0 7112 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_122
timestamp 1698175906
transform 1 0 7504 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_126
timestamp 1698175906
transform 1 0 7728 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_134
timestamp 1698175906
transform 1 0 8176 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_152
timestamp 1698175906
transform 1 0 9184 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_156
timestamp 1698175906
transform 1 0 9408 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_165
timestamp 1698175906
transform 1 0 9912 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_177
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_197
timestamp 1698175906
transform 1 0 11704 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_240
timestamp 1698175906
transform 1 0 14112 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 14336 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_259
timestamp 1698175906
transform 1 0 15176 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_291
timestamp 1698175906
transform 1 0 16968 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_307
timestamp 1698175906
transform 1 0 17864 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 2240 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 4032 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 4480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_88
timestamp 1698175906
transform 1 0 5600 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_118
timestamp 1698175906
transform 1 0 7280 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_120
timestamp 1698175906
transform 1 0 7392 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_129
timestamp 1698175906
transform 1 0 7896 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698175906
transform 1 0 8344 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 8456 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_144
timestamp 1698175906
transform 1 0 8736 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_163
timestamp 1698175906
transform 1 0 9800 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_167
timestamp 1698175906
transform 1 0 10024 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_169
timestamp 1698175906
transform 1 0 10136 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_205
timestamp 1698175906
transform 1 0 12152 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698175906
transform 1 0 16128 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_115
timestamp 1698175906
transform 1 0 7112 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_130
timestamp 1698175906
transform 1 0 7952 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_138
timestamp 1698175906
transform 1 0 8400 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_148
timestamp 1698175906
transform 1 0 8960 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_164
timestamp 1698175906
transform 1 0 9856 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698175906
transform 1 0 10304 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 10416 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698175906
transform 1 0 14168 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 2240 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 4032 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 4480 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_88
timestamp 1698175906
transform 1 0 5600 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_92
timestamp 1698175906
transform 1 0 5824 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_131
timestamp 1698175906
transform 1 0 8008 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_135
timestamp 1698175906
transform 1 0 8232 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 8456 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_155
timestamp 1698175906
transform 1 0 9352 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_159
timestamp 1698175906
transform 1 0 9576 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_233
timestamp 1698175906
transform 1 0 13720 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_265
timestamp 1698175906
transform 1 0 15512 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_273
timestamp 1698175906
transform 1 0 15960 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698175906
transform 1 0 16184 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 16296 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 18256 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 18704 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 2240 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 2464 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_115
timestamp 1698175906
transform 1 0 7112 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_119
timestamp 1698175906
transform 1 0 7336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_125
timestamp 1698175906
transform 1 0 7672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_162
timestamp 1698175906
transform 1 0 9744 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_166
timestamp 1698175906
transform 1 0 9968 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 10416 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_177
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_181
timestamp 1698175906
transform 1 0 10808 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_191
timestamp 1698175906
transform 1 0 11368 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_197
timestamp 1698175906
transform 1 0 11704 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_199
timestamp 1698175906
transform 1 0 11816 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698175906
transform 1 0 14168 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 18648 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_88
timestamp 1698175906
transform 1 0 5600 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_90
timestamp 1698175906
transform 1 0 5712 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_120
timestamp 1698175906
transform 1 0 7392 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_124
timestamp 1698175906
transform 1 0 7616 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_157
timestamp 1698175906
transform 1 0 9464 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_159
timestamp 1698175906
transform 1 0 9576 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_165
timestamp 1698175906
transform 1 0 9912 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_202
timestamp 1698175906
transform 1 0 11984 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_206
timestamp 1698175906
transform 1 0 12208 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_249
timestamp 1698175906
transform 1 0 14616 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_265
timestamp 1698175906
transform 1 0 15512 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_273
timestamp 1698175906
transform 1 0 15960 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 16184 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 16296 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_123
timestamp 1698175906
transform 1 0 7560 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_131
timestamp 1698175906
transform 1 0 8008 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_135
timestamp 1698175906
transform 1 0 8232 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_166
timestamp 1698175906
transform 1 0 9968 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_170
timestamp 1698175906
transform 1 0 10192 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698175906
transform 1 0 10416 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_190
timestamp 1698175906
transform 1 0 11312 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_206
timestamp 1698175906
transform 1 0 12208 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_210
timestamp 1698175906
transform 1 0 12432 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_214
timestamp 1698175906
transform 1 0 12656 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_227
timestamp 1698175906
transform 1 0 13384 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698175906
transform 1 0 14280 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 18648 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_158
timestamp 1698175906
transform 1 0 9520 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_162
timestamp 1698175906
transform 1 0 9744 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_192
timestamp 1698175906
transform 1 0 11424 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_196
timestamp 1698175906
transform 1 0 11648 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_204
timestamp 1698175906
transform 1 0 12096 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698175906
transform 1 0 12320 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_314
timestamp 1698175906
transform 1 0 18256 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_322
timestamp 1698175906
transform 1 0 18704 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_139
timestamp 1698175906
transform 1 0 8456 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_147
timestamp 1698175906
transform 1 0 8904 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_158
timestamp 1698175906
transform 1 0 9520 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_162
timestamp 1698175906
transform 1 0 9744 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_189
timestamp 1698175906
transform 1 0 11256 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_205
timestamp 1698175906
transform 1 0 12152 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 16128 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18760 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 13160 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 10472 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 9800 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 18760 0 -1 14112
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 18760 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18760 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform -1 0 10192 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 9016 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 8736 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 2240 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 9464 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 18760 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 18760 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 12096 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform -1 0 2240 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform -1 0 2240 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698175906
transform -1 0 2240 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13440 400 13496 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 20600 10416 21000 10472 0 FreeSans 224 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 13104 0 13160 400 0 FreeSans 224 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 0 8400 400 8456 0 FreeSans 224 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 10416 0 10472 400 0 FreeSans 224 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 9744 20600 9800 21000 0 FreeSans 224 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 20600 13440 21000 13496 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 20600 12096 21000 12152 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 9408 20600 9464 21000 0 FreeSans 224 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 9072 20600 9128 21000 0 FreeSans 224 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 11424 400 11480 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 9408 0 9464 400 0 FreeSans 224 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 11760 20600 11816 21000 0 FreeSans 224 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 20600 10752 21000 10808 0 FreeSans 224 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 20600 9408 21000 9464 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 20600 12432 21000 12488 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 9744 400 9800 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 0 12096 400 12152 0 FreeSans 224 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 0 12432 400 12488 0 FreeSans 224 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 8260 12936 8260 12936 0 _000_
rlabel metal2 7224 8092 7224 8092 0 _001_
rlabel metal2 9856 6916 9856 6916 0 _002_
rlabel metal2 8820 13356 8820 13356 0 _003_
rlabel metal3 10836 11228 10836 11228 0 _004_
rlabel metal2 13636 10948 13636 10948 0 _005_
rlabel metal2 12684 12572 12684 12572 0 _006_
rlabel metal3 7196 11508 7196 11508 0 _007_
rlabel metal2 8148 6636 8148 6636 0 _008_
rlabel metal2 9268 7280 9268 7280 0 _009_
rlabel metal2 12152 10724 12152 10724 0 _010_
rlabel metal2 12684 7448 12684 7448 0 _011_
rlabel metal2 6356 9828 6356 9828 0 _012_
rlabel metal2 7756 12068 7756 12068 0 _013_
rlabel metal2 10724 13720 10724 13720 0 _014_
rlabel metal3 7224 10836 7224 10836 0 _015_
rlabel metal2 7420 8876 7420 8876 0 _016_
rlabel metal2 11172 9436 11172 9436 0 _017_
rlabel metal2 11060 7504 11060 7504 0 _018_
rlabel metal2 13524 9212 13524 9212 0 _019_
rlabel metal2 7700 12516 7700 12516 0 _020_
rlabel metal2 11060 12908 11060 12908 0 _021_
rlabel metal2 13132 12768 13132 12768 0 _022_
rlabel metal2 13412 8652 13412 8652 0 _023_
rlabel metal2 13468 8624 13468 8624 0 _024_
rlabel metal2 11620 10430 11620 10430 0 _025_
rlabel metal2 8960 12348 8960 12348 0 _026_
rlabel metal2 8988 12796 8988 12796 0 _027_
rlabel metal2 8484 10598 8484 10598 0 _028_
rlabel metal2 8652 12796 8652 12796 0 _029_
rlabel metal2 11368 10612 11368 10612 0 _030_
rlabel metal2 8036 8960 8036 8960 0 _031_
rlabel metal2 7868 8624 7868 8624 0 _032_
rlabel metal2 7588 8848 7588 8848 0 _033_
rlabel metal2 10668 7840 10668 7840 0 _034_
rlabel metal2 9800 7756 9800 7756 0 _035_
rlabel metal2 10500 8204 10500 8204 0 _036_
rlabel metal2 10164 7700 10164 7700 0 _037_
rlabel metal2 9772 13076 9772 13076 0 _038_
rlabel metal2 11172 11256 11172 11256 0 _039_
rlabel metal2 11900 10780 11900 10780 0 _040_
rlabel metal2 11564 11004 11564 11004 0 _041_
rlabel metal2 13692 11200 13692 11200 0 _042_
rlabel metal2 12964 12376 12964 12376 0 _043_
rlabel metal2 12124 11060 12124 11060 0 _044_
rlabel metal2 7476 11368 7476 11368 0 _045_
rlabel metal2 9044 7028 9044 7028 0 _046_
rlabel metal2 9128 7252 9128 7252 0 _047_
rlabel metal2 9380 7588 9380 7588 0 _048_
rlabel metal3 12516 10780 12516 10780 0 _049_
rlabel metal2 12628 7840 12628 7840 0 _050_
rlabel metal2 12992 7700 12992 7700 0 _051_
rlabel metal3 6720 9548 6720 9548 0 _052_
rlabel metal2 11564 9016 11564 9016 0 _053_
rlabel metal2 10164 9436 10164 9436 0 _054_
rlabel metal2 7308 11508 7308 11508 0 _055_
rlabel metal2 7672 11956 7672 11956 0 _056_
rlabel metal3 9492 11620 9492 11620 0 _057_
rlabel metal2 11900 9296 11900 9296 0 _058_
rlabel metal2 10332 11200 10332 11200 0 _059_
rlabel metal3 10388 11060 10388 11060 0 _060_
rlabel metal3 8372 11284 8372 11284 0 _061_
rlabel metal2 12012 8988 12012 8988 0 _062_
rlabel metal3 10444 9492 10444 9492 0 _063_
rlabel metal2 8792 11844 8792 11844 0 _064_
rlabel metal2 8960 9212 8960 9212 0 _065_
rlabel metal2 9688 11060 9688 11060 0 _066_
rlabel metal2 11060 11032 11060 11032 0 _067_
rlabel metal3 10444 9716 10444 9716 0 _068_
rlabel metal2 10948 11200 10948 11200 0 _069_
rlabel metal2 13524 12516 13524 12516 0 _070_
rlabel metal2 11228 13440 11228 13440 0 _071_
rlabel metal2 11004 13524 11004 13524 0 _072_
rlabel metal2 7616 9268 7616 9268 0 _073_
rlabel metal3 9184 9996 9184 9996 0 _074_
rlabel metal2 11508 10472 11508 10472 0 _075_
rlabel metal3 12712 8708 12712 8708 0 _076_
rlabel metal3 12040 12460 12040 12460 0 _077_
rlabel metal3 10514 9212 10514 9212 0 _078_
rlabel metal2 8820 10836 8820 10836 0 _079_
rlabel metal3 8848 9604 8848 9604 0 _080_
rlabel metal3 8288 9716 8288 9716 0 _081_
rlabel metal2 10108 9352 10108 9352 0 _082_
rlabel metal2 10892 8036 10892 8036 0 _083_
rlabel metal2 12740 7812 12740 7812 0 _084_
rlabel metal2 11788 8288 11788 8288 0 _085_
rlabel metal3 12264 8036 12264 8036 0 _086_
rlabel metal2 13356 9688 13356 9688 0 _087_
rlabel metal2 13832 9492 13832 9492 0 _088_
rlabel metal2 8708 12376 8708 12376 0 _089_
rlabel metal2 7476 12124 7476 12124 0 _090_
rlabel metal2 11396 12740 11396 12740 0 _091_
rlabel metal3 12908 12348 12908 12348 0 _092_
rlabel metal2 13356 12880 13356 12880 0 _093_
rlabel metal3 1239 13468 1239 13468 0 clk
rlabel metal2 9800 10836 9800 10836 0 clknet_0_clk
rlabel metal2 10668 7112 10668 7112 0 clknet_1_0__leaf_clk
rlabel metal2 13160 10780 13160 10780 0 clknet_1_1__leaf_clk
rlabel metal3 8344 10780 8344 10780 0 dut16.count\[0\]
rlabel metal2 7420 9716 7420 9716 0 dut16.count\[1\]
rlabel metal2 12740 9044 12740 9044 0 dut16.count\[2\]
rlabel metal2 12096 8092 12096 8092 0 dut16.count\[3\]
rlabel metal2 14756 10724 14756 10724 0 net1
rlabel metal2 11732 11536 11732 11536 0 net10
rlabel metal2 9632 12684 9632 12684 0 net11
rlabel metal2 9324 13104 9324 13104 0 net12
rlabel metal2 8904 7308 8904 7308 0 net13
rlabel metal2 13356 11088 13356 11088 0 net14
rlabel metal3 14476 8876 14476 8876 0 net15
rlabel metal3 3178 11564 3178 11564 0 net16
rlabel metal3 9380 6524 9380 6524 0 net17
rlabel metal3 15246 13188 15246 13188 0 net18
rlabel metal2 11872 13076 11872 13076 0 net19
rlabel metal2 13244 3178 13244 3178 0 net2
rlabel metal2 15092 10920 15092 10920 0 net20
rlabel metal2 14700 9380 14700 9380 0 net21
rlabel metal2 13748 12768 13748 12768 0 net22
rlabel metal2 11340 14056 11340 14056 0 net23
rlabel metal2 5516 9884 5516 9884 0 net24
rlabel metal2 6020 12320 6020 12320 0 net25
rlabel metal2 2156 12908 2156 12908 0 net26
rlabel metal3 3178 8820 3178 8820 0 net3
rlabel metal2 10948 6776 10948 6776 0 net4
rlabel metal2 9856 13580 9856 13580 0 net5
rlabel metal2 18956 13272 18956 13272 0 net6
rlabel metal2 18956 11984 18956 11984 0 net7
rlabel metal2 14980 11116 14980 11116 0 net8
rlabel metal2 14196 13104 14196 13104 0 net9
rlabel metal3 20321 10444 20321 10444 0 segm[0]
rlabel metal2 13132 1211 13132 1211 0 segm[10]
rlabel metal3 679 8428 679 8428 0 segm[11]
rlabel metal2 10444 1099 10444 1099 0 segm[12]
rlabel metal2 10388 19012 10388 19012 0 segm[13]
rlabel metal2 19964 13664 19964 13664 0 segm[1]
rlabel metal2 20020 12180 20020 12180 0 segm[2]
rlabel metal3 20321 11452 20321 11452 0 segm[3]
rlabel metal2 19964 12936 19964 12936 0 segm[4]
rlabel metal2 20020 11900 20020 11900 0 segm[5]
rlabel metal2 9436 19845 9436 19845 0 segm[6]
rlabel metal3 9352 18340 9352 18340 0 segm[7]
rlabel metal2 9100 1099 9100 1099 0 segm[8]
rlabel metal2 20020 11172 20020 11172 0 segm[9]
rlabel metal2 20020 8820 20020 8820 0 sel[0]
rlabel metal3 679 11452 679 11452 0 sel[10]
rlabel metal2 9436 1211 9436 1211 0 sel[11]
rlabel metal2 20020 13356 20020 13356 0 sel[1]
rlabel metal2 11788 19873 11788 19873 0 sel[2]
rlabel metal2 20020 10752 20020 10752 0 sel[3]
rlabel metal2 20020 9548 20020 9548 0 sel[4]
rlabel metal2 20020 12628 20020 12628 0 sel[5]
rlabel metal2 11116 19845 11116 19845 0 sel[6]
rlabel metal3 679 9772 679 9772 0 sel[7]
rlabel metal3 679 12124 679 12124 0 sel[8]
rlabel metal3 679 12460 679 12460 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
