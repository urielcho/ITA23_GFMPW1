magic
tech gf180mcuD
magscale 1 5
timestamp 1699642795
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 11215 19137 11241 19143
rect 11215 19105 11241 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 10705 18999 10711 19025
rect 10737 18999 10743 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 11383 18745 11409 18751
rect 11383 18713 11409 18719
rect 13119 18745 13145 18751
rect 13119 18713 13145 18719
rect 11097 18607 11103 18633
rect 11129 18607 11135 18633
rect 12609 18607 12615 18633
rect 12641 18607 12647 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 855 18185 881 18191
rect 855 18153 881 18159
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 10767 14041 10793 14047
rect 10767 14009 10793 14015
rect 10823 13929 10849 13935
rect 10823 13897 10849 13903
rect 10767 13817 10793 13823
rect 10767 13785 10793 13791
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 10935 13537 10961 13543
rect 10935 13505 10961 13511
rect 11103 13537 11129 13543
rect 11103 13505 11129 13511
rect 10761 13455 10767 13481
rect 10793 13455 10799 13481
rect 11265 13455 11271 13481
rect 11297 13455 11303 13481
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 10873 13231 10879 13257
rect 10905 13231 10911 13257
rect 11943 13201 11969 13207
rect 11943 13169 11969 13175
rect 11999 13201 12025 13207
rect 11999 13169 12025 13175
rect 13287 13201 13313 13207
rect 13287 13169 13313 13175
rect 13343 13201 13369 13207
rect 13343 13169 13369 13175
rect 11831 13145 11857 13151
rect 9361 13119 9367 13145
rect 9393 13119 9399 13145
rect 11831 13113 11857 13119
rect 13175 13145 13201 13151
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 13175 13113 13201 13119
rect 9753 13063 9759 13089
rect 9785 13063 9791 13089
rect 19945 13063 19951 13089
rect 19977 13063 19983 13089
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 967 12809 993 12815
rect 20007 12809 20033 12815
rect 9585 12783 9591 12809
rect 9617 12783 9623 12809
rect 12385 12783 12391 12809
rect 12417 12783 12423 12809
rect 14009 12783 14015 12809
rect 14041 12783 14047 12809
rect 967 12777 993 12783
rect 20007 12777 20033 12783
rect 9759 12753 9785 12759
rect 2137 12727 2143 12753
rect 2169 12727 2175 12753
rect 8129 12727 8135 12753
rect 8161 12727 8167 12753
rect 9759 12721 9785 12727
rect 9927 12753 9953 12759
rect 10929 12727 10935 12753
rect 10961 12727 10967 12753
rect 12609 12727 12615 12753
rect 12641 12727 12647 12753
rect 18825 12727 18831 12753
rect 18857 12727 18863 12753
rect 9927 12721 9953 12727
rect 8521 12671 8527 12697
rect 8553 12671 8559 12697
rect 11321 12671 11327 12697
rect 11353 12671 11359 12697
rect 12945 12671 12951 12697
rect 12977 12671 12983 12697
rect 9871 12641 9897 12647
rect 9871 12609 9897 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 9647 12473 9673 12479
rect 9647 12441 9673 12447
rect 11439 12473 11465 12479
rect 11825 12447 11831 12473
rect 11857 12447 11863 12473
rect 11439 12441 11465 12447
rect 8359 12417 8385 12423
rect 9759 12417 9785 12423
rect 9361 12391 9367 12417
rect 9393 12391 9399 12417
rect 8359 12385 8385 12391
rect 9759 12385 9785 12391
rect 8247 12361 8273 12367
rect 8073 12335 8079 12361
rect 8105 12335 8111 12361
rect 8247 12329 8273 12335
rect 8415 12361 8441 12367
rect 9815 12361 9841 12367
rect 9473 12335 9479 12361
rect 9505 12335 9511 12361
rect 8415 12329 8441 12335
rect 9815 12329 9841 12335
rect 11383 12361 11409 12367
rect 11383 12329 11409 12335
rect 11495 12361 11521 12367
rect 11495 12329 11521 12335
rect 11719 12361 11745 12367
rect 11937 12335 11943 12361
rect 11969 12335 11975 12361
rect 12665 12335 12671 12361
rect 12697 12335 12703 12361
rect 11719 12329 11745 12335
rect 6673 12279 6679 12305
rect 6705 12279 6711 12305
rect 7737 12279 7743 12305
rect 7769 12279 7775 12305
rect 13001 12279 13007 12305
rect 13033 12279 13039 12305
rect 14065 12279 14071 12305
rect 14097 12279 14103 12305
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 9087 12081 9113 12087
rect 9087 12049 9113 12055
rect 9591 12081 9617 12087
rect 9591 12049 9617 12055
rect 13735 12081 13761 12087
rect 13735 12049 13761 12055
rect 7743 12025 7769 12031
rect 7743 11993 7769 11999
rect 12839 12025 12865 12031
rect 12839 11993 12865 11999
rect 13287 12025 13313 12031
rect 13287 11993 13313 11999
rect 20007 12025 20033 12031
rect 20007 11993 20033 11999
rect 7687 11969 7713 11975
rect 7687 11937 7713 11943
rect 7855 11969 7881 11975
rect 7855 11937 7881 11943
rect 9423 11969 9449 11975
rect 9423 11937 9449 11943
rect 13119 11969 13145 11975
rect 13119 11937 13145 11943
rect 13567 11969 13593 11975
rect 13567 11937 13593 11943
rect 13679 11969 13705 11975
rect 18825 11943 18831 11969
rect 18857 11943 18863 11969
rect 13679 11937 13705 11943
rect 7519 11913 7545 11919
rect 7519 11881 7545 11887
rect 9143 11913 9169 11919
rect 9143 11881 9169 11887
rect 9311 11913 9337 11919
rect 9311 11881 9337 11887
rect 13231 11913 13257 11919
rect 13231 11881 13257 11887
rect 13343 11913 13369 11919
rect 13343 11881 13369 11887
rect 13735 11913 13761 11919
rect 13735 11881 13761 11887
rect 9087 11857 9113 11863
rect 9087 11825 9113 11831
rect 9759 11857 9785 11863
rect 12783 11857 12809 11863
rect 9921 11831 9927 11857
rect 9953 11831 9959 11857
rect 9759 11825 9785 11831
rect 12783 11825 12809 11831
rect 12895 11857 12921 11863
rect 12895 11825 12921 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 8241 11663 8247 11689
rect 8273 11663 8279 11689
rect 9087 11633 9113 11639
rect 9087 11601 9113 11607
rect 11887 11633 11913 11639
rect 11887 11601 11913 11607
rect 11943 11633 11969 11639
rect 11943 11601 11969 11607
rect 11775 11577 11801 11583
rect 8129 11551 8135 11577
rect 8161 11551 8167 11577
rect 9305 11551 9311 11577
rect 9337 11551 9343 11577
rect 18825 11551 18831 11577
rect 18857 11551 18863 11577
rect 11775 11545 11801 11551
rect 9697 11495 9703 11521
rect 9729 11495 9735 11521
rect 10761 11495 10767 11521
rect 10793 11495 10799 11521
rect 9143 11465 9169 11471
rect 9143 11433 9169 11439
rect 20007 11465 20033 11471
rect 20007 11433 20033 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 9479 11297 9505 11303
rect 9479 11265 9505 11271
rect 10319 11297 10345 11303
rect 10319 11265 10345 11271
rect 967 11241 993 11247
rect 7239 11241 7265 11247
rect 7065 11215 7071 11241
rect 7097 11215 7103 11241
rect 967 11209 993 11215
rect 7239 11209 7265 11215
rect 7463 11241 7489 11247
rect 7463 11209 7489 11215
rect 8751 11241 8777 11247
rect 8751 11209 8777 11215
rect 9871 11241 9897 11247
rect 20007 11241 20033 11247
rect 12329 11215 12335 11241
rect 12361 11215 12367 11241
rect 9871 11209 9897 11215
rect 20007 11209 20033 11215
rect 7631 11185 7657 11191
rect 9311 11185 9337 11191
rect 2137 11159 2143 11185
rect 2169 11159 2175 11185
rect 7513 11159 7519 11185
rect 7545 11159 7551 11185
rect 7793 11159 7799 11185
rect 7825 11159 7831 11185
rect 7631 11153 7657 11159
rect 9311 11153 9337 11159
rect 9815 11185 9841 11191
rect 9815 11153 9841 11159
rect 10151 11185 10177 11191
rect 13231 11185 13257 11191
rect 10929 11159 10935 11185
rect 10961 11159 10967 11185
rect 18937 11159 18943 11185
rect 18969 11159 18975 11185
rect 10151 11153 10177 11159
rect 13231 11153 13257 11159
rect 7407 11129 7433 11135
rect 7407 11097 7433 11103
rect 9031 11129 9057 11135
rect 9031 11097 9057 11103
rect 9199 11129 9225 11135
rect 9199 11097 9225 11103
rect 10263 11129 10289 11135
rect 11265 11103 11271 11129
rect 11297 11103 11303 11129
rect 10263 11097 10289 11103
rect 7127 11073 7153 11079
rect 7127 11041 7153 11047
rect 8863 11073 8889 11079
rect 8863 11041 8889 11047
rect 8975 11073 9001 11079
rect 8975 11041 9001 11047
rect 9927 11073 9953 11079
rect 9927 11041 9953 11047
rect 10319 11073 10345 11079
rect 10319 11041 10345 11047
rect 13119 11073 13145 11079
rect 13119 11041 13145 11047
rect 13175 11073 13201 11079
rect 13175 11041 13201 11047
rect 13343 11073 13369 11079
rect 13343 11041 13369 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 7799 10905 7825 10911
rect 7799 10873 7825 10879
rect 8191 10905 8217 10911
rect 8191 10873 8217 10879
rect 9087 10905 9113 10911
rect 9087 10873 9113 10879
rect 12615 10905 12641 10911
rect 12615 10873 12641 10879
rect 7743 10849 7769 10855
rect 7009 10823 7015 10849
rect 7041 10823 7047 10849
rect 7743 10817 7769 10823
rect 7855 10849 7881 10855
rect 7855 10817 7881 10823
rect 8303 10849 8329 10855
rect 9199 10849 9225 10855
rect 8913 10823 8919 10849
rect 8945 10823 8951 10849
rect 13449 10823 13455 10849
rect 13481 10823 13487 10849
rect 14849 10823 14855 10849
rect 14881 10823 14887 10849
rect 15185 10823 15191 10849
rect 15217 10823 15223 10849
rect 8303 10817 8329 10823
rect 9199 10817 9225 10823
rect 8079 10793 8105 10799
rect 2137 10767 2143 10793
rect 2169 10767 2175 10793
rect 7401 10767 7407 10793
rect 7433 10767 7439 10793
rect 8079 10761 8105 10767
rect 8191 10793 8217 10799
rect 9143 10793 9169 10799
rect 8801 10767 8807 10793
rect 8833 10767 8839 10793
rect 8191 10761 8217 10767
rect 9143 10761 9169 10767
rect 9423 10793 9449 10799
rect 12727 10793 12753 10799
rect 9697 10767 9703 10793
rect 9729 10767 9735 10793
rect 9423 10761 9449 10767
rect 12727 10761 12753 10767
rect 12951 10793 12977 10799
rect 12951 10761 12977 10767
rect 13057 10761 13063 10787
rect 13089 10761 13095 10787
rect 14737 10767 14743 10793
rect 14769 10767 14775 10793
rect 15073 10767 15079 10793
rect 15105 10767 15111 10793
rect 18825 10767 18831 10793
rect 18857 10767 18863 10793
rect 967 10737 993 10743
rect 12671 10737 12697 10743
rect 20007 10737 20033 10743
rect 5945 10711 5951 10737
rect 5977 10711 5983 10737
rect 11657 10711 11663 10737
rect 11689 10711 11695 10737
rect 14513 10711 14519 10737
rect 14545 10711 14551 10737
rect 967 10705 993 10711
rect 12671 10705 12697 10711
rect 20007 10705 20033 10711
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 7351 10513 7377 10519
rect 7351 10481 7377 10487
rect 967 10457 993 10463
rect 7463 10457 7489 10463
rect 11271 10457 11297 10463
rect 4993 10431 4999 10457
rect 5025 10431 5031 10457
rect 7961 10431 7967 10457
rect 7993 10431 7999 10457
rect 967 10425 993 10431
rect 7463 10425 7489 10431
rect 11271 10425 11297 10431
rect 20007 10457 20033 10463
rect 20007 10425 20033 10431
rect 7575 10401 7601 10407
rect 10879 10401 10905 10407
rect 2137 10375 2143 10401
rect 2169 10375 2175 10401
rect 6449 10375 6455 10401
rect 6481 10375 6487 10401
rect 6841 10375 6847 10401
rect 6873 10375 6879 10401
rect 7121 10375 7127 10401
rect 7153 10375 7159 10401
rect 10033 10375 10039 10401
rect 10065 10375 10071 10401
rect 7575 10369 7601 10375
rect 10879 10369 10905 10375
rect 11215 10401 11241 10407
rect 11215 10369 11241 10375
rect 11551 10401 11577 10407
rect 11657 10375 11663 10401
rect 11689 10375 11695 10401
rect 14625 10375 14631 10401
rect 14657 10375 14663 10401
rect 14961 10375 14967 10401
rect 14993 10375 14999 10401
rect 18825 10375 18831 10401
rect 18857 10375 18863 10401
rect 11551 10369 11577 10375
rect 10711 10345 10737 10351
rect 6057 10319 6063 10345
rect 6089 10319 6095 10345
rect 6729 10319 6735 10345
rect 6761 10319 6767 10345
rect 7233 10319 7239 10345
rect 7265 10319 7271 10345
rect 12889 10319 12895 10345
rect 12921 10319 12927 10345
rect 10711 10313 10737 10319
rect 10655 10289 10681 10295
rect 11327 10289 11353 10295
rect 7289 10263 7295 10289
rect 7321 10263 7327 10289
rect 11041 10263 11047 10289
rect 11073 10263 11079 10289
rect 14737 10263 14743 10289
rect 14769 10263 14775 10289
rect 15073 10263 15079 10289
rect 15105 10263 15111 10289
rect 10655 10257 10681 10263
rect 11327 10257 11353 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 8359 10121 8385 10127
rect 8359 10089 8385 10095
rect 14519 10121 14545 10127
rect 14519 10089 14545 10095
rect 6735 10065 6761 10071
rect 6735 10033 6761 10039
rect 6791 10065 6817 10071
rect 6791 10033 6817 10039
rect 6847 10065 6873 10071
rect 6847 10033 6873 10039
rect 7351 10065 7377 10071
rect 10655 10065 10681 10071
rect 7737 10039 7743 10065
rect 7769 10039 7775 10065
rect 10481 10039 10487 10065
rect 10513 10039 10519 10065
rect 7351 10033 7377 10039
rect 10655 10033 10681 10039
rect 10711 10065 10737 10071
rect 10711 10033 10737 10039
rect 10823 10065 10849 10071
rect 11881 10039 11887 10065
rect 11913 10039 11919 10065
rect 10823 10033 10849 10039
rect 7239 10009 7265 10015
rect 8415 10009 8441 10015
rect 9479 10009 9505 10015
rect 10319 10009 10345 10015
rect 14463 10009 14489 10015
rect 2137 9983 2143 10009
rect 2169 9983 2175 10009
rect 7121 9983 7127 10009
rect 7153 9983 7159 10009
rect 7457 9983 7463 10009
rect 7489 9983 7495 10009
rect 7849 9983 7855 10009
rect 7881 9983 7887 10009
rect 8857 9983 8863 10009
rect 8889 9983 8895 10009
rect 9249 9983 9255 10009
rect 9281 9983 9287 10009
rect 9865 9983 9871 10009
rect 9897 9983 9903 10009
rect 9977 9983 9983 10009
rect 10009 9983 10015 10009
rect 11993 9983 11999 10009
rect 12025 9983 12031 10009
rect 12889 9983 12895 10009
rect 12921 9983 12927 10009
rect 18825 9983 18831 10009
rect 18857 9983 18863 10009
rect 7239 9977 7265 9983
rect 8415 9977 8441 9983
rect 9479 9977 9505 9983
rect 10319 9977 10345 9983
rect 14463 9977 14489 9983
rect 7295 9953 7321 9959
rect 20007 9953 20033 9959
rect 9081 9927 9087 9953
rect 9113 9927 9119 9953
rect 9641 9927 9647 9953
rect 9673 9927 9679 9953
rect 13225 9927 13231 9953
rect 13257 9927 13263 9953
rect 14289 9927 14295 9953
rect 14321 9927 14327 9953
rect 7295 9921 7321 9927
rect 20007 9921 20033 9927
rect 967 9897 993 9903
rect 14519 9897 14545 9903
rect 8857 9871 8863 9897
rect 8889 9871 8895 9897
rect 967 9865 993 9871
rect 14519 9865 14545 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 6735 9729 6761 9735
rect 6735 9697 6761 9703
rect 9311 9729 9337 9735
rect 9311 9697 9337 9703
rect 10263 9729 10289 9735
rect 10263 9697 10289 9703
rect 20007 9729 20033 9735
rect 20007 9697 20033 9703
rect 9697 9647 9703 9673
rect 9729 9647 9735 9673
rect 8639 9617 8665 9623
rect 6897 9591 6903 9617
rect 6929 9591 6935 9617
rect 8353 9591 8359 9617
rect 8385 9591 8391 9617
rect 8639 9585 8665 9591
rect 8695 9617 8721 9623
rect 8695 9585 8721 9591
rect 8919 9617 8945 9623
rect 8919 9585 8945 9591
rect 9087 9617 9113 9623
rect 9087 9585 9113 9591
rect 9423 9617 9449 9623
rect 10207 9617 10233 9623
rect 9865 9591 9871 9617
rect 9897 9591 9903 9617
rect 9423 9585 9449 9591
rect 10207 9585 10233 9591
rect 12223 9617 12249 9623
rect 12223 9585 12249 9591
rect 13623 9617 13649 9623
rect 13623 9585 13649 9591
rect 13791 9617 13817 9623
rect 18825 9591 18831 9617
rect 18857 9591 18863 9617
rect 13791 9585 13817 9591
rect 9031 9561 9057 9567
rect 8241 9535 8247 9561
rect 8273 9535 8279 9561
rect 9031 9529 9057 9535
rect 9199 9561 9225 9567
rect 9199 9529 9225 9535
rect 10151 9561 10177 9567
rect 10151 9529 10177 9535
rect 13735 9561 13761 9567
rect 13735 9529 13761 9535
rect 6791 9505 6817 9511
rect 6791 9473 6817 9479
rect 8751 9505 8777 9511
rect 12385 9479 12391 9505
rect 12417 9479 12423 9505
rect 8751 9473 8777 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 9927 9337 9953 9343
rect 9927 9305 9953 9311
rect 11103 9337 11129 9343
rect 11103 9305 11129 9311
rect 12055 9337 12081 9343
rect 12055 9305 12081 9311
rect 12783 9337 12809 9343
rect 12783 9305 12809 9311
rect 13119 9337 13145 9343
rect 13119 9305 13145 9311
rect 13231 9337 13257 9343
rect 13231 9305 13257 9311
rect 7295 9281 7321 9287
rect 7295 9249 7321 9255
rect 7351 9281 7377 9287
rect 7351 9249 7377 9255
rect 9479 9281 9505 9287
rect 9479 9249 9505 9255
rect 10039 9281 10065 9287
rect 10039 9249 10065 9255
rect 10095 9281 10121 9287
rect 10095 9249 10121 9255
rect 11719 9281 11745 9287
rect 11719 9249 11745 9255
rect 11775 9281 11801 9287
rect 11775 9249 11801 9255
rect 11887 9281 11913 9287
rect 11887 9249 11913 9255
rect 12671 9281 12697 9287
rect 12671 9249 12697 9255
rect 13623 9281 13649 9287
rect 13623 9249 13649 9255
rect 13679 9281 13705 9287
rect 13679 9249 13705 9255
rect 13903 9281 13929 9287
rect 13903 9249 13929 9255
rect 13959 9281 13985 9287
rect 13959 9249 13985 9255
rect 7183 9225 7209 9231
rect 6673 9199 6679 9225
rect 6705 9199 6711 9225
rect 7065 9199 7071 9225
rect 7097 9199 7103 9225
rect 7183 9193 7209 9199
rect 9591 9225 9617 9231
rect 9591 9193 9617 9199
rect 11159 9225 11185 9231
rect 11159 9193 11185 9199
rect 11271 9225 11297 9231
rect 11271 9193 11297 9199
rect 11439 9225 11465 9231
rect 11439 9193 11465 9199
rect 12111 9225 12137 9231
rect 12111 9193 12137 9199
rect 13007 9225 13033 9231
rect 13007 9193 13033 9199
rect 13455 9225 13481 9231
rect 13455 9193 13481 9199
rect 13511 9225 13537 9231
rect 13511 9193 13537 9199
rect 13791 9225 13817 9231
rect 18825 9199 18831 9225
rect 18857 9199 18863 9225
rect 13791 9193 13817 9199
rect 9759 9169 9785 9175
rect 5609 9143 5615 9169
rect 5641 9143 5647 9169
rect 9759 9137 9785 9143
rect 12727 9169 12753 9175
rect 12727 9137 12753 9143
rect 13175 9169 13201 9175
rect 13175 9137 13201 9143
rect 20007 9169 20033 9175
rect 20007 9137 20033 9143
rect 11551 9113 11577 9119
rect 11551 9081 11577 9087
rect 12055 9113 12081 9119
rect 12055 9081 12081 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 967 8889 993 8895
rect 967 8857 993 8863
rect 10095 8889 10121 8895
rect 11097 8863 11103 8889
rect 11129 8863 11135 8889
rect 12161 8863 12167 8889
rect 12193 8863 12199 8889
rect 12721 8863 12727 8889
rect 12753 8863 12759 8889
rect 13785 8863 13791 8889
rect 13817 8863 13823 8889
rect 19945 8863 19951 8889
rect 19977 8863 19983 8889
rect 10095 8857 10121 8863
rect 6903 8833 6929 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 6903 8801 6929 8807
rect 7015 8833 7041 8839
rect 7015 8801 7041 8807
rect 7183 8833 7209 8839
rect 7457 8807 7463 8833
rect 7489 8807 7495 8833
rect 10705 8807 10711 8833
rect 10737 8807 10743 8833
rect 12329 8807 12335 8833
rect 12361 8807 12367 8833
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 7183 8801 7209 8807
rect 9417 8751 9423 8777
rect 9449 8751 9455 8777
rect 7127 8721 7153 8727
rect 9591 8721 9617 8727
rect 7345 8695 7351 8721
rect 7377 8695 7383 8721
rect 7127 8689 7153 8695
rect 9591 8689 9617 8695
rect 10151 8721 10177 8727
rect 10151 8689 10177 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 7407 8553 7433 8559
rect 7407 8521 7433 8527
rect 8079 8553 8105 8559
rect 8079 8521 8105 8527
rect 9983 8553 10009 8559
rect 9983 8521 10009 8527
rect 10151 8553 10177 8559
rect 10313 8527 10319 8553
rect 10345 8527 10351 8553
rect 10151 8521 10177 8527
rect 6729 8471 6735 8497
rect 6761 8471 6767 8497
rect 13001 8471 13007 8497
rect 13033 8471 13039 8497
rect 19665 8471 19671 8497
rect 19697 8471 19703 8497
rect 8191 8441 8217 8447
rect 9815 8441 9841 8447
rect 2137 8415 2143 8441
rect 2169 8415 2175 8441
rect 7065 8415 7071 8441
rect 7097 8415 7103 8441
rect 9473 8415 9479 8441
rect 9505 8415 9511 8441
rect 12609 8415 12615 8441
rect 12641 8415 12647 8441
rect 18937 8415 18943 8441
rect 18969 8415 18975 8441
rect 8191 8409 8217 8415
rect 9815 8409 9841 8415
rect 967 8385 993 8391
rect 7519 8385 7545 8391
rect 5665 8359 5671 8385
rect 5697 8359 5703 8385
rect 967 8353 993 8359
rect 7519 8353 7545 8359
rect 8135 8385 8161 8391
rect 8135 8353 8161 8359
rect 8303 8385 8329 8391
rect 8303 8353 8329 8359
rect 9143 8385 9169 8391
rect 9361 8359 9367 8385
rect 9393 8359 9399 8385
rect 14065 8359 14071 8385
rect 14097 8359 14103 8385
rect 9143 8353 9169 8359
rect 7351 8329 7377 8335
rect 7351 8297 7377 8303
rect 8415 8329 8441 8335
rect 8415 8297 8441 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 8577 8079 8583 8105
rect 8609 8079 8615 8105
rect 9641 8079 9647 8105
rect 9673 8079 9679 8105
rect 8185 8023 8191 8049
rect 8217 8023 8223 8049
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 8919 7769 8945 7775
rect 8919 7737 8945 7743
rect 9087 7713 9113 7719
rect 7233 7687 7239 7713
rect 7265 7687 7271 7713
rect 10761 7687 10767 7713
rect 10793 7687 10799 7713
rect 9087 7681 9113 7687
rect 6841 7631 6847 7657
rect 6873 7631 6879 7657
rect 11097 7631 11103 7657
rect 11129 7631 11135 7657
rect 8297 7575 8303 7601
rect 8329 7575 8335 7601
rect 9697 7575 9703 7601
rect 9729 7575 9735 7601
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 20119 2449 20145 2455
rect 20119 2417 20145 2423
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 8521 1751 8527 1777
rect 8553 1751 8559 1777
rect 9031 1665 9057 1671
rect 9031 1633 9057 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 11215 19111 11241 19137
rect 12783 19111 12809 19137
rect 10711 18999 10737 19025
rect 12279 18999 12305 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 11383 18719 11409 18745
rect 13119 18719 13145 18745
rect 11103 18607 11129 18633
rect 12615 18607 12641 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 855 18159 881 18185
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 10767 14015 10793 14041
rect 10823 13903 10849 13929
rect 10767 13791 10793 13817
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 10935 13511 10961 13537
rect 11103 13511 11129 13537
rect 10767 13455 10793 13481
rect 11271 13455 11297 13481
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 10879 13231 10905 13257
rect 11943 13175 11969 13201
rect 11999 13175 12025 13201
rect 13287 13175 13313 13201
rect 13343 13175 13369 13201
rect 9367 13119 9393 13145
rect 11831 13119 11857 13145
rect 13175 13119 13201 13145
rect 18831 13119 18857 13145
rect 9759 13063 9785 13089
rect 19951 13063 19977 13089
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 967 12783 993 12809
rect 9591 12783 9617 12809
rect 12391 12783 12417 12809
rect 14015 12783 14041 12809
rect 20007 12783 20033 12809
rect 2143 12727 2169 12753
rect 8135 12727 8161 12753
rect 9759 12727 9785 12753
rect 9927 12727 9953 12753
rect 10935 12727 10961 12753
rect 12615 12727 12641 12753
rect 18831 12727 18857 12753
rect 8527 12671 8553 12697
rect 11327 12671 11353 12697
rect 12951 12671 12977 12697
rect 9871 12615 9897 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 9647 12447 9673 12473
rect 11439 12447 11465 12473
rect 11831 12447 11857 12473
rect 8359 12391 8385 12417
rect 9367 12391 9393 12417
rect 9759 12391 9785 12417
rect 8079 12335 8105 12361
rect 8247 12335 8273 12361
rect 8415 12335 8441 12361
rect 9479 12335 9505 12361
rect 9815 12335 9841 12361
rect 11383 12335 11409 12361
rect 11495 12335 11521 12361
rect 11719 12335 11745 12361
rect 11943 12335 11969 12361
rect 12671 12335 12697 12361
rect 6679 12279 6705 12305
rect 7743 12279 7769 12305
rect 13007 12279 13033 12305
rect 14071 12279 14097 12305
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 9087 12055 9113 12081
rect 9591 12055 9617 12081
rect 13735 12055 13761 12081
rect 7743 11999 7769 12025
rect 12839 11999 12865 12025
rect 13287 11999 13313 12025
rect 20007 11999 20033 12025
rect 7687 11943 7713 11969
rect 7855 11943 7881 11969
rect 9423 11943 9449 11969
rect 13119 11943 13145 11969
rect 13567 11943 13593 11969
rect 13679 11943 13705 11969
rect 18831 11943 18857 11969
rect 7519 11887 7545 11913
rect 9143 11887 9169 11913
rect 9311 11887 9337 11913
rect 13231 11887 13257 11913
rect 13343 11887 13369 11913
rect 13735 11887 13761 11913
rect 9087 11831 9113 11857
rect 9759 11831 9785 11857
rect 9927 11831 9953 11857
rect 12783 11831 12809 11857
rect 12895 11831 12921 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 8247 11663 8273 11689
rect 9087 11607 9113 11633
rect 11887 11607 11913 11633
rect 11943 11607 11969 11633
rect 8135 11551 8161 11577
rect 9311 11551 9337 11577
rect 11775 11551 11801 11577
rect 18831 11551 18857 11577
rect 9703 11495 9729 11521
rect 10767 11495 10793 11521
rect 9143 11439 9169 11465
rect 20007 11439 20033 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 9479 11271 9505 11297
rect 10319 11271 10345 11297
rect 967 11215 993 11241
rect 7071 11215 7097 11241
rect 7239 11215 7265 11241
rect 7463 11215 7489 11241
rect 8751 11215 8777 11241
rect 9871 11215 9897 11241
rect 12335 11215 12361 11241
rect 20007 11215 20033 11241
rect 2143 11159 2169 11185
rect 7519 11159 7545 11185
rect 7631 11159 7657 11185
rect 7799 11159 7825 11185
rect 9311 11159 9337 11185
rect 9815 11159 9841 11185
rect 10151 11159 10177 11185
rect 10935 11159 10961 11185
rect 13231 11159 13257 11185
rect 18943 11159 18969 11185
rect 7407 11103 7433 11129
rect 9031 11103 9057 11129
rect 9199 11103 9225 11129
rect 10263 11103 10289 11129
rect 11271 11103 11297 11129
rect 7127 11047 7153 11073
rect 8863 11047 8889 11073
rect 8975 11047 9001 11073
rect 9927 11047 9953 11073
rect 10319 11047 10345 11073
rect 13119 11047 13145 11073
rect 13175 11047 13201 11073
rect 13343 11047 13369 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 7799 10879 7825 10905
rect 8191 10879 8217 10905
rect 9087 10879 9113 10905
rect 12615 10879 12641 10905
rect 7015 10823 7041 10849
rect 7743 10823 7769 10849
rect 7855 10823 7881 10849
rect 8303 10823 8329 10849
rect 8919 10823 8945 10849
rect 9199 10823 9225 10849
rect 13455 10823 13481 10849
rect 14855 10823 14881 10849
rect 15191 10823 15217 10849
rect 2143 10767 2169 10793
rect 7407 10767 7433 10793
rect 8079 10767 8105 10793
rect 8191 10767 8217 10793
rect 8807 10767 8833 10793
rect 9143 10767 9169 10793
rect 9423 10767 9449 10793
rect 9703 10767 9729 10793
rect 12727 10767 12753 10793
rect 12951 10767 12977 10793
rect 13063 10761 13089 10787
rect 14743 10767 14769 10793
rect 15079 10767 15105 10793
rect 18831 10767 18857 10793
rect 967 10711 993 10737
rect 5951 10711 5977 10737
rect 11663 10711 11689 10737
rect 12671 10711 12697 10737
rect 14519 10711 14545 10737
rect 20007 10711 20033 10737
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 7351 10487 7377 10513
rect 967 10431 993 10457
rect 4999 10431 5025 10457
rect 7463 10431 7489 10457
rect 7967 10431 7993 10457
rect 11271 10431 11297 10457
rect 20007 10431 20033 10457
rect 2143 10375 2169 10401
rect 6455 10375 6481 10401
rect 6847 10375 6873 10401
rect 7127 10375 7153 10401
rect 7575 10375 7601 10401
rect 10039 10375 10065 10401
rect 10879 10375 10905 10401
rect 11215 10375 11241 10401
rect 11551 10375 11577 10401
rect 11663 10375 11689 10401
rect 14631 10375 14657 10401
rect 14967 10375 14993 10401
rect 18831 10375 18857 10401
rect 6063 10319 6089 10345
rect 6735 10319 6761 10345
rect 7239 10319 7265 10345
rect 10711 10319 10737 10345
rect 12895 10319 12921 10345
rect 7295 10263 7321 10289
rect 10655 10263 10681 10289
rect 11047 10263 11073 10289
rect 11327 10263 11353 10289
rect 14743 10263 14769 10289
rect 15079 10263 15105 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 8359 10095 8385 10121
rect 14519 10095 14545 10121
rect 6735 10039 6761 10065
rect 6791 10039 6817 10065
rect 6847 10039 6873 10065
rect 7351 10039 7377 10065
rect 7743 10039 7769 10065
rect 10487 10039 10513 10065
rect 10655 10039 10681 10065
rect 10711 10039 10737 10065
rect 10823 10039 10849 10065
rect 11887 10039 11913 10065
rect 2143 9983 2169 10009
rect 7127 9983 7153 10009
rect 7239 9983 7265 10009
rect 7463 9983 7489 10009
rect 7855 9983 7881 10009
rect 8415 9983 8441 10009
rect 8863 9983 8889 10009
rect 9255 9983 9281 10009
rect 9479 9983 9505 10009
rect 9871 9983 9897 10009
rect 9983 9983 10009 10009
rect 10319 9983 10345 10009
rect 11999 9983 12025 10009
rect 12895 9983 12921 10009
rect 14463 9983 14489 10009
rect 18831 9983 18857 10009
rect 7295 9927 7321 9953
rect 9087 9927 9113 9953
rect 9647 9927 9673 9953
rect 13231 9927 13257 9953
rect 14295 9927 14321 9953
rect 20007 9927 20033 9953
rect 967 9871 993 9897
rect 8863 9871 8889 9897
rect 14519 9871 14545 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 6735 9703 6761 9729
rect 9311 9703 9337 9729
rect 10263 9703 10289 9729
rect 20007 9703 20033 9729
rect 9703 9647 9729 9673
rect 6903 9591 6929 9617
rect 8359 9591 8385 9617
rect 8639 9591 8665 9617
rect 8695 9591 8721 9617
rect 8919 9591 8945 9617
rect 9087 9591 9113 9617
rect 9423 9591 9449 9617
rect 9871 9591 9897 9617
rect 10207 9591 10233 9617
rect 12223 9591 12249 9617
rect 13623 9591 13649 9617
rect 13791 9591 13817 9617
rect 18831 9591 18857 9617
rect 8247 9535 8273 9561
rect 9031 9535 9057 9561
rect 9199 9535 9225 9561
rect 10151 9535 10177 9561
rect 13735 9535 13761 9561
rect 6791 9479 6817 9505
rect 8751 9479 8777 9505
rect 12391 9479 12417 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 9927 9311 9953 9337
rect 11103 9311 11129 9337
rect 12055 9311 12081 9337
rect 12783 9311 12809 9337
rect 13119 9311 13145 9337
rect 13231 9311 13257 9337
rect 7295 9255 7321 9281
rect 7351 9255 7377 9281
rect 9479 9255 9505 9281
rect 10039 9255 10065 9281
rect 10095 9255 10121 9281
rect 11719 9255 11745 9281
rect 11775 9255 11801 9281
rect 11887 9255 11913 9281
rect 12671 9255 12697 9281
rect 13623 9255 13649 9281
rect 13679 9255 13705 9281
rect 13903 9255 13929 9281
rect 13959 9255 13985 9281
rect 6679 9199 6705 9225
rect 7071 9199 7097 9225
rect 7183 9199 7209 9225
rect 9591 9199 9617 9225
rect 11159 9199 11185 9225
rect 11271 9199 11297 9225
rect 11439 9199 11465 9225
rect 12111 9199 12137 9225
rect 13007 9199 13033 9225
rect 13455 9199 13481 9225
rect 13511 9199 13537 9225
rect 13791 9199 13817 9225
rect 18831 9199 18857 9225
rect 5615 9143 5641 9169
rect 9759 9143 9785 9169
rect 12727 9143 12753 9169
rect 13175 9143 13201 9169
rect 20007 9143 20033 9169
rect 11551 9087 11577 9113
rect 12055 9087 12081 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 967 8863 993 8889
rect 10095 8863 10121 8889
rect 11103 8863 11129 8889
rect 12167 8863 12193 8889
rect 12727 8863 12753 8889
rect 13791 8863 13817 8889
rect 19951 8863 19977 8889
rect 2143 8807 2169 8833
rect 6903 8807 6929 8833
rect 7015 8807 7041 8833
rect 7183 8807 7209 8833
rect 7463 8807 7489 8833
rect 10711 8807 10737 8833
rect 12335 8807 12361 8833
rect 18831 8807 18857 8833
rect 9423 8751 9449 8777
rect 7127 8695 7153 8721
rect 7351 8695 7377 8721
rect 9591 8695 9617 8721
rect 10151 8695 10177 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7407 8527 7433 8553
rect 8079 8527 8105 8553
rect 9983 8527 10009 8553
rect 10151 8527 10177 8553
rect 10319 8527 10345 8553
rect 6735 8471 6761 8497
rect 13007 8471 13033 8497
rect 19671 8471 19697 8497
rect 2143 8415 2169 8441
rect 7071 8415 7097 8441
rect 8191 8415 8217 8441
rect 9479 8415 9505 8441
rect 9815 8415 9841 8441
rect 12615 8415 12641 8441
rect 18943 8415 18969 8441
rect 967 8359 993 8385
rect 5671 8359 5697 8385
rect 7519 8359 7545 8385
rect 8135 8359 8161 8385
rect 8303 8359 8329 8385
rect 9143 8359 9169 8385
rect 9367 8359 9393 8385
rect 14071 8359 14097 8385
rect 7351 8303 7377 8329
rect 8415 8303 8441 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 8583 8079 8609 8105
rect 9647 8079 9673 8105
rect 8191 8023 8217 8049
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 8919 7743 8945 7769
rect 7239 7687 7265 7713
rect 9087 7687 9113 7713
rect 10767 7687 10793 7713
rect 6847 7631 6873 7657
rect 11103 7631 11129 7657
rect 8303 7575 8329 7601
rect 9703 7575 9729 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 20119 2423 20145 2449
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 8527 1751 8553 1777
rect 9031 1639 9057 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 10752 20600 10808 21000
rect 11088 20600 11144 21000
rect 11424 20600 11480 21000
rect 12096 20600 12152 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 10710 19025 10738 19031
rect 10710 18999 10711 19025
rect 10737 18999 10738 19025
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 854 18186 882 18191
rect 854 18139 882 18158
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 10150 13818 10178 13823
rect 10094 13790 10150 13818
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 10094 13258 10122 13790
rect 10150 13785 10178 13790
rect 10710 13482 10738 18999
rect 10766 18746 10794 20600
rect 11102 19138 11130 20600
rect 11214 19138 11242 19143
rect 11102 19137 11242 19138
rect 11102 19111 11215 19137
rect 11241 19111 11242 19137
rect 11102 19110 11242 19111
rect 11214 19105 11242 19110
rect 11438 19138 11466 20600
rect 11438 19105 11466 19110
rect 10766 18713 10794 18718
rect 11382 18746 11410 18751
rect 11382 18699 11410 18718
rect 12110 18746 12138 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 12110 18713 12138 18718
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 11102 18633 11130 18639
rect 11102 18607 11103 18633
rect 11129 18607 11130 18633
rect 10766 14042 10794 14047
rect 10766 13995 10794 14014
rect 11102 14042 11130 18607
rect 10822 13929 10850 13935
rect 10822 13903 10823 13929
rect 10849 13903 10850 13929
rect 10766 13818 10794 13823
rect 10766 13771 10794 13790
rect 10766 13482 10794 13487
rect 10710 13481 10794 13482
rect 10710 13455 10767 13481
rect 10793 13455 10794 13481
rect 10710 13454 10794 13455
rect 10766 13449 10794 13454
rect 9926 13230 10122 13258
rect 10822 13258 10850 13903
rect 10934 13538 10962 13543
rect 11102 13538 11130 14014
rect 8750 13146 8778 13151
rect 9366 13146 9394 13151
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 966 12809 994 12815
rect 966 12783 967 12809
rect 993 12783 994 12809
rect 966 12474 994 12783
rect 966 12441 994 12446
rect 2142 12753 2170 12759
rect 2142 12727 2143 12753
rect 2169 12727 2170 12753
rect 2142 12306 2170 12727
rect 8134 12753 8162 12759
rect 8134 12727 8135 12753
rect 8161 12727 8162 12753
rect 7910 12362 7938 12367
rect 8078 12362 8106 12367
rect 8134 12362 8162 12727
rect 8526 12697 8554 12703
rect 8526 12671 8527 12697
rect 8553 12671 8554 12697
rect 8526 12474 8554 12671
rect 8526 12441 8554 12446
rect 8358 12418 8386 12423
rect 8358 12371 8386 12390
rect 7854 12334 7910 12362
rect 2142 12273 2170 12278
rect 6678 12306 6706 12311
rect 6678 12259 6706 12278
rect 7742 12305 7770 12311
rect 7742 12279 7743 12305
rect 7769 12279 7770 12305
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 7742 12025 7770 12279
rect 7742 11999 7743 12025
rect 7769 11999 7770 12025
rect 7742 11993 7770 11999
rect 7686 11970 7714 11975
rect 7518 11913 7546 11919
rect 7518 11887 7519 11913
rect 7545 11887 7546 11913
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 7518 11298 7546 11887
rect 7518 11265 7546 11270
rect 966 11242 994 11247
rect 7070 11242 7098 11247
rect 966 11195 994 11214
rect 7014 11241 7098 11242
rect 7014 11215 7071 11241
rect 7097 11215 7098 11241
rect 7014 11214 7098 11215
rect 2142 11186 2170 11191
rect 2142 11139 2170 11158
rect 5950 11186 5978 11191
rect 2142 10793 2170 10799
rect 2142 10767 2143 10793
rect 2169 10767 2170 10793
rect 966 10738 994 10743
rect 966 10691 994 10710
rect 2142 10514 2170 10767
rect 5950 10737 5978 11158
rect 7014 10849 7042 11214
rect 7070 11209 7098 11214
rect 7238 11242 7266 11247
rect 7462 11242 7490 11247
rect 7238 11241 7490 11242
rect 7238 11215 7239 11241
rect 7265 11215 7463 11241
rect 7489 11215 7490 11241
rect 7238 11214 7490 11215
rect 7238 11209 7266 11214
rect 7462 11209 7490 11214
rect 7518 11186 7546 11191
rect 7518 11139 7546 11158
rect 7630 11185 7658 11191
rect 7630 11159 7631 11185
rect 7657 11159 7658 11185
rect 7406 11130 7434 11135
rect 7406 11083 7434 11102
rect 7014 10823 7015 10849
rect 7041 10823 7042 10849
rect 7014 10817 7042 10823
rect 7126 11073 7154 11079
rect 7126 11047 7127 11073
rect 7153 11047 7154 11073
rect 5950 10711 5951 10737
rect 5977 10711 5978 10737
rect 5950 10705 5978 10711
rect 6454 10794 6482 10799
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 2142 10481 2170 10486
rect 966 10458 994 10463
rect 966 10411 994 10430
rect 4998 10457 5026 10463
rect 4998 10431 4999 10457
rect 5025 10431 5026 10457
rect 2142 10402 2170 10407
rect 2142 10355 2170 10374
rect 4998 10402 5026 10431
rect 4998 10369 5026 10374
rect 6454 10401 6482 10766
rect 7126 10626 7154 11047
rect 7630 10962 7658 11159
rect 7686 11130 7714 11942
rect 7854 11969 7882 12334
rect 7910 12329 7938 12334
rect 7966 12361 8162 12362
rect 7966 12335 8079 12361
rect 8105 12335 8162 12361
rect 7966 12334 8162 12335
rect 8246 12362 8274 12367
rect 7854 11943 7855 11969
rect 7881 11943 7882 11969
rect 7854 11937 7882 11943
rect 7686 11097 7714 11102
rect 7798 11185 7826 11191
rect 7798 11159 7799 11185
rect 7825 11159 7826 11185
rect 7462 10934 7658 10962
rect 7350 10906 7378 10911
rect 7126 10593 7154 10598
rect 7182 10794 7210 10799
rect 6454 10375 6455 10401
rect 6481 10375 6482 10401
rect 6454 10369 6482 10375
rect 6734 10514 6762 10519
rect 6062 10345 6090 10351
rect 6062 10319 6063 10345
rect 6089 10319 6090 10345
rect 6062 10066 6090 10319
rect 6734 10345 6762 10486
rect 6846 10402 6874 10407
rect 6846 10355 6874 10374
rect 7126 10402 7154 10407
rect 7126 10355 7154 10374
rect 6734 10319 6735 10345
rect 6761 10319 6762 10345
rect 6734 10313 6762 10319
rect 6902 10178 6930 10183
rect 6846 10150 6902 10178
rect 6062 10033 6090 10038
rect 6734 10065 6762 10071
rect 6734 10039 6735 10065
rect 6761 10039 6762 10065
rect 2142 10010 2170 10015
rect 2142 9963 2170 9982
rect 5614 10010 5642 10015
rect 966 9898 994 9903
rect 966 9851 994 9870
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 5614 9169 5642 9982
rect 6734 9954 6762 10039
rect 6790 10066 6818 10071
rect 6790 10019 6818 10038
rect 6846 10065 6874 10150
rect 6902 10145 6930 10150
rect 6846 10039 6847 10065
rect 6873 10039 6874 10065
rect 6846 10033 6874 10039
rect 7126 10010 7154 10015
rect 7126 9963 7154 9982
rect 6734 9730 6762 9926
rect 6734 9729 6874 9730
rect 6734 9703 6735 9729
rect 6761 9703 6874 9729
rect 6734 9702 6874 9703
rect 6734 9697 6762 9702
rect 6790 9505 6818 9511
rect 6790 9479 6791 9505
rect 6817 9479 6818 9505
rect 6790 9338 6818 9479
rect 6678 9310 6818 9338
rect 6678 9225 6706 9310
rect 6678 9199 6679 9225
rect 6705 9199 6706 9225
rect 6678 9193 6706 9199
rect 5614 9143 5615 9169
rect 5641 9143 5642 9169
rect 5614 9137 5642 9143
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 966 8890 994 8895
rect 966 8843 994 8862
rect 2142 8834 2170 8839
rect 2142 8787 2170 8806
rect 5670 8834 5698 8839
rect 6846 8834 6874 9702
rect 6902 9618 6930 9623
rect 6902 9571 6930 9590
rect 7182 9338 7210 10766
rect 7350 10513 7378 10878
rect 7406 10794 7434 10799
rect 7406 10747 7434 10766
rect 7350 10487 7351 10513
rect 7377 10487 7378 10513
rect 7350 10481 7378 10487
rect 7462 10457 7490 10934
rect 7798 10905 7826 11159
rect 7798 10879 7799 10905
rect 7825 10879 7826 10905
rect 7798 10873 7826 10879
rect 7854 10962 7882 10967
rect 7742 10850 7770 10855
rect 7462 10431 7463 10457
rect 7489 10431 7490 10457
rect 7238 10345 7266 10351
rect 7238 10319 7239 10345
rect 7265 10319 7266 10345
rect 7238 10009 7266 10319
rect 7294 10289 7322 10295
rect 7294 10263 7295 10289
rect 7321 10263 7322 10289
rect 7294 10178 7322 10263
rect 7294 10145 7322 10150
rect 7350 10066 7378 10071
rect 7350 10019 7378 10038
rect 7238 9983 7239 10009
rect 7265 9983 7266 10009
rect 7238 9898 7266 9983
rect 7462 10010 7490 10431
rect 7574 10822 7742 10850
rect 7574 10401 7602 10822
rect 7742 10803 7770 10822
rect 7854 10849 7882 10934
rect 7854 10823 7855 10849
rect 7881 10823 7882 10849
rect 7854 10817 7882 10823
rect 7966 10794 7994 12334
rect 8078 12329 8106 12334
rect 8246 12315 8274 12334
rect 8414 12362 8442 12367
rect 8414 12315 8442 12334
rect 8246 11970 8274 11975
rect 8246 11689 8274 11942
rect 8246 11663 8247 11689
rect 8273 11663 8274 11689
rect 8246 11657 8274 11663
rect 8134 11578 8162 11583
rect 7574 10375 7575 10401
rect 7601 10375 7602 10401
rect 7574 10066 7602 10375
rect 7854 10626 7882 10631
rect 7574 10033 7602 10038
rect 7742 10065 7770 10071
rect 7742 10039 7743 10065
rect 7769 10039 7770 10065
rect 7462 9963 7490 9982
rect 7238 9865 7266 9870
rect 7294 9953 7322 9959
rect 7294 9927 7295 9953
rect 7321 9927 7322 9953
rect 7294 9618 7322 9927
rect 7406 9954 7434 9959
rect 7294 9585 7322 9590
rect 7350 9898 7378 9903
rect 7070 9310 7210 9338
rect 7070 9225 7098 9310
rect 7294 9281 7322 9287
rect 7294 9255 7295 9281
rect 7321 9255 7322 9281
rect 7070 9199 7071 9225
rect 7097 9199 7098 9225
rect 7014 8890 7042 8895
rect 6902 8834 6930 8839
rect 6846 8833 6930 8834
rect 6846 8807 6903 8833
rect 6929 8807 6930 8833
rect 6846 8806 6930 8807
rect 966 8442 994 8447
rect 966 8385 994 8414
rect 2142 8442 2170 8447
rect 2142 8395 2170 8414
rect 966 8359 967 8385
rect 993 8359 994 8385
rect 966 8353 994 8359
rect 5670 8385 5698 8806
rect 6902 8801 6930 8806
rect 7014 8833 7042 8862
rect 7014 8807 7015 8833
rect 7041 8807 7042 8833
rect 7014 8801 7042 8807
rect 6846 8722 6874 8727
rect 6734 8694 6846 8722
rect 6734 8497 6762 8694
rect 6846 8689 6874 8694
rect 6734 8471 6735 8497
rect 6761 8471 6762 8497
rect 6734 8465 6762 8471
rect 5670 8359 5671 8385
rect 5697 8359 5698 8385
rect 5670 8353 5698 8359
rect 7070 8441 7098 9199
rect 7182 9225 7210 9231
rect 7182 9199 7183 9225
rect 7209 9199 7210 9225
rect 7182 8833 7210 9199
rect 7182 8807 7183 8833
rect 7209 8807 7210 8833
rect 7182 8801 7210 8807
rect 7294 8834 7322 9255
rect 7350 9281 7378 9870
rect 7350 9255 7351 9281
rect 7377 9255 7378 9281
rect 7350 9249 7378 9255
rect 7294 8801 7322 8806
rect 7126 8722 7154 8727
rect 7126 8675 7154 8694
rect 7350 8721 7378 8727
rect 7350 8695 7351 8721
rect 7377 8695 7378 8721
rect 7070 8415 7071 8441
rect 7097 8415 7098 8441
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 6846 8050 6874 8055
rect 6846 7657 6874 8022
rect 7070 8050 7098 8415
rect 7350 8442 7378 8695
rect 7406 8553 7434 9926
rect 7742 9954 7770 10039
rect 7854 10009 7882 10598
rect 7966 10457 7994 10766
rect 8078 11550 8134 11578
rect 8078 10962 8106 11550
rect 8134 11531 8162 11550
rect 8750 11242 8778 13118
rect 9254 13145 9394 13146
rect 9254 13119 9367 13145
rect 9393 13119 9394 13145
rect 9254 13118 9394 13119
rect 9086 12418 9114 12423
rect 9086 12081 9114 12390
rect 9086 12055 9087 12081
rect 9113 12055 9114 12081
rect 9086 12049 9114 12055
rect 9142 11914 9170 11933
rect 9142 11881 9170 11886
rect 9086 11858 9114 11863
rect 9086 11802 9114 11830
rect 8750 11195 8778 11214
rect 8974 11774 9114 11802
rect 9142 11802 9170 11807
rect 8974 11130 9002 11774
rect 9086 11634 9114 11639
rect 9142 11634 9170 11774
rect 9086 11633 9170 11634
rect 9086 11607 9087 11633
rect 9113 11607 9170 11633
rect 9086 11606 9170 11607
rect 9086 11601 9114 11606
rect 9254 11578 9282 13118
rect 9366 13113 9394 13118
rect 9758 13089 9786 13095
rect 9758 13063 9759 13089
rect 9785 13063 9786 13089
rect 9590 12809 9618 12815
rect 9590 12783 9591 12809
rect 9617 12783 9618 12809
rect 9366 12417 9394 12423
rect 9366 12391 9367 12417
rect 9393 12391 9394 12417
rect 9310 11913 9338 11919
rect 9310 11887 9311 11913
rect 9337 11887 9338 11913
rect 9310 11746 9338 11887
rect 9366 11858 9394 12391
rect 9478 12362 9506 12367
rect 9590 12362 9618 12783
rect 9758 12753 9786 13063
rect 9758 12727 9759 12753
rect 9785 12727 9786 12753
rect 9758 12721 9786 12727
rect 9926 12753 9954 13230
rect 10822 13225 10850 13230
rect 10878 13537 11130 13538
rect 10878 13511 10935 13537
rect 10961 13511 11103 13537
rect 11129 13511 11130 13537
rect 10878 13510 11130 13511
rect 10878 13257 10906 13510
rect 10934 13505 10962 13510
rect 11102 13505 11130 13510
rect 11270 13482 11298 13487
rect 11270 13435 11298 13454
rect 12278 13482 12306 18999
rect 13118 18746 13146 18751
rect 13118 18699 13146 18718
rect 12614 18633 12642 18639
rect 12614 18607 12615 18633
rect 12641 18607 12642 18633
rect 12614 13454 12642 18607
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 12278 13449 12306 13454
rect 12390 13426 12642 13454
rect 10878 13231 10879 13257
rect 10905 13231 10906 13257
rect 10878 13225 10906 13231
rect 11998 13258 12026 13263
rect 11942 13202 11970 13207
rect 11942 13155 11970 13174
rect 11998 13201 12026 13230
rect 11998 13175 11999 13201
rect 12025 13175 12026 13201
rect 11830 13146 11858 13151
rect 11718 13145 11858 13146
rect 11718 13119 11831 13145
rect 11857 13119 11858 13145
rect 11718 13118 11858 13119
rect 9926 12727 9927 12753
rect 9953 12727 9954 12753
rect 9926 12721 9954 12727
rect 10934 12753 10962 12759
rect 10934 12727 10935 12753
rect 10961 12727 10962 12753
rect 9870 12642 9898 12647
rect 9814 12641 9898 12642
rect 9814 12615 9871 12641
rect 9897 12615 9898 12641
rect 9814 12614 9898 12615
rect 9646 12474 9674 12479
rect 9646 12427 9674 12446
rect 9758 12418 9786 12423
rect 9758 12371 9786 12390
rect 9478 12361 9618 12362
rect 9478 12335 9479 12361
rect 9505 12335 9618 12361
rect 9478 12334 9618 12335
rect 9814 12361 9842 12614
rect 9870 12609 9898 12614
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9814 12335 9815 12361
rect 9841 12335 9842 12361
rect 9366 11825 9394 11830
rect 9422 11969 9450 11975
rect 9422 11943 9423 11969
rect 9449 11943 9450 11969
rect 9310 11713 9338 11718
rect 9310 11578 9338 11583
rect 9254 11577 9338 11578
rect 9254 11551 9311 11577
rect 9337 11551 9338 11577
rect 9254 11550 9338 11551
rect 9142 11465 9170 11471
rect 9142 11439 9143 11465
rect 9169 11439 9170 11465
rect 8862 11074 8890 11079
rect 8974 11074 9002 11102
rect 8078 10793 8106 10934
rect 8806 11073 8890 11074
rect 8806 11047 8863 11073
rect 8889 11047 8890 11073
rect 8806 11046 8890 11047
rect 8806 11018 8834 11046
rect 8862 11041 8890 11046
rect 8918 11073 9002 11074
rect 8918 11047 8975 11073
rect 9001 11047 9002 11073
rect 8918 11046 9002 11047
rect 8190 10906 8218 10911
rect 8190 10859 8218 10878
rect 8078 10767 8079 10793
rect 8105 10767 8106 10793
rect 8078 10761 8106 10767
rect 8134 10850 8162 10855
rect 8134 10794 8162 10822
rect 8302 10850 8330 10855
rect 8190 10794 8218 10799
rect 8134 10793 8274 10794
rect 8134 10767 8191 10793
rect 8217 10767 8274 10793
rect 8134 10766 8274 10767
rect 8190 10761 8218 10766
rect 7966 10431 7967 10457
rect 7993 10431 7994 10457
rect 7966 10425 7994 10431
rect 7854 9983 7855 10009
rect 7881 9983 7882 10009
rect 7854 9977 7882 9983
rect 7742 9921 7770 9926
rect 8246 9561 8274 10766
rect 8302 10122 8330 10822
rect 8806 10793 8834 10990
rect 8862 10962 8890 10967
rect 8918 10962 8946 11046
rect 8974 11041 9002 11046
rect 9030 11129 9058 11135
rect 9030 11103 9031 11129
rect 9057 11103 9058 11129
rect 8918 10934 9002 10962
rect 8862 10850 8890 10934
rect 8918 10850 8946 10855
rect 8862 10849 8946 10850
rect 8862 10823 8919 10849
rect 8945 10823 8946 10849
rect 8862 10822 8946 10823
rect 8918 10817 8946 10822
rect 8806 10767 8807 10793
rect 8833 10767 8834 10793
rect 8806 10761 8834 10767
rect 8358 10122 8386 10127
rect 8302 10121 8386 10122
rect 8302 10095 8359 10121
rect 8385 10095 8386 10121
rect 8302 10094 8386 10095
rect 8358 10066 8386 10094
rect 8358 10033 8386 10038
rect 8862 10066 8890 10071
rect 8414 10010 8442 10015
rect 8414 10009 8722 10010
rect 8414 9983 8415 10009
rect 8441 9983 8722 10009
rect 8414 9982 8722 9983
rect 8414 9977 8442 9982
rect 8638 9842 8666 9847
rect 8246 9535 8247 9561
rect 8273 9535 8274 9561
rect 8246 9529 8274 9535
rect 8358 9617 8386 9623
rect 8358 9591 8359 9617
rect 8385 9591 8386 9617
rect 8078 9506 8106 9511
rect 7462 8834 7490 8839
rect 7462 8787 7490 8806
rect 7406 8527 7407 8553
rect 7433 8527 7434 8553
rect 7406 8521 7434 8527
rect 8078 8553 8106 9478
rect 8358 9282 8386 9591
rect 8638 9617 8666 9814
rect 8638 9591 8639 9617
rect 8665 9591 8666 9617
rect 8638 9585 8666 9591
rect 8694 9617 8722 9982
rect 8862 10009 8890 10038
rect 8862 9983 8863 10009
rect 8889 9983 8890 10009
rect 8862 9977 8890 9983
rect 8862 9898 8890 9903
rect 8862 9851 8890 9870
rect 8694 9591 8695 9617
rect 8721 9591 8722 9617
rect 8358 9249 8386 9254
rect 8694 9226 8722 9591
rect 8918 9618 8946 9623
rect 8974 9618 9002 10934
rect 9030 10234 9058 11103
rect 9086 11018 9114 11023
rect 9086 10905 9114 10990
rect 9086 10879 9087 10905
rect 9113 10879 9114 10905
rect 9086 10873 9114 10879
rect 9142 10906 9170 11439
rect 9198 11130 9226 11135
rect 9198 11083 9226 11102
rect 9142 10873 9170 10878
rect 9198 10850 9226 10855
rect 9198 10803 9226 10822
rect 9142 10794 9170 10799
rect 9086 10793 9170 10794
rect 9086 10767 9143 10793
rect 9169 10767 9170 10793
rect 9086 10766 9170 10767
rect 9086 10738 9114 10766
rect 9142 10761 9170 10766
rect 9254 10794 9282 11550
rect 9310 11545 9338 11550
rect 9422 11578 9450 11943
rect 9478 11802 9506 12334
rect 9590 12082 9618 12087
rect 9814 12082 9842 12335
rect 9590 12081 9842 12082
rect 9590 12055 9591 12081
rect 9617 12055 9842 12081
rect 9590 12054 9842 12055
rect 9590 12049 9618 12054
rect 9478 11769 9506 11774
rect 9758 11857 9786 11863
rect 9926 11858 9954 11877
rect 9758 11831 9759 11857
rect 9785 11831 9786 11857
rect 9758 11746 9786 11831
rect 9758 11634 9786 11718
rect 9422 11298 9450 11550
rect 9646 11606 9786 11634
rect 9814 11830 9926 11858
rect 9646 11410 9674 11606
rect 9702 11522 9730 11527
rect 9702 11475 9730 11494
rect 9646 11382 9786 11410
rect 9478 11298 9506 11303
rect 9422 11297 9506 11298
rect 9422 11271 9479 11297
rect 9505 11271 9506 11297
rect 9422 11270 9506 11271
rect 9478 11265 9506 11270
rect 9702 11242 9730 11247
rect 9310 11186 9338 11191
rect 9310 11139 9338 11158
rect 9254 10761 9282 10766
rect 9422 10794 9450 10799
rect 9422 10747 9450 10766
rect 9702 10793 9730 11214
rect 9702 10767 9703 10793
rect 9729 10767 9730 10793
rect 9702 10761 9730 10767
rect 9758 11074 9786 11382
rect 9814 11185 9842 11830
rect 9926 11825 9954 11830
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9926 11690 9954 11695
rect 9870 11522 9898 11527
rect 9870 11241 9898 11494
rect 9870 11215 9871 11241
rect 9897 11215 9898 11241
rect 9870 11209 9898 11215
rect 9814 11159 9815 11185
rect 9841 11159 9842 11185
rect 9814 11153 9842 11159
rect 9926 11074 9954 11662
rect 10766 11522 10794 11527
rect 10710 11521 10794 11522
rect 10710 11495 10767 11521
rect 10793 11495 10794 11521
rect 10710 11494 10794 11495
rect 10318 11298 10346 11303
rect 10150 11297 10346 11298
rect 10150 11271 10319 11297
rect 10345 11271 10346 11297
rect 10150 11270 10346 11271
rect 10150 11185 10178 11270
rect 10318 11265 10346 11270
rect 10150 11159 10151 11185
rect 10177 11159 10178 11185
rect 10150 11153 10178 11159
rect 10710 11186 10738 11494
rect 10766 11489 10794 11494
rect 9086 10705 9114 10710
rect 9030 10201 9058 10206
rect 9198 10234 9226 10239
rect 9198 10094 9226 10206
rect 8918 9617 9002 9618
rect 8918 9591 8919 9617
rect 8945 9591 9002 9617
rect 8918 9590 9002 9591
rect 9086 10066 9114 10071
rect 9198 10066 9282 10094
rect 9086 9953 9114 10038
rect 9086 9927 9087 9953
rect 9113 9927 9114 9953
rect 9086 9617 9114 9927
rect 9254 10009 9282 10066
rect 9702 10066 9730 10071
rect 9254 9983 9255 10009
rect 9281 9983 9282 10009
rect 9254 9730 9282 9983
rect 9478 10010 9506 10015
rect 9478 9963 9506 9982
rect 9254 9697 9282 9702
rect 9310 9954 9338 9959
rect 9310 9729 9338 9926
rect 9646 9954 9674 9959
rect 9646 9907 9674 9926
rect 9310 9703 9311 9729
rect 9337 9703 9338 9729
rect 9310 9697 9338 9703
rect 9702 9673 9730 10038
rect 9702 9647 9703 9673
rect 9729 9647 9730 9673
rect 9702 9641 9730 9647
rect 9086 9591 9087 9617
rect 9113 9591 9114 9617
rect 8918 9585 8946 9590
rect 9086 9585 9114 9591
rect 9422 9617 9450 9623
rect 9422 9591 9423 9617
rect 9449 9591 9450 9617
rect 9030 9561 9058 9567
rect 9030 9535 9031 9561
rect 9057 9535 9058 9561
rect 8750 9506 8778 9511
rect 8750 9459 8778 9478
rect 9030 9506 9058 9535
rect 9030 9473 9058 9478
rect 9198 9561 9226 9567
rect 9198 9535 9199 9561
rect 9225 9535 9226 9561
rect 8694 9193 8722 9198
rect 8078 8527 8079 8553
rect 8105 8527 8106 8553
rect 8078 8521 8106 8527
rect 8302 8890 8330 8895
rect 7350 8409 7378 8414
rect 8190 8442 8218 8447
rect 8302 8442 8330 8862
rect 8190 8441 8274 8442
rect 8190 8415 8191 8441
rect 8217 8415 8274 8441
rect 8190 8414 8274 8415
rect 8190 8409 8218 8414
rect 7518 8386 7546 8391
rect 7518 8339 7546 8358
rect 8134 8386 8162 8391
rect 8134 8339 8162 8358
rect 7350 8330 7378 8335
rect 7070 8017 7098 8022
rect 7238 8329 7378 8330
rect 7238 8303 7351 8329
rect 7377 8303 7378 8329
rect 7238 8302 7378 8303
rect 7238 7713 7266 8302
rect 7350 8297 7378 8302
rect 8190 8050 8218 8055
rect 8190 8003 8218 8022
rect 7238 7687 7239 7713
rect 7265 7687 7266 7713
rect 7238 7681 7266 7687
rect 6846 7631 6847 7657
rect 6873 7631 6874 7657
rect 6846 7625 6874 7631
rect 8246 7602 8274 8414
rect 8302 8385 8330 8414
rect 9198 8442 9226 9535
rect 9422 9338 9450 9591
rect 9422 9305 9450 9310
rect 9702 9338 9730 9343
rect 9758 9338 9786 11046
rect 9814 11073 9954 11074
rect 9814 11047 9927 11073
rect 9953 11047 9954 11073
rect 9814 11046 9954 11047
rect 9814 10962 9842 11046
rect 9926 11041 9954 11046
rect 10262 11129 10290 11135
rect 10262 11103 10263 11129
rect 10289 11103 10290 11129
rect 10262 11074 10290 11103
rect 10262 11041 10290 11046
rect 10318 11074 10346 11079
rect 10318 11073 10402 11074
rect 10318 11047 10319 11073
rect 10345 11047 10402 11073
rect 10318 11046 10402 11047
rect 10318 11041 10346 11046
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 9814 10929 9842 10934
rect 9870 10906 9898 10911
rect 9870 10290 9898 10878
rect 10038 10402 10066 10407
rect 10038 10355 10066 10374
rect 9814 10262 9898 10290
rect 10262 10290 10290 10295
rect 9814 9618 9842 10262
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9982 10066 10010 10071
rect 9870 10010 9898 10015
rect 9870 10009 9954 10010
rect 9870 9983 9871 10009
rect 9897 9983 9954 10009
rect 9870 9982 9954 9983
rect 9870 9977 9898 9982
rect 9870 9618 9898 9623
rect 9814 9617 9898 9618
rect 9814 9591 9871 9617
rect 9897 9591 9898 9617
rect 9814 9590 9898 9591
rect 9926 9618 9954 9982
rect 9982 10009 10010 10038
rect 9982 9983 9983 10009
rect 10009 9983 10010 10009
rect 9982 9977 10010 9983
rect 10262 9730 10290 10262
rect 10374 10066 10402 11046
rect 10710 10346 10738 11158
rect 10934 11185 10962 12727
rect 11326 12698 11354 12703
rect 11326 12697 11466 12698
rect 11326 12671 11327 12697
rect 11353 12671 11466 12697
rect 11326 12670 11466 12671
rect 11326 12665 11354 12670
rect 11438 12473 11466 12670
rect 11438 12447 11439 12473
rect 11465 12447 11466 12473
rect 11438 12441 11466 12447
rect 11382 12361 11410 12367
rect 11382 12335 11383 12361
rect 11409 12335 11410 12361
rect 10934 11159 10935 11185
rect 10961 11159 10962 11185
rect 10878 10794 10906 10799
rect 10878 10401 10906 10766
rect 10878 10375 10879 10401
rect 10905 10375 10906 10401
rect 10710 10345 10794 10346
rect 10710 10319 10711 10345
rect 10737 10319 10794 10345
rect 10710 10318 10794 10319
rect 10710 10313 10738 10318
rect 10654 10290 10682 10295
rect 10654 10243 10682 10262
rect 10486 10066 10514 10071
rect 10654 10066 10682 10071
rect 10374 10065 10682 10066
rect 10374 10039 10487 10065
rect 10513 10039 10655 10065
rect 10681 10039 10682 10065
rect 10374 10038 10682 10039
rect 10318 10009 10346 10015
rect 10318 9983 10319 10009
rect 10345 9983 10346 10009
rect 10318 9842 10346 9983
rect 10486 9954 10514 10038
rect 10654 10033 10682 10038
rect 10710 10066 10738 10071
rect 10710 10019 10738 10038
rect 10486 9921 10514 9926
rect 10318 9809 10346 9814
rect 10710 9842 10738 9847
rect 10766 9842 10794 10318
rect 10822 10066 10850 10071
rect 10878 10066 10906 10375
rect 10822 10065 10906 10066
rect 10822 10039 10823 10065
rect 10849 10039 10906 10065
rect 10822 10038 10906 10039
rect 10822 10033 10850 10038
rect 10738 9814 10794 9842
rect 10710 9809 10738 9814
rect 10262 9683 10290 9702
rect 10206 9618 10234 9623
rect 9926 9590 10122 9618
rect 9870 9562 9898 9590
rect 9870 9529 9898 9534
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9926 9338 9954 9343
rect 9758 9337 9954 9338
rect 9758 9311 9927 9337
rect 9953 9311 9954 9337
rect 9758 9310 9954 9311
rect 9478 9282 9506 9287
rect 9702 9282 9730 9310
rect 9926 9305 9954 9310
rect 10038 9282 10066 9287
rect 9702 9254 9786 9282
rect 9478 9235 9506 9254
rect 9422 9226 9450 9231
rect 9422 8778 9450 9198
rect 9590 9226 9618 9231
rect 9590 9179 9618 9198
rect 9758 9169 9786 9254
rect 9758 9143 9759 9169
rect 9785 9143 9786 9169
rect 9758 9137 9786 9143
rect 9982 9254 10038 9282
rect 9982 8890 10010 9254
rect 10038 9235 10066 9254
rect 10094 9282 10122 9590
rect 10206 9571 10234 9590
rect 10150 9562 10178 9567
rect 10150 9515 10178 9534
rect 10318 9282 10346 9287
rect 10094 9281 10318 9282
rect 10094 9255 10095 9281
rect 10121 9255 10318 9281
rect 10094 9254 10318 9255
rect 10094 9249 10122 9254
rect 10094 8890 10122 8895
rect 9982 8889 10122 8890
rect 9982 8863 10095 8889
rect 10121 8863 10122 8889
rect 9982 8862 10122 8863
rect 9198 8409 9226 8414
rect 9366 8777 9450 8778
rect 9366 8751 9423 8777
rect 9449 8751 9450 8777
rect 9366 8750 9450 8751
rect 8302 8359 8303 8385
rect 8329 8359 8330 8385
rect 8302 8353 8330 8359
rect 9142 8385 9170 8391
rect 9142 8359 9143 8385
rect 9169 8359 9170 8385
rect 8414 8330 8442 8335
rect 8414 8329 8610 8330
rect 8414 8303 8415 8329
rect 8441 8303 8610 8329
rect 8414 8302 8610 8303
rect 8414 8297 8442 8302
rect 8582 8106 8610 8302
rect 8582 8105 8946 8106
rect 8582 8079 8583 8105
rect 8609 8079 8946 8105
rect 8582 8078 8946 8079
rect 8582 8073 8610 8078
rect 8918 7769 8946 8078
rect 8918 7743 8919 7769
rect 8945 7743 8946 7769
rect 8918 7737 8946 7743
rect 9086 7714 9114 7719
rect 9142 7714 9170 8359
rect 9366 8385 9394 8750
rect 9422 8745 9450 8750
rect 9590 8722 9618 8727
rect 9590 8721 9674 8722
rect 9590 8695 9591 8721
rect 9617 8695 9674 8721
rect 9590 8694 9674 8695
rect 9590 8689 9618 8694
rect 9646 8554 9674 8694
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9366 8359 9367 8385
rect 9393 8359 9394 8385
rect 9366 8353 9394 8359
rect 9478 8441 9506 8447
rect 9478 8415 9479 8441
rect 9505 8415 9506 8441
rect 9478 7994 9506 8415
rect 9646 8105 9674 8526
rect 9982 8554 10010 8559
rect 10094 8554 10122 8862
rect 10150 8722 10178 8727
rect 10150 8721 10234 8722
rect 10150 8695 10151 8721
rect 10177 8695 10234 8721
rect 10150 8694 10234 8695
rect 10150 8689 10178 8694
rect 9982 8553 10122 8554
rect 9982 8527 9983 8553
rect 10009 8527 10122 8553
rect 9982 8526 10122 8527
rect 10150 8554 10178 8559
rect 10206 8554 10234 8694
rect 10262 8554 10290 8559
rect 10206 8526 10262 8554
rect 9982 8521 10010 8526
rect 10150 8507 10178 8526
rect 10262 8521 10290 8526
rect 10318 8553 10346 9254
rect 10710 8833 10738 8839
rect 10710 8807 10711 8833
rect 10737 8807 10738 8833
rect 10710 8666 10738 8807
rect 10766 8666 10794 8671
rect 10710 8638 10766 8666
rect 10766 8633 10794 8638
rect 10934 8666 10962 11159
rect 11214 11858 11242 11863
rect 11382 11858 11410 12335
rect 11242 11830 11410 11858
rect 11494 12361 11522 12367
rect 11494 12335 11495 12361
rect 11521 12335 11522 12361
rect 11214 10401 11242 11830
rect 11494 11802 11522 12335
rect 11718 12361 11746 13118
rect 11830 13113 11858 13118
rect 11998 12978 12026 13175
rect 11830 12950 12026 12978
rect 12390 13202 12418 13426
rect 13342 13258 13370 13263
rect 11830 12473 11858 12950
rect 12390 12809 12418 13174
rect 13286 13202 13314 13207
rect 13286 13155 13314 13174
rect 13342 13201 13370 13230
rect 13342 13175 13343 13201
rect 13369 13175 13370 13201
rect 12390 12783 12391 12809
rect 12417 12783 12418 12809
rect 12390 12777 12418 12783
rect 13174 13145 13202 13151
rect 13174 13119 13175 13145
rect 13201 13119 13202 13145
rect 12614 12754 12642 12759
rect 12614 12753 12698 12754
rect 12614 12727 12615 12753
rect 12641 12727 12698 12753
rect 12614 12726 12698 12727
rect 12614 12721 12642 12726
rect 11830 12447 11831 12473
rect 11857 12447 11858 12473
rect 11830 12441 11858 12447
rect 11718 12335 11719 12361
rect 11745 12335 11746 12361
rect 11718 12329 11746 12335
rect 11942 12362 11970 12367
rect 11494 11769 11522 11774
rect 11886 11634 11914 11639
rect 11886 11587 11914 11606
rect 11942 11633 11970 12334
rect 12670 12361 12698 12726
rect 12950 12698 12978 12703
rect 12950 12697 13090 12698
rect 12950 12671 12951 12697
rect 12977 12671 13090 12697
rect 12950 12670 13090 12671
rect 12950 12665 12978 12670
rect 12670 12335 12671 12361
rect 12697 12335 12698 12361
rect 11942 11607 11943 11633
rect 11969 11607 11970 11633
rect 11774 11578 11802 11583
rect 11550 11577 11802 11578
rect 11550 11551 11775 11577
rect 11801 11551 11802 11577
rect 11550 11550 11802 11551
rect 11270 11129 11298 11135
rect 11270 11103 11271 11129
rect 11297 11103 11298 11129
rect 11270 10457 11298 11103
rect 11270 10431 11271 10457
rect 11297 10431 11298 10457
rect 11270 10425 11298 10431
rect 11214 10375 11215 10401
rect 11241 10375 11242 10401
rect 11214 10369 11242 10375
rect 11550 10401 11578 11550
rect 11774 11545 11802 11550
rect 11550 10375 11551 10401
rect 11577 10375 11578 10401
rect 11550 10369 11578 10375
rect 11662 10737 11690 10743
rect 11662 10711 11663 10737
rect 11689 10711 11690 10737
rect 11662 10402 11690 10711
rect 11662 10355 11690 10374
rect 11046 10289 11074 10295
rect 11046 10263 11047 10289
rect 11073 10263 11074 10289
rect 11046 10178 11074 10263
rect 11326 10289 11354 10295
rect 11326 10263 11327 10289
rect 11353 10263 11354 10289
rect 11326 10178 11354 10263
rect 11046 10150 11354 10178
rect 11102 9337 11130 9343
rect 11102 9311 11103 9337
rect 11129 9311 11130 9337
rect 11102 8889 11130 9311
rect 11158 9338 11186 9343
rect 11158 9225 11186 9310
rect 11326 9338 11354 10150
rect 11886 10066 11914 10071
rect 11942 10066 11970 11607
rect 12334 11634 12362 11639
rect 12334 11241 12362 11606
rect 12334 11215 12335 11241
rect 12361 11215 12362 11241
rect 12334 11209 12362 11215
rect 12614 11074 12642 11079
rect 12614 10905 12642 11046
rect 12614 10879 12615 10905
rect 12641 10879 12642 10905
rect 12614 10873 12642 10879
rect 12670 10906 12698 12335
rect 13006 12306 13034 12311
rect 12838 12305 13034 12306
rect 12838 12279 13007 12305
rect 13033 12279 13034 12305
rect 12838 12278 13034 12279
rect 12838 12025 12866 12278
rect 13006 12273 13034 12278
rect 12838 11999 12839 12025
rect 12865 11999 12866 12025
rect 12838 11993 12866 11999
rect 13062 12026 13090 12670
rect 13062 11993 13090 11998
rect 13118 11970 13146 11975
rect 13174 11970 13202 13119
rect 13342 12642 13370 13175
rect 14070 13146 14098 13151
rect 14014 12809 14042 12815
rect 14014 12783 14015 12809
rect 14041 12783 14042 12809
rect 14014 12754 14042 12783
rect 13790 12726 14014 12754
rect 13342 12614 13426 12642
rect 13398 12586 13426 12614
rect 13398 12558 13482 12586
rect 13286 12026 13314 12031
rect 13286 11979 13314 11998
rect 13118 11969 13202 11970
rect 13118 11943 13119 11969
rect 13145 11943 13202 11969
rect 13118 11942 13202 11943
rect 13454 11970 13482 12558
rect 13734 12082 13762 12087
rect 13118 11937 13146 11942
rect 13454 11937 13482 11942
rect 13566 12081 13762 12082
rect 13566 12055 13735 12081
rect 13761 12055 13762 12081
rect 13566 12054 13762 12055
rect 13566 11969 13594 12054
rect 13734 12049 13762 12054
rect 13566 11943 13567 11969
rect 13593 11943 13594 11969
rect 13566 11937 13594 11943
rect 13678 11970 13706 11975
rect 12726 11914 12754 11919
rect 12726 11018 12754 11886
rect 13230 11914 13258 11933
rect 13678 11923 13706 11942
rect 13230 11881 13258 11886
rect 13342 11913 13370 11919
rect 13342 11887 13343 11913
rect 13369 11887 13370 11913
rect 12782 11858 12810 11863
rect 12838 11858 12866 11863
rect 12782 11857 12838 11858
rect 12782 11831 12783 11857
rect 12809 11831 12838 11857
rect 12782 11830 12838 11831
rect 12782 11825 12810 11830
rect 12726 10985 12754 10990
rect 12670 10878 12810 10906
rect 12726 10793 12754 10799
rect 12726 10767 12727 10793
rect 12753 10767 12754 10793
rect 11886 10065 11970 10066
rect 11886 10039 11887 10065
rect 11913 10039 11970 10065
rect 11886 10038 11970 10039
rect 11886 10033 11914 10038
rect 11942 9338 11970 10038
rect 12670 10737 12698 10743
rect 12670 10711 12671 10737
rect 12697 10711 12698 10737
rect 11998 10009 12026 10015
rect 11998 9983 11999 10009
rect 12025 9983 12026 10009
rect 11998 9618 12026 9983
rect 12670 9954 12698 10711
rect 12726 10738 12754 10767
rect 12782 10794 12810 10878
rect 12782 10761 12810 10766
rect 12726 10705 12754 10710
rect 12838 10514 12866 11830
rect 12894 11857 12922 11863
rect 12894 11831 12895 11857
rect 12921 11831 12922 11857
rect 12894 11802 12922 11831
rect 13286 11858 13314 11863
rect 13342 11858 13370 11887
rect 13734 11914 13762 11919
rect 13790 11914 13818 12726
rect 14014 12721 14042 12726
rect 14070 12305 14098 13118
rect 18830 13146 18858 13151
rect 18830 13099 18858 13118
rect 19950 13089 19978 13095
rect 19950 13063 19951 13089
rect 19977 13063 19978 13089
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 19950 12810 19978 13063
rect 19950 12777 19978 12782
rect 20006 12809 20034 12815
rect 20006 12783 20007 12809
rect 20033 12783 20034 12809
rect 18830 12754 18858 12759
rect 18830 12707 18858 12726
rect 20006 12474 20034 12783
rect 20006 12441 20034 12446
rect 14070 12279 14071 12305
rect 14097 12279 14098 12305
rect 14070 12273 14098 12279
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 18830 11970 18858 11975
rect 13734 11913 13818 11914
rect 13734 11887 13735 11913
rect 13761 11887 13818 11913
rect 13734 11886 13818 11887
rect 18774 11969 18858 11970
rect 18774 11943 18831 11969
rect 18857 11943 18858 11969
rect 18774 11942 18858 11943
rect 13734 11881 13762 11886
rect 13314 11830 13370 11858
rect 13286 11825 13314 11830
rect 12894 11769 12922 11774
rect 13230 11802 13258 11807
rect 13230 11185 13258 11774
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 13230 11159 13231 11185
rect 13257 11159 13258 11185
rect 13230 11153 13258 11159
rect 13118 11074 13146 11079
rect 12670 9921 12698 9926
rect 12726 10486 12866 10514
rect 12950 10793 12978 10799
rect 12950 10767 12951 10793
rect 12977 10767 12978 10793
rect 11998 9585 12026 9590
rect 12222 9618 12250 9623
rect 12222 9571 12250 9590
rect 12390 9506 12418 9511
rect 12390 9459 12418 9478
rect 12054 9338 12082 9343
rect 11942 9310 12026 9338
rect 11326 9305 11354 9310
rect 11158 9199 11159 9225
rect 11185 9199 11186 9225
rect 11158 9193 11186 9199
rect 11270 9282 11298 9287
rect 11270 9225 11298 9254
rect 11718 9282 11746 9287
rect 11718 9235 11746 9254
rect 11774 9281 11802 9287
rect 11774 9255 11775 9281
rect 11801 9255 11802 9281
rect 11270 9199 11271 9225
rect 11297 9199 11298 9225
rect 11270 9193 11298 9199
rect 11438 9226 11466 9231
rect 11102 8863 11103 8889
rect 11129 8863 11130 8889
rect 11102 8857 11130 8863
rect 10934 8633 10962 8638
rect 11102 8666 11130 8671
rect 10318 8527 10319 8553
rect 10345 8527 10346 8553
rect 10318 8521 10346 8527
rect 10766 8554 10794 8559
rect 9646 8079 9647 8105
rect 9673 8079 9674 8105
rect 9646 8073 9674 8079
rect 9814 8441 9842 8447
rect 9814 8415 9815 8441
rect 9841 8415 9842 8441
rect 9814 7994 9842 8415
rect 9478 7966 9842 7994
rect 9086 7713 9170 7714
rect 9086 7687 9087 7713
rect 9113 7687 9170 7713
rect 9086 7686 9170 7687
rect 9086 7681 9114 7686
rect 8302 7602 8330 7607
rect 8246 7601 8330 7602
rect 8246 7575 8303 7601
rect 8329 7575 8330 7601
rect 8246 7574 8330 7575
rect 9702 7602 9730 7607
rect 9814 7602 9842 7966
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 10766 7713 10794 8526
rect 10766 7687 10767 7713
rect 10793 7687 10794 7713
rect 10766 7681 10794 7687
rect 11102 7657 11130 8638
rect 11438 8554 11466 9198
rect 11774 9226 11802 9255
rect 11886 9282 11914 9287
rect 11886 9235 11914 9254
rect 11998 9226 12026 9310
rect 12054 9337 12194 9338
rect 12054 9311 12055 9337
rect 12081 9311 12194 9337
rect 12054 9310 12194 9311
rect 12054 9305 12082 9310
rect 12110 9226 12138 9231
rect 11998 9225 12138 9226
rect 11998 9199 12111 9225
rect 12137 9199 12138 9225
rect 11998 9198 12138 9199
rect 11774 9193 11802 9198
rect 12110 9193 12138 9198
rect 11550 9114 11578 9119
rect 11550 9067 11578 9086
rect 12054 9114 12082 9119
rect 12054 9067 12082 9086
rect 12166 8946 12194 9310
rect 12670 9282 12698 9287
rect 12726 9282 12754 10486
rect 12950 10458 12978 10767
rect 13006 10794 13034 10799
rect 13034 10787 13090 10794
rect 13034 10766 13063 10787
rect 13006 10761 13034 10766
rect 13062 10761 13063 10766
rect 13089 10761 13090 10787
rect 12838 10430 12978 10458
rect 12838 9898 12866 10430
rect 12838 9865 12866 9870
rect 12894 10346 12922 10351
rect 13062 10346 13090 10761
rect 12894 10345 13090 10346
rect 12894 10319 12895 10345
rect 12921 10319 13090 10345
rect 12894 10318 13090 10319
rect 12894 10009 12922 10318
rect 12894 9983 12895 10009
rect 12921 9983 12922 10009
rect 12782 9338 12810 9343
rect 12782 9291 12810 9310
rect 12698 9254 12754 9282
rect 12670 9235 12698 9254
rect 12166 8889 12194 8918
rect 12166 8863 12167 8889
rect 12193 8863 12194 8889
rect 12166 8857 12194 8863
rect 12726 9169 12754 9175
rect 12726 9143 12727 9169
rect 12753 9143 12754 9169
rect 12726 8889 12754 9143
rect 12726 8863 12727 8889
rect 12753 8863 12754 8889
rect 12726 8857 12754 8863
rect 12334 8833 12362 8839
rect 12334 8807 12335 8833
rect 12361 8807 12362 8833
rect 12334 8666 12362 8807
rect 12334 8633 12362 8638
rect 12614 8666 12642 8671
rect 11438 8521 11466 8526
rect 12614 8441 12642 8638
rect 12894 8666 12922 9983
rect 13118 9394 13146 11046
rect 13174 11073 13202 11079
rect 13174 11047 13175 11073
rect 13201 11047 13202 11073
rect 13174 10962 13202 11047
rect 13342 11073 13370 11079
rect 13342 11047 13343 11073
rect 13369 11047 13370 11073
rect 13342 10962 13370 11047
rect 13174 10934 13314 10962
rect 13342 10934 13538 10962
rect 13286 10906 13314 10934
rect 13286 10878 13482 10906
rect 13454 10849 13482 10878
rect 13454 10823 13455 10849
rect 13481 10823 13482 10849
rect 13454 10817 13482 10823
rect 13510 10094 13538 10934
rect 14854 10850 14882 10855
rect 14854 10803 14882 10822
rect 15190 10849 15218 10855
rect 15190 10823 15191 10849
rect 15217 10823 15218 10849
rect 14742 10793 14770 10799
rect 14742 10767 14743 10793
rect 14769 10767 14770 10793
rect 14518 10738 14546 10743
rect 14462 10710 14518 10738
rect 14462 10178 14490 10710
rect 14518 10691 14546 10710
rect 14742 10738 14770 10767
rect 14742 10705 14770 10710
rect 15078 10793 15106 10799
rect 15078 10767 15079 10793
rect 15105 10767 15106 10793
rect 15078 10738 15106 10767
rect 15190 10794 15218 10823
rect 18774 10850 18802 11942
rect 18830 11937 18858 11942
rect 20006 11802 20034 11999
rect 20006 11769 20034 11774
rect 18830 11578 18858 11583
rect 18830 11531 18858 11550
rect 20006 11466 20034 11471
rect 20006 11419 20034 11438
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 18774 10817 18802 10822
rect 18942 11185 18970 11191
rect 18942 11159 18943 11185
rect 18969 11159 18970 11185
rect 15190 10761 15218 10766
rect 18830 10794 18858 10799
rect 18830 10747 18858 10766
rect 15078 10705 15106 10710
rect 18942 10738 18970 11159
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 18942 10705 18970 10710
rect 20006 10794 20034 10799
rect 20006 10737 20034 10766
rect 20006 10711 20007 10737
rect 20033 10711 20034 10737
rect 20006 10705 20034 10711
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 20006 10458 20034 10463
rect 20006 10411 20034 10430
rect 14630 10402 14658 10407
rect 14966 10402 14994 10407
rect 14462 10145 14490 10150
rect 14518 10401 14994 10402
rect 14518 10375 14631 10401
rect 14657 10375 14967 10401
rect 14993 10375 14994 10401
rect 14518 10374 14994 10375
rect 14518 10121 14546 10374
rect 14630 10369 14658 10374
rect 14742 10290 14770 10295
rect 14742 10243 14770 10262
rect 14518 10095 14519 10121
rect 14545 10095 14546 10121
rect 14518 10094 14546 10095
rect 13510 10066 13650 10094
rect 13230 9954 13258 9959
rect 13230 9907 13258 9926
rect 13622 9617 13650 10066
rect 13622 9591 13623 9617
rect 13649 9591 13650 9617
rect 13622 9585 13650 9591
rect 13734 10066 13762 10071
rect 13734 9561 13762 10038
rect 14294 10066 14546 10094
rect 13734 9535 13735 9561
rect 13761 9535 13762 9561
rect 13734 9529 13762 9535
rect 13790 10010 13818 10015
rect 13790 9618 13818 9982
rect 14294 9953 14322 10066
rect 14462 10010 14490 10015
rect 14462 9963 14490 9982
rect 14966 10010 14994 10374
rect 18830 10402 18858 10407
rect 18830 10355 18858 10374
rect 14966 9977 14994 9982
rect 15078 10289 15106 10295
rect 15078 10263 15079 10289
rect 15105 10263 15106 10289
rect 14294 9927 14295 9953
rect 14321 9927 14322 9953
rect 14294 9921 14322 9927
rect 14518 9898 14546 9903
rect 14518 9851 14546 9870
rect 15078 9618 15106 10263
rect 20006 10066 20034 10071
rect 18830 10010 18858 10015
rect 18830 9963 18858 9982
rect 20006 9953 20034 10038
rect 20006 9927 20007 9953
rect 20033 9927 20034 9953
rect 20006 9921 20034 9927
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 20006 9786 20034 9791
rect 20006 9729 20034 9758
rect 20006 9703 20007 9729
rect 20033 9703 20034 9729
rect 20006 9697 20034 9703
rect 13790 9617 13986 9618
rect 13790 9591 13791 9617
rect 13817 9591 13986 9617
rect 13790 9590 13986 9591
rect 13118 9337 13146 9366
rect 13678 9506 13706 9511
rect 13678 9450 13706 9478
rect 13790 9450 13818 9590
rect 13678 9422 13818 9450
rect 13118 9311 13119 9337
rect 13145 9311 13146 9337
rect 13118 9305 13146 9311
rect 13230 9338 13258 9343
rect 13230 9291 13258 9310
rect 13622 9281 13650 9287
rect 13622 9255 13623 9281
rect 13649 9255 13650 9281
rect 13006 9226 13034 9231
rect 13006 9179 13034 9198
rect 13454 9226 13482 9231
rect 13454 9179 13482 9198
rect 13510 9225 13538 9231
rect 13510 9199 13511 9225
rect 13537 9199 13538 9225
rect 12894 8633 12922 8638
rect 13174 9169 13202 9175
rect 13174 9143 13175 9169
rect 13201 9143 13202 9169
rect 13006 8498 13034 8503
rect 13174 8498 13202 9143
rect 13510 9170 13538 9199
rect 13510 9137 13538 9142
rect 13622 8890 13650 9255
rect 13678 9281 13706 9422
rect 13678 9255 13679 9281
rect 13705 9255 13706 9281
rect 13678 9249 13706 9255
rect 13902 9281 13930 9287
rect 13902 9255 13903 9281
rect 13929 9255 13930 9281
rect 13790 9226 13818 9231
rect 13790 9179 13818 9198
rect 13790 8890 13818 8895
rect 13622 8862 13790 8890
rect 13790 8843 13818 8862
rect 13902 8834 13930 9255
rect 13958 9281 13986 9590
rect 15078 9585 15106 9590
rect 18830 9618 18858 9623
rect 18830 9571 18858 9590
rect 13958 9255 13959 9281
rect 13985 9255 13986 9281
rect 13958 9249 13986 9255
rect 20006 9450 20034 9455
rect 18830 9225 18858 9231
rect 18830 9199 18831 9225
rect 18857 9199 18858 9225
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 18830 8946 18858 9199
rect 20006 9169 20034 9422
rect 20006 9143 20007 9169
rect 20033 9143 20034 9169
rect 20006 9137 20034 9143
rect 18830 8913 18858 8918
rect 19950 9114 19978 9119
rect 18942 8890 18970 8895
rect 14070 8834 14098 8839
rect 13902 8806 14070 8834
rect 13006 8497 13202 8498
rect 13006 8471 13007 8497
rect 13033 8471 13202 8497
rect 13006 8470 13202 8471
rect 13006 8465 13034 8470
rect 12614 8415 12615 8441
rect 12641 8415 12642 8441
rect 12614 8409 12642 8415
rect 14070 8385 14098 8806
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 18942 8441 18970 8862
rect 19950 8889 19978 9086
rect 19950 8863 19951 8889
rect 19977 8863 19978 8889
rect 19950 8857 19978 8863
rect 19670 8778 19698 8783
rect 19670 8497 19698 8750
rect 19670 8471 19671 8497
rect 19697 8471 19698 8497
rect 19670 8465 19698 8471
rect 18942 8415 18943 8441
rect 18969 8415 18970 8441
rect 18942 8409 18970 8415
rect 14070 8359 14071 8385
rect 14097 8359 14098 8385
rect 14070 8353 14098 8359
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 11102 7631 11103 7657
rect 11129 7631 11130 7657
rect 11102 7625 11130 7631
rect 9702 7601 9842 7602
rect 9702 7575 9703 7601
rect 9729 7575 9842 7601
rect 9702 7574 9842 7575
rect 8302 7546 8442 7574
rect 9702 7569 9730 7574
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 8414 4214 8442 7546
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 8414 4186 8554 4214
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8526 1777 8554 4186
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 20118 2449 20146 2455
rect 20118 2423 20119 2449
rect 20145 2423 20146 2449
rect 20118 2394 20146 2423
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 20118 2361 20146 2366
rect 9918 2333 10050 2338
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 8526 1751 8527 1777
rect 8553 1751 8554 1777
rect 8526 1745 8554 1751
rect 8414 1722 8442 1727
rect 8414 400 8442 1694
rect 9030 1722 9058 1727
rect 9030 1665 9058 1694
rect 9030 1639 9031 1665
rect 9057 1639 9058 1665
rect 9030 1633 9058 1639
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 8400 0 8456 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 854 18185 882 18186
rect 854 18159 855 18185
rect 855 18159 881 18185
rect 881 18159 882 18185
rect 854 18158 882 18159
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 10150 13790 10178 13818
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 11438 19110 11466 19138
rect 10766 18718 10794 18746
rect 11382 18745 11410 18746
rect 11382 18719 11383 18745
rect 11383 18719 11409 18745
rect 11409 18719 11410 18745
rect 11382 18718 11410 18719
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 12110 18718 12138 18746
rect 10766 14041 10794 14042
rect 10766 14015 10767 14041
rect 10767 14015 10793 14041
rect 10793 14015 10794 14041
rect 10766 14014 10794 14015
rect 11102 14014 11130 14042
rect 10766 13817 10794 13818
rect 10766 13791 10767 13817
rect 10767 13791 10793 13817
rect 10793 13791 10794 13817
rect 10766 13790 10794 13791
rect 10822 13230 10850 13258
rect 8750 13118 8778 13146
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 966 12446 994 12474
rect 8526 12446 8554 12474
rect 8358 12417 8386 12418
rect 8358 12391 8359 12417
rect 8359 12391 8385 12417
rect 8385 12391 8386 12417
rect 8358 12390 8386 12391
rect 7910 12334 7938 12362
rect 2142 12278 2170 12306
rect 6678 12305 6706 12306
rect 6678 12279 6679 12305
rect 6679 12279 6705 12305
rect 6705 12279 6706 12305
rect 6678 12278 6706 12279
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 7686 11969 7714 11970
rect 7686 11943 7687 11969
rect 7687 11943 7713 11969
rect 7713 11943 7714 11969
rect 7686 11942 7714 11943
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 7518 11270 7546 11298
rect 966 11241 994 11242
rect 966 11215 967 11241
rect 967 11215 993 11241
rect 993 11215 994 11241
rect 966 11214 994 11215
rect 2142 11185 2170 11186
rect 2142 11159 2143 11185
rect 2143 11159 2169 11185
rect 2169 11159 2170 11185
rect 2142 11158 2170 11159
rect 5950 11158 5978 11186
rect 966 10737 994 10738
rect 966 10711 967 10737
rect 967 10711 993 10737
rect 993 10711 994 10737
rect 966 10710 994 10711
rect 7518 11185 7546 11186
rect 7518 11159 7519 11185
rect 7519 11159 7545 11185
rect 7545 11159 7546 11185
rect 7518 11158 7546 11159
rect 7406 11129 7434 11130
rect 7406 11103 7407 11129
rect 7407 11103 7433 11129
rect 7433 11103 7434 11129
rect 7406 11102 7434 11103
rect 6454 10766 6482 10794
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 2142 10486 2170 10514
rect 966 10457 994 10458
rect 966 10431 967 10457
rect 967 10431 993 10457
rect 993 10431 994 10457
rect 966 10430 994 10431
rect 2142 10401 2170 10402
rect 2142 10375 2143 10401
rect 2143 10375 2169 10401
rect 2169 10375 2170 10401
rect 2142 10374 2170 10375
rect 4998 10374 5026 10402
rect 8246 12361 8274 12362
rect 8246 12335 8247 12361
rect 8247 12335 8273 12361
rect 8273 12335 8274 12361
rect 8246 12334 8274 12335
rect 7686 11102 7714 11130
rect 7350 10878 7378 10906
rect 7126 10598 7154 10626
rect 7182 10766 7210 10794
rect 6734 10486 6762 10514
rect 6846 10401 6874 10402
rect 6846 10375 6847 10401
rect 6847 10375 6873 10401
rect 6873 10375 6874 10401
rect 6846 10374 6874 10375
rect 7126 10401 7154 10402
rect 7126 10375 7127 10401
rect 7127 10375 7153 10401
rect 7153 10375 7154 10401
rect 7126 10374 7154 10375
rect 6902 10150 6930 10178
rect 6062 10038 6090 10066
rect 2142 10009 2170 10010
rect 2142 9983 2143 10009
rect 2143 9983 2169 10009
rect 2169 9983 2170 10009
rect 2142 9982 2170 9983
rect 5614 9982 5642 10010
rect 966 9897 994 9898
rect 966 9871 967 9897
rect 967 9871 993 9897
rect 993 9871 994 9897
rect 966 9870 994 9871
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 6790 10065 6818 10066
rect 6790 10039 6791 10065
rect 6791 10039 6817 10065
rect 6817 10039 6818 10065
rect 6790 10038 6818 10039
rect 7126 10009 7154 10010
rect 7126 9983 7127 10009
rect 7127 9983 7153 10009
rect 7153 9983 7154 10009
rect 7126 9982 7154 9983
rect 6734 9926 6762 9954
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 966 8889 994 8890
rect 966 8863 967 8889
rect 967 8863 993 8889
rect 993 8863 994 8889
rect 966 8862 994 8863
rect 2142 8833 2170 8834
rect 2142 8807 2143 8833
rect 2143 8807 2169 8833
rect 2169 8807 2170 8833
rect 2142 8806 2170 8807
rect 5670 8806 5698 8834
rect 6902 9617 6930 9618
rect 6902 9591 6903 9617
rect 6903 9591 6929 9617
rect 6929 9591 6930 9617
rect 6902 9590 6930 9591
rect 7406 10793 7434 10794
rect 7406 10767 7407 10793
rect 7407 10767 7433 10793
rect 7433 10767 7434 10793
rect 7406 10766 7434 10767
rect 7854 10934 7882 10962
rect 7294 10150 7322 10178
rect 7350 10065 7378 10066
rect 7350 10039 7351 10065
rect 7351 10039 7377 10065
rect 7377 10039 7378 10065
rect 7350 10038 7378 10039
rect 7742 10849 7770 10850
rect 7742 10823 7743 10849
rect 7743 10823 7769 10849
rect 7769 10823 7770 10849
rect 7742 10822 7770 10823
rect 8414 12361 8442 12362
rect 8414 12335 8415 12361
rect 8415 12335 8441 12361
rect 8441 12335 8442 12361
rect 8414 12334 8442 12335
rect 8246 11942 8274 11970
rect 7966 10766 7994 10794
rect 7854 10598 7882 10626
rect 7574 10038 7602 10066
rect 7462 10009 7490 10010
rect 7462 9983 7463 10009
rect 7463 9983 7489 10009
rect 7489 9983 7490 10009
rect 7462 9982 7490 9983
rect 7238 9870 7266 9898
rect 7406 9926 7434 9954
rect 7294 9590 7322 9618
rect 7350 9870 7378 9898
rect 7014 8862 7042 8890
rect 966 8414 994 8442
rect 2142 8441 2170 8442
rect 2142 8415 2143 8441
rect 2143 8415 2169 8441
rect 2169 8415 2170 8441
rect 2142 8414 2170 8415
rect 6846 8694 6874 8722
rect 7294 8806 7322 8834
rect 7126 8721 7154 8722
rect 7126 8695 7127 8721
rect 7127 8695 7153 8721
rect 7153 8695 7154 8721
rect 7126 8694 7154 8695
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 6846 8022 6874 8050
rect 8134 11577 8162 11578
rect 8134 11551 8135 11577
rect 8135 11551 8161 11577
rect 8161 11551 8162 11577
rect 8134 11550 8162 11551
rect 9086 12390 9114 12418
rect 9142 11913 9170 11914
rect 9142 11887 9143 11913
rect 9143 11887 9169 11913
rect 9169 11887 9170 11913
rect 9142 11886 9170 11887
rect 9086 11857 9114 11858
rect 9086 11831 9087 11857
rect 9087 11831 9113 11857
rect 9113 11831 9114 11857
rect 9086 11830 9114 11831
rect 8750 11241 8778 11242
rect 8750 11215 8751 11241
rect 8751 11215 8777 11241
rect 8777 11215 8778 11241
rect 8750 11214 8778 11215
rect 9142 11774 9170 11802
rect 11270 13481 11298 13482
rect 11270 13455 11271 13481
rect 11271 13455 11297 13481
rect 11297 13455 11298 13481
rect 11270 13454 11298 13455
rect 13118 18745 13146 18746
rect 13118 18719 13119 18745
rect 13119 18719 13145 18745
rect 13145 18719 13146 18745
rect 13118 18718 13146 18719
rect 12278 13454 12306 13482
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 11998 13230 12026 13258
rect 11942 13201 11970 13202
rect 11942 13175 11943 13201
rect 11943 13175 11969 13201
rect 11969 13175 11970 13201
rect 11942 13174 11970 13175
rect 9646 12473 9674 12474
rect 9646 12447 9647 12473
rect 9647 12447 9673 12473
rect 9673 12447 9674 12473
rect 9646 12446 9674 12447
rect 9758 12417 9786 12418
rect 9758 12391 9759 12417
rect 9759 12391 9785 12417
rect 9785 12391 9786 12417
rect 9758 12390 9786 12391
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9366 11830 9394 11858
rect 9310 11718 9338 11746
rect 8974 11102 9002 11130
rect 8078 10934 8106 10962
rect 8806 10990 8834 11018
rect 8190 10905 8218 10906
rect 8190 10879 8191 10905
rect 8191 10879 8217 10905
rect 8217 10879 8218 10905
rect 8190 10878 8218 10879
rect 8134 10822 8162 10850
rect 8302 10849 8330 10850
rect 8302 10823 8303 10849
rect 8303 10823 8329 10849
rect 8329 10823 8330 10849
rect 8302 10822 8330 10823
rect 7742 9926 7770 9954
rect 8862 10934 8890 10962
rect 8358 10038 8386 10066
rect 8862 10038 8890 10066
rect 8638 9814 8666 9842
rect 8078 9478 8106 9506
rect 7462 8833 7490 8834
rect 7462 8807 7463 8833
rect 7463 8807 7489 8833
rect 7489 8807 7490 8833
rect 7462 8806 7490 8807
rect 8862 9897 8890 9898
rect 8862 9871 8863 9897
rect 8863 9871 8889 9897
rect 8889 9871 8890 9897
rect 8862 9870 8890 9871
rect 8358 9254 8386 9282
rect 9086 10990 9114 11018
rect 9198 11129 9226 11130
rect 9198 11103 9199 11129
rect 9199 11103 9225 11129
rect 9225 11103 9226 11129
rect 9198 11102 9226 11103
rect 9142 10878 9170 10906
rect 9198 10849 9226 10850
rect 9198 10823 9199 10849
rect 9199 10823 9225 10849
rect 9225 10823 9226 10849
rect 9198 10822 9226 10823
rect 9478 11774 9506 11802
rect 9758 11718 9786 11746
rect 9422 11550 9450 11578
rect 9926 11857 9954 11858
rect 9926 11831 9927 11857
rect 9927 11831 9953 11857
rect 9953 11831 9954 11857
rect 9926 11830 9954 11831
rect 9702 11521 9730 11522
rect 9702 11495 9703 11521
rect 9703 11495 9729 11521
rect 9729 11495 9730 11521
rect 9702 11494 9730 11495
rect 9702 11214 9730 11242
rect 9310 11185 9338 11186
rect 9310 11159 9311 11185
rect 9311 11159 9337 11185
rect 9337 11159 9338 11185
rect 9310 11158 9338 11159
rect 9254 10766 9282 10794
rect 9422 10793 9450 10794
rect 9422 10767 9423 10793
rect 9423 10767 9449 10793
rect 9449 10767 9450 10793
rect 9422 10766 9450 10767
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 9926 11662 9954 11690
rect 9870 11494 9898 11522
rect 10710 11158 10738 11186
rect 9758 11046 9786 11074
rect 9086 10710 9114 10738
rect 9030 10206 9058 10234
rect 9198 10206 9226 10234
rect 9086 10038 9114 10066
rect 9702 10038 9730 10066
rect 9478 10009 9506 10010
rect 9478 9983 9479 10009
rect 9479 9983 9505 10009
rect 9505 9983 9506 10009
rect 9478 9982 9506 9983
rect 9254 9702 9282 9730
rect 9310 9926 9338 9954
rect 9646 9953 9674 9954
rect 9646 9927 9647 9953
rect 9647 9927 9673 9953
rect 9673 9927 9674 9953
rect 9646 9926 9674 9927
rect 8750 9505 8778 9506
rect 8750 9479 8751 9505
rect 8751 9479 8777 9505
rect 8777 9479 8778 9505
rect 8750 9478 8778 9479
rect 9030 9478 9058 9506
rect 8694 9198 8722 9226
rect 8302 8862 8330 8890
rect 7350 8414 7378 8442
rect 7518 8385 7546 8386
rect 7518 8359 7519 8385
rect 7519 8359 7545 8385
rect 7545 8359 7546 8385
rect 7518 8358 7546 8359
rect 8134 8385 8162 8386
rect 8134 8359 8135 8385
rect 8135 8359 8161 8385
rect 8161 8359 8162 8385
rect 8134 8358 8162 8359
rect 7070 8022 7098 8050
rect 8190 8049 8218 8050
rect 8190 8023 8191 8049
rect 8191 8023 8217 8049
rect 8217 8023 8218 8049
rect 8190 8022 8218 8023
rect 8302 8414 8330 8442
rect 9422 9310 9450 9338
rect 9702 9310 9730 9338
rect 10262 11046 10290 11074
rect 9814 10934 9842 10962
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 9870 10878 9898 10906
rect 10038 10401 10066 10402
rect 10038 10375 10039 10401
rect 10039 10375 10065 10401
rect 10065 10375 10066 10401
rect 10038 10374 10066 10375
rect 10262 10262 10290 10290
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9982 10038 10010 10066
rect 10878 10766 10906 10794
rect 10654 10289 10682 10290
rect 10654 10263 10655 10289
rect 10655 10263 10681 10289
rect 10681 10263 10682 10289
rect 10654 10262 10682 10263
rect 10710 10065 10738 10066
rect 10710 10039 10711 10065
rect 10711 10039 10737 10065
rect 10737 10039 10738 10065
rect 10710 10038 10738 10039
rect 10486 9926 10514 9954
rect 10318 9814 10346 9842
rect 10710 9814 10738 9842
rect 10262 9729 10290 9730
rect 10262 9703 10263 9729
rect 10263 9703 10289 9729
rect 10289 9703 10290 9729
rect 10262 9702 10290 9703
rect 9870 9534 9898 9562
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9478 9281 9506 9282
rect 9478 9255 9479 9281
rect 9479 9255 9505 9281
rect 9505 9255 9506 9281
rect 9478 9254 9506 9255
rect 9422 9198 9450 9226
rect 9590 9225 9618 9226
rect 9590 9199 9591 9225
rect 9591 9199 9617 9225
rect 9617 9199 9618 9225
rect 9590 9198 9618 9199
rect 10038 9281 10066 9282
rect 10038 9255 10039 9281
rect 10039 9255 10065 9281
rect 10065 9255 10066 9281
rect 10038 9254 10066 9255
rect 10206 9617 10234 9618
rect 10206 9591 10207 9617
rect 10207 9591 10233 9617
rect 10233 9591 10234 9617
rect 10206 9590 10234 9591
rect 10150 9561 10178 9562
rect 10150 9535 10151 9561
rect 10151 9535 10177 9561
rect 10177 9535 10178 9561
rect 10150 9534 10178 9535
rect 10318 9254 10346 9282
rect 9198 8414 9226 8442
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 9646 8526 9674 8554
rect 10150 8553 10178 8554
rect 10150 8527 10151 8553
rect 10151 8527 10177 8553
rect 10177 8527 10178 8553
rect 10150 8526 10178 8527
rect 10262 8526 10290 8554
rect 10766 8638 10794 8666
rect 11214 11830 11242 11858
rect 13342 13230 13370 13258
rect 12390 13174 12418 13202
rect 13286 13201 13314 13202
rect 13286 13175 13287 13201
rect 13287 13175 13313 13201
rect 13313 13175 13314 13201
rect 13286 13174 13314 13175
rect 11942 12361 11970 12362
rect 11942 12335 11943 12361
rect 11943 12335 11969 12361
rect 11969 12335 11970 12361
rect 11942 12334 11970 12335
rect 11494 11774 11522 11802
rect 11886 11633 11914 11634
rect 11886 11607 11887 11633
rect 11887 11607 11913 11633
rect 11913 11607 11914 11633
rect 11886 11606 11914 11607
rect 11662 10401 11690 10402
rect 11662 10375 11663 10401
rect 11663 10375 11689 10401
rect 11689 10375 11690 10401
rect 11662 10374 11690 10375
rect 11158 9310 11186 9338
rect 12334 11606 12362 11634
rect 12614 11046 12642 11074
rect 13062 11998 13090 12026
rect 14070 13118 14098 13146
rect 14014 12726 14042 12754
rect 13286 12025 13314 12026
rect 13286 11999 13287 12025
rect 13287 11999 13313 12025
rect 13313 11999 13314 12025
rect 13286 11998 13314 11999
rect 13454 11942 13482 11970
rect 13678 11969 13706 11970
rect 13678 11943 13679 11969
rect 13679 11943 13705 11969
rect 13705 11943 13706 11969
rect 13678 11942 13706 11943
rect 12726 11886 12754 11914
rect 13230 11913 13258 11914
rect 13230 11887 13231 11913
rect 13231 11887 13257 11913
rect 13257 11887 13258 11913
rect 13230 11886 13258 11887
rect 12838 11830 12866 11858
rect 12726 10990 12754 11018
rect 11326 9310 11354 9338
rect 12782 10766 12810 10794
rect 12726 10710 12754 10738
rect 18830 13145 18858 13146
rect 18830 13119 18831 13145
rect 18831 13119 18857 13145
rect 18857 13119 18858 13145
rect 18830 13118 18858 13119
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 19950 12782 19978 12810
rect 18830 12753 18858 12754
rect 18830 12727 18831 12753
rect 18831 12727 18857 12753
rect 18857 12727 18858 12753
rect 18830 12726 18858 12727
rect 20006 12446 20034 12474
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 13286 11830 13314 11858
rect 12894 11774 12922 11802
rect 13230 11774 13258 11802
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 13118 11073 13146 11074
rect 13118 11047 13119 11073
rect 13119 11047 13145 11073
rect 13145 11047 13146 11073
rect 13118 11046 13146 11047
rect 12670 9926 12698 9954
rect 11998 9590 12026 9618
rect 12222 9617 12250 9618
rect 12222 9591 12223 9617
rect 12223 9591 12249 9617
rect 12249 9591 12250 9617
rect 12222 9590 12250 9591
rect 12390 9505 12418 9506
rect 12390 9479 12391 9505
rect 12391 9479 12417 9505
rect 12417 9479 12418 9505
rect 12390 9478 12418 9479
rect 11270 9254 11298 9282
rect 11718 9281 11746 9282
rect 11718 9255 11719 9281
rect 11719 9255 11745 9281
rect 11745 9255 11746 9281
rect 11718 9254 11746 9255
rect 11438 9225 11466 9226
rect 11438 9199 11439 9225
rect 11439 9199 11465 9225
rect 11465 9199 11466 9225
rect 11438 9198 11466 9199
rect 10934 8638 10962 8666
rect 11102 8638 11130 8666
rect 10766 8526 10794 8554
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 11886 9281 11914 9282
rect 11886 9255 11887 9281
rect 11887 9255 11913 9281
rect 11913 9255 11914 9281
rect 11886 9254 11914 9255
rect 11774 9198 11802 9226
rect 11550 9113 11578 9114
rect 11550 9087 11551 9113
rect 11551 9087 11577 9113
rect 11577 9087 11578 9113
rect 11550 9086 11578 9087
rect 12054 9113 12082 9114
rect 12054 9087 12055 9113
rect 12055 9087 12081 9113
rect 12081 9087 12082 9113
rect 12054 9086 12082 9087
rect 13006 10766 13034 10794
rect 12838 9870 12866 9898
rect 12782 9337 12810 9338
rect 12782 9311 12783 9337
rect 12783 9311 12809 9337
rect 12809 9311 12810 9337
rect 12782 9310 12810 9311
rect 12670 9281 12698 9282
rect 12670 9255 12671 9281
rect 12671 9255 12697 9281
rect 12697 9255 12698 9281
rect 12670 9254 12698 9255
rect 12166 8918 12194 8946
rect 12334 8638 12362 8666
rect 12614 8638 12642 8666
rect 11438 8526 11466 8554
rect 14854 10849 14882 10850
rect 14854 10823 14855 10849
rect 14855 10823 14881 10849
rect 14881 10823 14882 10849
rect 14854 10822 14882 10823
rect 14518 10737 14546 10738
rect 14518 10711 14519 10737
rect 14519 10711 14545 10737
rect 14545 10711 14546 10737
rect 14518 10710 14546 10711
rect 14742 10710 14770 10738
rect 20006 11774 20034 11802
rect 18830 11577 18858 11578
rect 18830 11551 18831 11577
rect 18831 11551 18857 11577
rect 18857 11551 18858 11577
rect 18830 11550 18858 11551
rect 20006 11465 20034 11466
rect 20006 11439 20007 11465
rect 20007 11439 20033 11465
rect 20033 11439 20034 11465
rect 20006 11438 20034 11439
rect 18774 10822 18802 10850
rect 15190 10766 15218 10794
rect 18830 10793 18858 10794
rect 18830 10767 18831 10793
rect 18831 10767 18857 10793
rect 18857 10767 18858 10793
rect 18830 10766 18858 10767
rect 15078 10710 15106 10738
rect 20006 11102 20034 11130
rect 18942 10710 18970 10738
rect 20006 10766 20034 10794
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 20006 10457 20034 10458
rect 20006 10431 20007 10457
rect 20007 10431 20033 10457
rect 20033 10431 20034 10457
rect 20006 10430 20034 10431
rect 14462 10150 14490 10178
rect 14742 10289 14770 10290
rect 14742 10263 14743 10289
rect 14743 10263 14769 10289
rect 14769 10263 14770 10289
rect 14742 10262 14770 10263
rect 13230 9953 13258 9954
rect 13230 9927 13231 9953
rect 13231 9927 13257 9953
rect 13257 9927 13258 9953
rect 13230 9926 13258 9927
rect 13734 10038 13762 10066
rect 13790 9982 13818 10010
rect 14462 10009 14490 10010
rect 14462 9983 14463 10009
rect 14463 9983 14489 10009
rect 14489 9983 14490 10009
rect 14462 9982 14490 9983
rect 18830 10401 18858 10402
rect 18830 10375 18831 10401
rect 18831 10375 18857 10401
rect 18857 10375 18858 10401
rect 18830 10374 18858 10375
rect 14966 9982 14994 10010
rect 14518 9897 14546 9898
rect 14518 9871 14519 9897
rect 14519 9871 14545 9897
rect 14545 9871 14546 9897
rect 14518 9870 14546 9871
rect 20006 10038 20034 10066
rect 18830 10009 18858 10010
rect 18830 9983 18831 10009
rect 18831 9983 18857 10009
rect 18857 9983 18858 10009
rect 18830 9982 18858 9983
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 20006 9758 20034 9786
rect 13118 9366 13146 9394
rect 13678 9478 13706 9506
rect 13230 9337 13258 9338
rect 13230 9311 13231 9337
rect 13231 9311 13257 9337
rect 13257 9311 13258 9337
rect 13230 9310 13258 9311
rect 13006 9225 13034 9226
rect 13006 9199 13007 9225
rect 13007 9199 13033 9225
rect 13033 9199 13034 9225
rect 13006 9198 13034 9199
rect 13454 9225 13482 9226
rect 13454 9199 13455 9225
rect 13455 9199 13481 9225
rect 13481 9199 13482 9225
rect 13454 9198 13482 9199
rect 12894 8638 12922 8666
rect 13510 9142 13538 9170
rect 13790 9225 13818 9226
rect 13790 9199 13791 9225
rect 13791 9199 13817 9225
rect 13817 9199 13818 9225
rect 13790 9198 13818 9199
rect 13790 8889 13818 8890
rect 13790 8863 13791 8889
rect 13791 8863 13817 8889
rect 13817 8863 13818 8889
rect 13790 8862 13818 8863
rect 15078 9590 15106 9618
rect 18830 9617 18858 9618
rect 18830 9591 18831 9617
rect 18831 9591 18857 9617
rect 18857 9591 18858 9617
rect 18830 9590 18858 9591
rect 20006 9422 20034 9450
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 18830 8918 18858 8946
rect 19950 9086 19978 9114
rect 18942 8862 18970 8890
rect 14070 8806 14098 8834
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 19670 8750 19698 8778
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 20118 2366 20146 2394
rect 10022 2338 10050 2339
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 8414 1694 8442 1722
rect 9030 1694 9058 1722
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 11433 19110 11438 19138
rect 11466 19110 12782 19138
rect 12810 19110 12815 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 10761 18718 10766 18746
rect 10794 18718 11382 18746
rect 11410 18718 11415 18746
rect 12105 18718 12110 18746
rect 12138 18718 13118 18746
rect 13146 18718 13151 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 0 18186 400 18200
rect 0 18158 854 18186
rect 882 18158 887 18186
rect 0 18144 400 18158
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 10761 14014 10766 14042
rect 10794 14014 11102 14042
rect 11130 14014 11135 14042
rect 10145 13790 10150 13818
rect 10178 13790 10766 13818
rect 10794 13790 10799 13818
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 11265 13454 11270 13482
rect 11298 13454 12278 13482
rect 12306 13454 12311 13482
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 10817 13230 10822 13258
rect 10850 13230 11998 13258
rect 12026 13230 13342 13258
rect 13370 13230 13375 13258
rect 11937 13174 11942 13202
rect 11970 13174 12390 13202
rect 12418 13174 12423 13202
rect 13281 13174 13286 13202
rect 13314 13174 13454 13202
rect 0 13146 400 13160
rect 13426 13146 13454 13174
rect 0 13118 8750 13146
rect 8778 13118 8783 13146
rect 13426 13118 14070 13146
rect 14098 13118 18830 13146
rect 18858 13118 18863 13146
rect 0 13104 400 13118
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 20600 12810 21000 12824
rect 19945 12782 19950 12810
rect 19978 12782 21000 12810
rect 20600 12768 21000 12782
rect 14009 12726 14014 12754
rect 14042 12726 18830 12754
rect 18858 12726 18863 12754
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 0 12474 400 12488
rect 20600 12474 21000 12488
rect 0 12446 966 12474
rect 994 12446 999 12474
rect 8521 12446 8526 12474
rect 8554 12446 9646 12474
rect 9674 12446 9679 12474
rect 20001 12446 20006 12474
rect 20034 12446 21000 12474
rect 0 12432 400 12446
rect 20600 12432 21000 12446
rect 7546 12390 8358 12418
rect 8386 12390 8391 12418
rect 9081 12390 9086 12418
rect 9114 12390 9758 12418
rect 9786 12390 9791 12418
rect 7546 12306 7574 12390
rect 7905 12334 7910 12362
rect 7938 12334 8246 12362
rect 8274 12334 8279 12362
rect 8409 12334 8414 12362
rect 8442 12334 11942 12362
rect 11970 12334 11975 12362
rect 2137 12278 2142 12306
rect 2170 12278 6678 12306
rect 6706 12278 7574 12306
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 13057 11998 13062 12026
rect 13090 11998 13286 12026
rect 13314 11998 13319 12026
rect 7681 11942 7686 11970
rect 7714 11942 8246 11970
rect 8274 11942 10010 11970
rect 13449 11942 13454 11970
rect 13482 11942 13678 11970
rect 13706 11942 13711 11970
rect 9982 11914 10010 11942
rect 9137 11886 9142 11914
rect 9170 11886 9954 11914
rect 9982 11886 12726 11914
rect 12754 11886 13230 11914
rect 13258 11886 13263 11914
rect 9926 11858 9954 11886
rect 9081 11830 9086 11858
rect 9114 11830 9366 11858
rect 9394 11830 9399 11858
rect 9921 11830 9926 11858
rect 9954 11830 11214 11858
rect 11242 11830 11247 11858
rect 12833 11830 12838 11858
rect 12866 11830 13286 11858
rect 13314 11830 13319 11858
rect 20600 11802 21000 11816
rect 9137 11774 9142 11802
rect 9170 11774 9478 11802
rect 9506 11774 9511 11802
rect 10094 11774 11494 11802
rect 11522 11774 12894 11802
rect 12922 11774 13230 11802
rect 13258 11774 13263 11802
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 9305 11718 9310 11746
rect 9338 11718 9758 11746
rect 9786 11718 9791 11746
rect 10094 11690 10122 11774
rect 20600 11760 21000 11774
rect 9921 11662 9926 11690
rect 9954 11662 10122 11690
rect 11881 11606 11886 11634
rect 11914 11606 12334 11634
rect 12362 11606 15974 11634
rect 15946 11578 15974 11606
rect 8129 11550 8134 11578
rect 8162 11550 9422 11578
rect 9450 11550 9455 11578
rect 15946 11550 18830 11578
rect 18858 11550 18863 11578
rect 9697 11494 9702 11522
rect 9730 11494 9870 11522
rect 9898 11494 9903 11522
rect 20600 11466 21000 11480
rect 20001 11438 20006 11466
rect 20034 11438 21000 11466
rect 20600 11424 21000 11438
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 7499 11270 7518 11298
rect 7546 11270 7551 11298
rect 961 11214 966 11242
rect 994 11214 999 11242
rect 8745 11214 8750 11242
rect 8778 11214 9702 11242
rect 9730 11214 9735 11242
rect 0 11130 400 11144
rect 966 11130 994 11214
rect 2137 11158 2142 11186
rect 2170 11158 5950 11186
rect 5978 11158 7518 11186
rect 7546 11158 7551 11186
rect 9305 11158 9310 11186
rect 9338 11158 10710 11186
rect 10738 11158 10743 11186
rect 20600 11130 21000 11144
rect 0 11102 994 11130
rect 7401 11102 7406 11130
rect 7434 11102 7686 11130
rect 7714 11102 7719 11130
rect 8969 11102 8974 11130
rect 9002 11102 9198 11130
rect 9226 11102 9231 11130
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 0 11088 400 11102
rect 20600 11088 21000 11102
rect 9753 11046 9758 11074
rect 9786 11046 10262 11074
rect 10290 11046 10295 11074
rect 12609 11046 12614 11074
rect 12642 11046 13118 11074
rect 13146 11046 13151 11074
rect 8801 10990 8806 11018
rect 8834 10990 9086 11018
rect 9114 10990 9119 11018
rect 12707 10990 12726 11018
rect 12754 10990 12759 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 7849 10934 7854 10962
rect 7882 10934 8078 10962
rect 8106 10934 8111 10962
rect 8857 10934 8862 10962
rect 8890 10934 9814 10962
rect 9842 10934 9847 10962
rect 7345 10878 7350 10906
rect 7378 10878 7518 10906
rect 7546 10878 8190 10906
rect 8218 10878 8223 10906
rect 9137 10878 9142 10906
rect 9170 10878 9870 10906
rect 9898 10878 9903 10906
rect 7737 10822 7742 10850
rect 7770 10822 8134 10850
rect 8162 10822 8167 10850
rect 8297 10822 8302 10850
rect 8330 10822 9198 10850
rect 9226 10822 9231 10850
rect 14849 10822 14854 10850
rect 14882 10822 18774 10850
rect 18802 10822 18807 10850
rect 0 10794 400 10808
rect 20600 10794 21000 10808
rect 0 10766 994 10794
rect 6449 10766 6454 10794
rect 6482 10766 7182 10794
rect 7210 10766 7406 10794
rect 7434 10766 7966 10794
rect 7994 10766 9254 10794
rect 9282 10766 9287 10794
rect 9417 10766 9422 10794
rect 9450 10766 10878 10794
rect 10906 10766 10911 10794
rect 12777 10766 12782 10794
rect 12810 10766 13006 10794
rect 13034 10766 13039 10794
rect 15185 10766 15190 10794
rect 15218 10766 18830 10794
rect 18858 10766 18863 10794
rect 20001 10766 20006 10794
rect 20034 10766 21000 10794
rect 0 10752 400 10766
rect 966 10738 994 10766
rect 20600 10752 21000 10766
rect 961 10710 966 10738
rect 994 10710 999 10738
rect 7854 10710 9086 10738
rect 9114 10710 9119 10738
rect 12707 10710 12726 10738
rect 12754 10710 12759 10738
rect 14513 10710 14518 10738
rect 14546 10710 14742 10738
rect 14770 10710 15078 10738
rect 15106 10710 18942 10738
rect 18970 10710 18975 10738
rect 7854 10626 7882 10710
rect 7121 10598 7126 10626
rect 7154 10598 7854 10626
rect 7882 10598 7887 10626
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 2137 10486 2142 10514
rect 2170 10486 6734 10514
rect 6762 10486 6767 10514
rect 0 10458 400 10472
rect 20600 10458 21000 10472
rect 0 10430 966 10458
rect 994 10430 999 10458
rect 20001 10430 20006 10458
rect 20034 10430 21000 10458
rect 0 10416 400 10430
rect 20600 10416 21000 10430
rect 2137 10374 2142 10402
rect 2170 10374 4998 10402
rect 5026 10374 6846 10402
rect 6874 10374 7126 10402
rect 7154 10374 7159 10402
rect 10033 10374 10038 10402
rect 10066 10374 11662 10402
rect 11690 10374 11695 10402
rect 15946 10374 18830 10402
rect 18858 10374 18863 10402
rect 15946 10290 15974 10374
rect 10257 10262 10262 10290
rect 10290 10262 10654 10290
rect 10682 10262 10687 10290
rect 14737 10262 14742 10290
rect 14770 10262 15974 10290
rect 9025 10206 9030 10234
rect 9058 10206 9198 10234
rect 9226 10206 9231 10234
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 6897 10150 6902 10178
rect 6930 10150 7294 10178
rect 7322 10150 7327 10178
rect 14457 10150 14462 10178
rect 14490 10150 14495 10178
rect 14462 10066 14490 10150
rect 20600 10122 21000 10136
rect 20006 10094 21000 10122
rect 20006 10066 20034 10094
rect 20600 10080 21000 10094
rect 6057 10038 6062 10066
rect 6090 10038 6790 10066
rect 6818 10038 6823 10066
rect 7345 10038 7350 10066
rect 7378 10038 7574 10066
rect 7602 10038 7607 10066
rect 8353 10038 8358 10066
rect 8386 10038 8862 10066
rect 8890 10038 8895 10066
rect 9081 10038 9086 10066
rect 9114 10038 9702 10066
rect 9730 10038 9982 10066
rect 10010 10038 10710 10066
rect 10738 10038 10743 10066
rect 13729 10038 13734 10066
rect 13762 10038 14490 10066
rect 20001 10038 20006 10066
rect 20034 10038 20039 10066
rect 2137 9982 2142 10010
rect 2170 9982 5614 10010
rect 5642 9982 7126 10010
rect 7154 9982 7159 10010
rect 7457 9982 7462 10010
rect 7490 9982 9478 10010
rect 9506 9982 9511 10010
rect 13785 9982 13790 10010
rect 13818 9982 14462 10010
rect 14490 9982 14495 10010
rect 14961 9982 14966 10010
rect 14994 9982 18830 10010
rect 18858 9982 18863 10010
rect 6729 9926 6734 9954
rect 6762 9926 7406 9954
rect 7434 9926 7742 9954
rect 7770 9926 7775 9954
rect 9305 9926 9310 9954
rect 9338 9926 9646 9954
rect 9674 9926 10486 9954
rect 10514 9926 10519 9954
rect 12665 9926 12670 9954
rect 12698 9926 13230 9954
rect 13258 9926 13263 9954
rect 961 9870 966 9898
rect 994 9870 999 9898
rect 7233 9870 7238 9898
rect 7266 9870 7350 9898
rect 7378 9870 8862 9898
rect 8890 9870 8895 9898
rect 12833 9870 12838 9898
rect 12866 9870 14518 9898
rect 14546 9870 14551 9898
rect 0 9786 400 9800
rect 966 9786 994 9870
rect 8633 9814 8638 9842
rect 8666 9814 10318 9842
rect 10346 9814 10710 9842
rect 10738 9814 10743 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 20600 9786 21000 9800
rect 0 9758 994 9786
rect 20001 9758 20006 9786
rect 20034 9758 21000 9786
rect 0 9744 400 9758
rect 20600 9744 21000 9758
rect 9249 9702 9254 9730
rect 9282 9702 10262 9730
rect 10290 9702 10295 9730
rect 6897 9590 6902 9618
rect 6930 9590 7294 9618
rect 7322 9590 7327 9618
rect 10201 9590 10206 9618
rect 10234 9590 11998 9618
rect 12026 9590 12222 9618
rect 12250 9590 12255 9618
rect 15073 9590 15078 9618
rect 15106 9590 18830 9618
rect 18858 9590 18863 9618
rect 9865 9534 9870 9562
rect 9898 9534 10150 9562
rect 10178 9534 10183 9562
rect 8073 9478 8078 9506
rect 8106 9478 8750 9506
rect 8778 9478 9030 9506
rect 9058 9478 9063 9506
rect 12385 9478 12390 9506
rect 12418 9478 13678 9506
rect 13706 9478 13711 9506
rect 20600 9450 21000 9464
rect 20001 9422 20006 9450
rect 20034 9422 21000 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 20600 9408 21000 9422
rect 11046 9366 13118 9394
rect 13146 9366 13151 9394
rect 11046 9338 11074 9366
rect 9417 9310 9422 9338
rect 9450 9310 9702 9338
rect 9730 9310 11074 9338
rect 11153 9310 11158 9338
rect 11186 9310 11326 9338
rect 11354 9310 12782 9338
rect 12810 9310 13230 9338
rect 13258 9310 13263 9338
rect 8353 9254 8358 9282
rect 8386 9254 9478 9282
rect 9506 9254 10038 9282
rect 10066 9254 10071 9282
rect 10313 9254 10318 9282
rect 10346 9254 11270 9282
rect 11298 9254 11718 9282
rect 11746 9254 11751 9282
rect 11881 9254 11886 9282
rect 11914 9254 12670 9282
rect 12698 9254 12703 9282
rect 8689 9198 8694 9226
rect 8722 9198 9422 9226
rect 9450 9198 9590 9226
rect 9618 9198 9623 9226
rect 11433 9198 11438 9226
rect 11466 9198 11774 9226
rect 11802 9198 11807 9226
rect 13001 9198 13006 9226
rect 13034 9198 13039 9226
rect 13449 9198 13454 9226
rect 13482 9198 13790 9226
rect 13818 9198 13823 9226
rect 13006 9170 13034 9198
rect 13006 9142 13510 9170
rect 13538 9142 13543 9170
rect 20600 9114 21000 9128
rect 11545 9086 11550 9114
rect 11578 9086 12054 9114
rect 12082 9086 12087 9114
rect 19945 9086 19950 9114
rect 19978 9086 21000 9114
rect 20600 9072 21000 9086
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 12161 8918 12166 8946
rect 12194 8918 18830 8946
rect 18858 8918 18863 8946
rect 961 8862 966 8890
rect 994 8862 999 8890
rect 7009 8862 7014 8890
rect 7042 8862 8302 8890
rect 8330 8862 8335 8890
rect 13785 8862 13790 8890
rect 13818 8862 18942 8890
rect 18970 8862 18975 8890
rect 0 8778 400 8792
rect 966 8778 994 8862
rect 2137 8806 2142 8834
rect 2170 8806 5670 8834
rect 5698 8806 7294 8834
rect 7322 8806 7462 8834
rect 7490 8806 7495 8834
rect 14065 8806 14070 8834
rect 14098 8806 18830 8834
rect 18858 8806 18863 8834
rect 20600 8778 21000 8792
rect 0 8750 994 8778
rect 19665 8750 19670 8778
rect 19698 8750 21000 8778
rect 0 8736 400 8750
rect 20600 8736 21000 8750
rect 6841 8694 6846 8722
rect 6874 8694 7126 8722
rect 7154 8694 7159 8722
rect 10761 8638 10766 8666
rect 10794 8638 10934 8666
rect 10962 8638 11102 8666
rect 11130 8638 12334 8666
rect 12362 8638 12614 8666
rect 12642 8638 12894 8666
rect 12922 8638 12927 8666
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 9641 8526 9646 8554
rect 9674 8526 10150 8554
rect 10178 8526 10183 8554
rect 10257 8526 10262 8554
rect 10290 8526 10766 8554
rect 10794 8526 11438 8554
rect 11466 8526 11471 8554
rect 0 8442 400 8456
rect 0 8414 966 8442
rect 994 8414 999 8442
rect 2137 8414 2142 8442
rect 2170 8414 7350 8442
rect 7378 8414 7383 8442
rect 8297 8414 8302 8442
rect 8330 8414 9198 8442
rect 9226 8414 9231 8442
rect 0 8400 400 8414
rect 7513 8358 7518 8386
rect 7546 8358 8134 8386
rect 8162 8358 8167 8386
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 6841 8022 6846 8050
rect 6874 8022 7070 8050
rect 7098 8022 8190 8050
rect 8218 8022 8223 8050
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 20600 2394 21000 2408
rect 20113 2366 20118 2394
rect 20146 2366 21000 2394
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 20600 2352 21000 2366
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 8409 1694 8414 1722
rect 8442 1694 9030 1722
rect 9058 1694 9063 1722
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 7518 11270 7546 11298
rect 12726 10990 12754 11018
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 7518 10878 7546 10906
rect 12726 10710 12754 10738
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 7518 11298 7546 11303
rect 7518 10906 7546 11270
rect 7518 10873 7546 10878
rect 9904 10990 10064 11746
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 10206 10064 10962
rect 12726 11018 12754 11023
rect 12726 10738 12754 10990
rect 12726 10705 12754 10710
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _072_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9744 0 -1 8624
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _073_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9184 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _074_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9240 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _075_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9128 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _076_
timestamp 1698175906
transform 1 0 9240 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _077_
timestamp 1698175906
transform -1 0 9912 0 -1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _078_
timestamp 1698175906
transform 1 0 10192 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _079_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9744 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _080_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8512 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _081_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9464 0 -1 10192
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _082_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8512 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _083_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9464 0 -1 10192
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _084_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7056 0 -1 10192
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _085_
timestamp 1698175906
transform 1 0 9016 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _086_
timestamp 1698175906
transform -1 0 8008 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _087_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _088_
timestamp 1698175906
transform 1 0 8008 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _089_
timestamp 1698175906
transform 1 0 13608 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _090_
timestamp 1698175906
transform 1 0 13160 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _091_
timestamp 1698175906
transform -1 0 8512 0 -1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _092_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8400 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _093_
timestamp 1698175906
transform -1 0 7896 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _094_
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _095_
timestamp 1698175906
transform 1 0 12152 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _096_
timestamp 1698175906
transform 1 0 14392 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _097_
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _098_
timestamp 1698175906
transform -1 0 13888 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _099_
timestamp 1698175906
transform 1 0 13048 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _100_
timestamp 1698175906
transform -1 0 10920 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _101_
timestamp 1698175906
transform -1 0 10024 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _102_
timestamp 1698175906
transform -1 0 14056 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _103_
timestamp 1698175906
transform 1 0 13048 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _104_
timestamp 1698175906
transform -1 0 13776 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _105_
timestamp 1698175906
transform 1 0 12600 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _106_
timestamp 1698175906
transform -1 0 12040 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _107_
timestamp 1698175906
transform 1 0 11144 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _108_
timestamp 1698175906
transform -1 0 8960 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8960 0 1 9408
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _110_
timestamp 1698175906
transform -1 0 7448 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _111_
timestamp 1698175906
transform -1 0 7280 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8512 0 -1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _113_
timestamp 1698175906
transform -1 0 7616 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7056 0 1 10192
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _115_
timestamp 1698175906
transform -1 0 6944 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _116_
timestamp 1698175906
transform -1 0 7952 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7336 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _118_
timestamp 1698175906
transform -1 0 7336 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _119_
timestamp 1698175906
transform 1 0 9744 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10024 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform 1 0 10080 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _122_
timestamp 1698175906
transform 1 0 9016 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10024 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1698175906
transform 1 0 10248 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _125_
timestamp 1698175906
transform 1 0 10584 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform 1 0 10808 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _127_
timestamp 1698175906
transform -1 0 10808 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _128_
timestamp 1698175906
transform -1 0 10360 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_
timestamp 1698175906
transform -1 0 12152 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _130_
timestamp 1698175906
transform -1 0 12208 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _131_
timestamp 1698175906
transform -1 0 11648 0 -1 9408
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform -1 0 9632 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _133_
timestamp 1698175906
transform -1 0 9128 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _134_
timestamp 1698175906
transform 1 0 8680 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _135_
timestamp 1698175906
transform -1 0 10192 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _136_
timestamp 1698175906
transform 1 0 9688 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1698175906
transform -1 0 12096 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform -1 0 12096 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _139_
timestamp 1698175906
transform 1 0 11312 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _140_
timestamp 1698175906
transform 1 0 11648 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _141_
timestamp 1698175906
transform -1 0 13440 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _142_
timestamp 1698175906
transform 1 0 12712 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _143_
timestamp 1698175906
transform -1 0 9688 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _144_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10640 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _145_
timestamp 1698175906
transform 1 0 10864 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _146_
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _147_
timestamp 1698175906
transform -1 0 11256 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _148_
timestamp 1698175906
transform 1 0 8120 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _149_
timestamp 1698175906
transform 1 0 8064 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _150_
timestamp 1698175906
transform 1 0 9240 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _151_
timestamp 1698175906
transform -1 0 7168 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _152_
timestamp 1698175906
transform 1 0 12488 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _153_
timestamp 1698175906
transform -1 0 8232 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _154_
timestamp 1698175906
transform 1 0 12768 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _155_
timestamp 1698175906
transform 1 0 12992 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _156_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9296 0 -1 13328
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _157_
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _158_
timestamp 1698175906
transform 1 0 12264 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _159_
timestamp 1698175906
transform 1 0 10808 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _160_
timestamp 1698175906
transform -1 0 7224 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _161_
timestamp 1698175906
transform 1 0 6776 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _162_
timestamp 1698175906
transform -1 0 6552 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _163_
timestamp 1698175906
transform -1 0 7504 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _166_
timestamp 1698175906
transform 1 0 14616 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _167_
timestamp 1698175906
transform 1 0 11032 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _168_
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _169_
timestamp 1698175906
transform -1 0 7616 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _170_
timestamp 1698175906
transform -1 0 7000 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _171_
timestamp 1698175906
transform 1 0 14840 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _172_
timestamp 1698175906
transform -1 0 11032 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _173_
timestamp 1698175906
transform 1 0 14952 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8736 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9632 0 -1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 11592 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_165 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9912 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698175906
transform 1 0 10136 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 12208 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 16128 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_317 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_333 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19320 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_341
timestamp 1698175906
transform 1 0 19768 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 10248 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698175906
transform 1 0 12208 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698175906
transform 1 0 10248 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 14168 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_104
timestamp 1698175906
transform 1 0 6496 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_108
timestamp 1698175906
transform 1 0 6720 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698175906
transform 1 0 8400 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_152
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_189
timestamp 1698175906
transform 1 0 11256 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_205
timestamp 1698175906
transform 1 0 12152 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 12376 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 16128 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_123
timestamp 1698175906
transform 1 0 7560 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_131
timestamp 1698175906
transform 1 0 8008 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_162
timestamp 1698175906
transform 1 0 9744 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_170
timestamp 1698175906
transform 1 0 10192 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 10416 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_177
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698175906
transform 1 0 14168 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 2240 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 4032 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 4480 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_117
timestamp 1698175906
transform 1 0 7224 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_124
timestamp 1698175906
transform 1 0 7616 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_128
timestamp 1698175906
transform 1 0 7840 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_174
timestamp 1698175906
transform 1 0 10416 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698175906
transform 1 0 12208 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_241
timestamp 1698175906
transform 1 0 14168 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_273
timestamp 1698175906
transform 1 0 15960 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698175906
transform 1 0 16184 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 16296 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_109
timestamp 1698175906
transform 1 0 6776 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_124
timestamp 1698175906
transform 1 0 7616 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_140
timestamp 1698175906
transform 1 0 8512 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_148
timestamp 1698175906
transform 1 0 8960 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_152
timestamp 1698175906
transform 1 0 9184 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_154
timestamp 1698175906
transform 1 0 9296 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_161
timestamp 1698175906
transform 1 0 9688 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_165
timestamp 1698175906
transform 1 0 9912 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698175906
transform 1 0 10248 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_177
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_236
timestamp 1698175906
transform 1 0 13888 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 14336 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_80
timestamp 1698175906
transform 1 0 5152 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_84
timestamp 1698175906
transform 1 0 5376 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_86
timestamp 1698175906
transform 1 0 5488 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_121
timestamp 1698175906
transform 1 0 7448 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_137
timestamp 1698175906
transform 1 0 8344 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 8456 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_150
timestamp 1698175906
transform 1 0 9072 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_154
timestamp 1698175906
transform 1 0 9296 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_164
timestamp 1698175906
transform 1 0 9856 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_170
timestamp 1698175906
transform 1 0 10192 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_178
timestamp 1698175906
transform 1 0 10640 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_182
timestamp 1698175906
transform 1 0 10864 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_184
timestamp 1698175906
transform 1 0 10976 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698175906
transform 1 0 12208 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_239
timestamp 1698175906
transform 1 0 14056 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_271
timestamp 1698175906
transform 1 0 15848 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 16296 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 18256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 18704 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_113
timestamp 1698175906
transform 1 0 7000 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_129
timestamp 1698175906
transform 1 0 7896 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_133
timestamp 1698175906
transform 1 0 8120 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698175906
transform 1 0 10360 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_177
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_193
timestamp 1698175906
transform 1 0 11480 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_201
timestamp 1698175906
transform 1 0 11928 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_211
timestamp 1698175906
transform 1 0 12488 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_227
timestamp 1698175906
transform 1 0 13384 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_236
timestamp 1698175906
transform 1 0 13888 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 14336 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 2240 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 4032 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 4480 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_104
timestamp 1698175906
transform 1 0 6496 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_112
timestamp 1698175906
transform 1 0 6944 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_123
timestamp 1698175906
transform 1 0 7560 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_131
timestamp 1698175906
transform 1 0 8008 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_135
timestamp 1698175906
transform 1 0 8232 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_182
timestamp 1698175906
transform 1 0 10864 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_198
timestamp 1698175906
transform 1 0 11760 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_205
timestamp 1698175906
transform 1 0 12152 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 12376 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_212
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_250
timestamp 1698175906
transform 1 0 14672 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_266
timestamp 1698175906
transform 1 0 15568 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_274
timestamp 1698175906
transform 1 0 16016 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 16240 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 18256 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 18704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698175906
transform 1 0 2240 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698175906
transform 1 0 2464 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 4536 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 4760 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 4872 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_113
timestamp 1698175906
transform 1 0 7000 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_259
timestamp 1698175906
transform 1 0 15176 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_291
timestamp 1698175906
transform 1 0 16968 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_307
timestamp 1698175906
transform 1 0 17864 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 18648 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 2240 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 4032 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 4480 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_88
timestamp 1698175906
transform 1 0 5600 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_92
timestamp 1698175906
transform 1 0 5824 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_122
timestamp 1698175906
transform 1 0 7504 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_138
timestamp 1698175906
transform 1 0 8400 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_142
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_157
timestamp 1698175906
transform 1 0 9464 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_159
timestamp 1698175906
transform 1 0 9576 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_261
timestamp 1698175906
transform 1 0 15288 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698175906
transform 1 0 16184 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 16296 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 2240 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 2464 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_111
timestamp 1698175906
transform 1 0 6888 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_129
timestamp 1698175906
transform 1 0 7896 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_137
timestamp 1698175906
transform 1 0 8344 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_141
timestamp 1698175906
transform 1 0 8568 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_143
timestamp 1698175906
transform 1 0 8680 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_159
timestamp 1698175906
transform 1 0 9576 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_161
timestamp 1698175906
transform 1 0 9688 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_177
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_210
timestamp 1698175906
transform 1 0 12432 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_218
timestamp 1698175906
transform 1 0 12880 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_220
timestamp 1698175906
transform 1 0 12992 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_229
timestamp 1698175906
transform 1 0 13496 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_104
timestamp 1698175906
transform 1 0 6496 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_120
timestamp 1698175906
transform 1 0 7392 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_128
timestamp 1698175906
transform 1 0 7840 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_130
timestamp 1698175906
transform 1 0 7952 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698175906
transform 1 0 8344 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 8456 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_146
timestamp 1698175906
transform 1 0 8848 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_148
timestamp 1698175906
transform 1 0 8960 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_182
timestamp 1698175906
transform 1 0 10864 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_203
timestamp 1698175906
transform 1 0 12040 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698175906
transform 1 0 12264 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698175906
transform 1 0 16128 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_115
timestamp 1698175906
transform 1 0 7112 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_119
timestamp 1698175906
transform 1 0 7336 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_129
timestamp 1698175906
transform 1 0 7896 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_145
timestamp 1698175906
transform 1 0 8792 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_147
timestamp 1698175906
transform 1 0 8904 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_167
timestamp 1698175906
transform 1 0 10024 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_209
timestamp 1698175906
transform 1 0 12376 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_213
timestamp 1698175906
transform 1 0 12600 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_236
timestamp 1698175906
transform 1 0 13888 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 14336 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_104
timestamp 1698175906
transform 1 0 6496 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_150
timestamp 1698175906
transform 1 0 9072 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_165
timestamp 1698175906
transform 1 0 9912 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_181
timestamp 1698175906
transform 1 0 10808 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_189
timestamp 1698175906
transform 1 0 11256 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_204
timestamp 1698175906
transform 1 0 12096 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698175906
transform 1 0 12320 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_241
timestamp 1698175906
transform 1 0 14168 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_273
timestamp 1698175906
transform 1 0 15960 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698175906
transform 1 0 16184 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 16296 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 2240 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 2464 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_123
timestamp 1698175906
transform 1 0 7560 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_131
timestamp 1698175906
transform 1 0 8008 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_161
timestamp 1698175906
transform 1 0 9688 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_167
timestamp 1698175906
transform 1 0 10024 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_177
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_181
timestamp 1698175906
transform 1 0 10808 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_240
timestamp 1698175906
transform 1 0 14112 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 14336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 18648 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698175906
transform 1 0 8288 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_150
timestamp 1698175906
transform 1 0 9072 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_185
timestamp 1698175906
transform 1 0 11032 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_193
timestamp 1698175906
transform 1 0 11480 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_197
timestamp 1698175906
transform 1 0 11704 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_204
timestamp 1698175906
transform 1 0 12096 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698175906
transform 1 0 12320 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_212
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_220
timestamp 1698175906
transform 1 0 12992 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_222
timestamp 1698175906
transform 1 0 13104 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_228
timestamp 1698175906
transform 1 0 13440 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_260
timestamp 1698175906
transform 1 0 15232 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 16128 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698175906
transform 1 0 10248 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_191
timestamp 1698175906
transform 1 0 11368 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_223
timestamp 1698175906
transform 1 0 13160 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_239
timestamp 1698175906
transform 1 0 14056 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698175906
transform 1 0 14280 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_174
timestamp 1698175906
transform 1 0 10416 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_183
timestamp 1698175906
transform 1 0 10920 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_199
timestamp 1698175906
transform 1 0 11816 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698175906
transform 1 0 12264 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 12376 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_6
timestamp 1698175906
transform 1 0 1008 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_22
timestamp 1698175906
transform 1 0 1904 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_30
timestamp 1698175906
transform 1 0 2352 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_174
timestamp 1698175906
transform 1 0 10416 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_178
timestamp 1698175906
transform 1 0 10640 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_180
timestamp 1698175906
transform 1 0 10752 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 14000 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 15792 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 16240 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita46_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19992 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita46_26
timestamp 1698175906
transform -1 0 1008 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 8456 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform -1 0 2240 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform -1 0 2240 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform -1 0 2240 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 10808 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 18760 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 18760 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform -1 0 2240 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 18760 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 18760 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 2240 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 18760 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 10640 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform -1 0 2240 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 18760 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13104 400 13160 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 8400 0 8456 400 0 FreeSans 224 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 0 10752 400 10808 0 FreeSans 224 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 0 10416 400 10472 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 0 11088 400 11144 0 FreeSans 224 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 20600 2352 21000 2408 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 11424 20600 11480 21000 0 FreeSans 224 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 0 18144 400 18200 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 10752 20600 10808 21000 0 FreeSans 224 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 20600 10416 21000 10472 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 20600 10080 21000 10136 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 0 8400 400 8456 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 0 8736 400 8792 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 20600 9744 21000 9800 0 FreeSans 224 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 0 12432 400 12488 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 20600 12432 21000 12488 0 FreeSans 224 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 20600 10752 21000 10808 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 9744 400 9800 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 12096 20600 12152 21000 0 FreeSans 224 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 20600 9072 21000 9128 0 FreeSans 224 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 20600 9408 21000 9464 0 FreeSans 224 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 11116 9100 11116 9100 0 _000_
rlabel metal2 11452 12572 11452 12572 0 _001_
rlabel metal2 12852 12152 12852 12152 0 _002_
rlabel metal2 10192 8708 10192 8708 0 _003_
rlabel metal2 8596 8204 8596 8204 0 _004_
rlabel metal3 9100 12460 9100 12460 0 _005_
rlabel metal2 9884 11368 9884 11368 0 _006_
rlabel metal2 6692 9268 6692 9268 0 _007_
rlabel metal3 13188 12012 13188 12012 0 _008_
rlabel metal2 7756 12152 7756 12152 0 _009_
rlabel metal3 12964 9940 12964 9940 0 _010_
rlabel metal2 13468 10864 13468 10864 0 _011_
rlabel metal2 9772 12908 9772 12908 0 _012_
rlabel metal2 13104 8484 13104 8484 0 _013_
rlabel metal2 12740 9016 12740 9016 0 _014_
rlabel metal2 11284 10780 11284 10780 0 _015_
rlabel metal2 6748 8596 6748 8596 0 _016_
rlabel metal2 7252 8008 7252 8008 0 _017_
rlabel metal3 6440 10052 6440 10052 0 _018_
rlabel metal2 7028 11032 7028 11032 0 _019_
rlabel metal2 11564 10976 11564 10976 0 _020_
rlabel metal3 8428 9492 8428 9492 0 _021_
rlabel metal2 8316 8400 8316 8400 0 _022_
rlabel metal2 7196 9016 7196 9016 0 _023_
rlabel metal3 7840 8372 7840 8372 0 _024_
rlabel metal2 6860 10108 6860 10108 0 _025_
rlabel metal2 7812 11032 7812 11032 0 _026_
rlabel metal2 7364 11228 7364 11228 0 _027_
rlabel metal3 8932 9268 8932 9268 0 _028_
rlabel metal2 10108 9436 10108 9436 0 _029_
rlabel metal2 9856 9604 9856 9604 0 _030_
rlabel metal2 9996 10024 9996 10024 0 _031_
rlabel metal3 9492 9940 9492 9940 0 _032_
rlabel metal2 10892 10584 10892 10584 0 _033_
rlabel metal3 13020 9324 13020 9324 0 _034_
rlabel metal2 9268 10038 9268 10038 0 _035_
rlabel metal3 11228 9604 11228 9604 0 _036_
rlabel metal3 10192 12348 10192 12348 0 _037_
rlabel metal3 11816 9100 11816 9100 0 _038_
rlabel metal2 8960 11060 8960 11060 0 _039_
rlabel metal2 8820 10920 8820 10920 0 _040_
rlabel metal2 9884 11060 9884 11060 0 _041_
rlabel metal2 10276 11088 10276 11088 0 _042_
rlabel metal3 10584 11844 10584 11844 0 _043_
rlabel metal3 13580 11956 13580 11956 0 _044_
rlabel metal2 11732 12740 11732 12740 0 _045_
rlabel metal3 12292 9268 12292 9268 0 _046_
rlabel metal2 13160 11956 13160 11956 0 _047_
rlabel metal2 8708 9800 8708 9800 0 _048_
rlabel metal2 9128 7700 9128 7700 0 _049_
rlabel metal2 9100 12236 9100 12236 0 _050_
rlabel metal2 9464 11284 9464 11284 0 _051_
rlabel metal2 9828 12208 9828 12208 0 _052_
rlabel metal2 10164 11228 10164 11228 0 _053_
rlabel metal2 8232 10780 8232 10780 0 _054_
rlabel metal2 7644 11060 7644 11060 0 _055_
rlabel metal3 8764 10836 8764 10836 0 _056_
rlabel metal2 7364 9576 7364 9576 0 _057_
rlabel metal3 7112 9604 7112 9604 0 _058_
rlabel metal2 7868 10304 7868 10304 0 _059_
rlabel metal2 7756 9996 7756 9996 0 _060_
rlabel metal3 12992 11900 12992 11900 0 _061_
rlabel metal2 13580 12012 13580 12012 0 _062_
rlabel metal2 7868 12152 7868 12152 0 _063_
rlabel metal4 7532 11088 7532 11088 0 _064_
rlabel metal2 12628 10976 12628 10976 0 _065_
rlabel metal2 13804 9800 13804 9800 0 _066_
rlabel metal2 12852 10164 12852 10164 0 _067_
rlabel metal2 13524 10514 13524 10514 0 _068_
rlabel metal2 10136 13804 10136 13804 0 _069_
rlabel metal3 13636 9212 13636 9212 0 _070_
rlabel metal2 13524 9184 13524 9184 0 _071_
rlabel metal2 8764 12180 8764 12180 0 clk
rlabel metal2 11676 10556 11676 10556 0 clknet_0_clk
rlabel metal2 7980 10612 7980 10612 0 clknet_1_0__leaf_clk
rlabel metal2 10724 8736 10724 8736 0 clknet_1_1__leaf_clk
rlabel metal2 9828 8008 9828 8008 0 dut46.count\[0\]
rlabel metal2 9660 8400 9660 8400 0 dut46.count\[1\]
rlabel metal2 9492 12068 9492 12068 0 dut46.count\[2\]
rlabel metal2 10332 9912 10332 9912 0 dut46.count\[3\]
rlabel metal2 18788 11396 18788 11396 0 net1
rlabel metal2 14812 10388 14812 10388 0 net10
rlabel metal3 4760 8428 4760 8428 0 net11
rlabel metal2 5684 8596 5684 8596 0 net12
rlabel metal2 15092 9940 15092 9940 0 net13
rlabel metal2 13636 9072 13636 9072 0 net14
rlabel metal3 15960 11592 15960 11592 0 net15
rlabel metal3 7966 12404 7966 12404 0 net16
rlabel metal2 14028 12768 14028 12768 0 net17
rlabel metal2 10752 13468 10752 13468 0 net18
rlabel metal2 15204 10808 15204 10808 0 net19
rlabel metal2 8540 2982 8540 2982 0 net2
rlabel metal2 5628 9576 5628 9576 0 net20
rlabel metal2 14084 12712 14084 12712 0 net21
rlabel metal2 12628 16030 12628 16030 0 net22
rlabel metal2 14084 8596 14084 8596 0 net23
rlabel metal2 18844 9072 18844 9072 0 net24
rlabel metal2 20132 2408 20132 2408 0 net25
rlabel metal3 623 18172 623 18172 0 net26
rlabel metal2 6748 10416 6748 10416 0 net3
rlabel metal2 5012 10416 5012 10416 0 net4
rlabel metal2 5964 10948 5964 10948 0 net5
rlabel metal3 11788 13468 11788 13468 0 net6
rlabel metal2 15092 10752 15092 10752 0 net7
rlabel metal3 10948 14028 10948 14028 0 net8
rlabel metal3 15358 10276 15358 10276 0 net9
rlabel metal2 20020 11900 20020 11900 0 segm[0]
rlabel metal2 8428 1043 8428 1043 0 segm[10]
rlabel metal3 679 10780 679 10780 0 segm[11]
rlabel metal3 679 10444 679 10444 0 segm[12]
rlabel metal3 679 11116 679 11116 0 segm[13]
rlabel metal2 11452 19873 11452 19873 0 segm[2]
rlabel metal2 20020 11172 20020 11172 0 segm[3]
rlabel metal2 10780 19677 10780 19677 0 segm[5]
rlabel metal3 20321 10444 20321 10444 0 segm[6]
rlabel metal3 20321 10108 20321 10108 0 segm[7]
rlabel metal3 679 8428 679 8428 0 segm[8]
rlabel metal3 679 8764 679 8764 0 segm[9]
rlabel metal2 20020 9744 20020 9744 0 sel[0]
rlabel metal2 19684 8624 19684 8624 0 sel[10]
rlabel metal3 20321 11452 20321 11452 0 sel[11]
rlabel metal3 679 12460 679 12460 0 sel[1]
rlabel metal2 20020 12628 20020 12628 0 sel[2]
rlabel metal2 11116 19873 11116 19873 0 sel[3]
rlabel metal2 20020 10752 20020 10752 0 sel[4]
rlabel metal3 679 9772 679 9772 0 sel[5]
rlabel metal2 19964 12936 19964 12936 0 sel[6]
rlabel metal2 12124 19677 12124 19677 0 sel[7]
rlabel metal2 19964 8988 19964 8988 0 sel[8]
rlabel metal2 20020 9296 20020 9296 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
