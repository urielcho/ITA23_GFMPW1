magic
tech gf180mcuD
magscale 1 10
timestamp 1699641132
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 22094 38274 22146 38286
rect 22094 38210 22146 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 14802 38110 14814 38162
rect 14866 38110 14878 38162
rect 18834 38110 18846 38162
rect 18898 38110 18910 38162
rect 16370 37998 16382 38050
rect 16434 37998 16446 38050
rect 18050 37998 18062 38050
rect 18114 37998 18126 38050
rect 21074 37998 21086 38050
rect 21138 37998 21150 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 18398 37490 18450 37502
rect 18398 37426 18450 37438
rect 21422 37490 21474 37502
rect 21422 37426 21474 37438
rect 26798 37490 26850 37502
rect 26798 37426 26850 37438
rect 17378 37214 17390 37266
rect 17442 37214 17454 37266
rect 20402 37214 20414 37266
rect 20466 37214 20478 37266
rect 25778 37214 25790 37266
rect 25842 37214 25854 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 16718 36706 16770 36718
rect 16718 36642 16770 36654
rect 15698 36430 15710 36482
rect 15762 36430 15774 36482
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 16146 28030 16158 28082
rect 16210 28030 16222 28082
rect 13234 27806 13246 27858
rect 13298 27806 13310 27858
rect 17714 27806 17726 27858
rect 17778 27806 17790 27858
rect 16830 27746 16882 27758
rect 21198 27746 21250 27758
rect 13906 27694 13918 27746
rect 13970 27694 13982 27746
rect 18498 27694 18510 27746
rect 18562 27694 18574 27746
rect 20626 27694 20638 27746
rect 20690 27694 20702 27746
rect 16830 27682 16882 27694
rect 21198 27682 21250 27694
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 20750 27186 20802 27198
rect 20290 27134 20302 27186
rect 20354 27134 20366 27186
rect 20750 27122 20802 27134
rect 22990 27074 23042 27086
rect 15474 27022 15486 27074
rect 15538 27022 15550 27074
rect 16594 27022 16606 27074
rect 16658 27022 16670 27074
rect 17378 27022 17390 27074
rect 17442 27022 17454 27074
rect 23314 27022 23326 27074
rect 23378 27022 23390 27074
rect 22990 27010 23042 27022
rect 14814 26962 14866 26974
rect 14814 26898 14866 26910
rect 14926 26962 14978 26974
rect 15698 26910 15710 26962
rect 15762 26910 15774 26962
rect 16370 26910 16382 26962
rect 16434 26910 16446 26962
rect 18162 26910 18174 26962
rect 18226 26910 18238 26962
rect 14926 26898 14978 26910
rect 15150 26850 15202 26862
rect 15150 26786 15202 26798
rect 23102 26850 23154 26862
rect 23102 26786 23154 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 16382 26514 16434 26526
rect 16382 26450 16434 26462
rect 18958 26514 19010 26526
rect 18958 26450 19010 26462
rect 19854 26514 19906 26526
rect 19854 26450 19906 26462
rect 16046 26402 16098 26414
rect 16046 26338 16098 26350
rect 16158 26402 16210 26414
rect 16158 26338 16210 26350
rect 19742 26402 19794 26414
rect 19742 26338 19794 26350
rect 20414 26402 20466 26414
rect 20414 26338 20466 26350
rect 20974 26402 21026 26414
rect 20974 26338 21026 26350
rect 18846 26290 18898 26302
rect 18846 26226 18898 26238
rect 19070 26290 19122 26302
rect 19070 26226 19122 26238
rect 19518 26290 19570 26302
rect 19518 26226 19570 26238
rect 20078 26290 20130 26302
rect 20078 26226 20130 26238
rect 20302 26290 20354 26302
rect 20302 26226 20354 26238
rect 20862 26290 20914 26302
rect 21298 26238 21310 26290
rect 21362 26238 21374 26290
rect 37650 26238 37662 26290
rect 37714 26238 37726 26290
rect 20862 26226 20914 26238
rect 24670 26178 24722 26190
rect 22082 26126 22094 26178
rect 22146 26126 22158 26178
rect 24210 26126 24222 26178
rect 24274 26126 24286 26178
rect 24670 26114 24722 26126
rect 25790 26178 25842 26190
rect 25790 26114 25842 26126
rect 20414 26066 20466 26078
rect 20414 26002 20466 26014
rect 40014 26066 40066 26078
rect 40014 26002 40066 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 21870 25730 21922 25742
rect 21870 25666 21922 25678
rect 1934 25618 1986 25630
rect 22206 25618 22258 25630
rect 27582 25618 27634 25630
rect 18722 25566 18734 25618
rect 18786 25566 18798 25618
rect 25554 25566 25566 25618
rect 25618 25566 25630 25618
rect 26674 25566 26686 25618
rect 26738 25566 26750 25618
rect 1934 25554 1986 25566
rect 22206 25554 22258 25566
rect 27582 25554 27634 25566
rect 20078 25506 20130 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 15810 25454 15822 25506
rect 15874 25454 15886 25506
rect 20078 25442 20130 25454
rect 21758 25506 21810 25518
rect 21758 25442 21810 25454
rect 22094 25506 22146 25518
rect 22642 25454 22654 25506
rect 22706 25454 22718 25506
rect 22094 25442 22146 25454
rect 20190 25394 20242 25406
rect 16594 25342 16606 25394
rect 16658 25342 16670 25394
rect 20190 25330 20242 25342
rect 20414 25394 20466 25406
rect 20414 25330 20466 25342
rect 21422 25394 21474 25406
rect 21422 25330 21474 25342
rect 22318 25394 22370 25406
rect 26238 25394 26290 25406
rect 23426 25342 23438 25394
rect 23490 25342 23502 25394
rect 26338 25342 26350 25394
rect 26402 25342 26414 25394
rect 22318 25330 22370 25342
rect 26238 25330 26290 25342
rect 19182 25282 19234 25294
rect 19182 25218 19234 25230
rect 25902 25282 25954 25294
rect 25902 25218 25954 25230
rect 26126 25282 26178 25294
rect 26126 25218 26178 25230
rect 27470 25282 27522 25294
rect 27470 25218 27522 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 15038 24946 15090 24958
rect 15038 24882 15090 24894
rect 17614 24946 17666 24958
rect 17614 24882 17666 24894
rect 18510 24946 18562 24958
rect 18510 24882 18562 24894
rect 18622 24946 18674 24958
rect 18622 24882 18674 24894
rect 23438 24946 23490 24958
rect 23438 24882 23490 24894
rect 24558 24946 24610 24958
rect 24558 24882 24610 24894
rect 25342 24946 25394 24958
rect 25342 24882 25394 24894
rect 26450 24782 26462 24834
rect 26514 24782 26526 24834
rect 18846 24722 18898 24734
rect 22654 24722 22706 24734
rect 24446 24722 24498 24734
rect 14018 24670 14030 24722
rect 14082 24670 14094 24722
rect 19058 24670 19070 24722
rect 19122 24670 19134 24722
rect 22866 24670 22878 24722
rect 22930 24670 22942 24722
rect 23426 24670 23438 24722
rect 23490 24670 23502 24722
rect 25666 24670 25678 24722
rect 25730 24670 25742 24722
rect 18846 24658 18898 24670
rect 22654 24658 22706 24670
rect 24446 24658 24498 24670
rect 14590 24610 14642 24622
rect 11106 24558 11118 24610
rect 11170 24558 11182 24610
rect 13234 24558 13246 24610
rect 13298 24558 13310 24610
rect 14590 24546 14642 24558
rect 17726 24610 17778 24622
rect 17726 24546 17778 24558
rect 18734 24610 18786 24622
rect 28578 24558 28590 24610
rect 28642 24558 28654 24610
rect 18734 24546 18786 24558
rect 14478 24498 14530 24510
rect 24334 24498 24386 24510
rect 23202 24446 23214 24498
rect 23266 24446 23278 24498
rect 14478 24434 14530 24446
rect 24334 24434 24386 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 14478 24050 14530 24062
rect 14478 23986 14530 23998
rect 19630 24050 19682 24062
rect 23538 23998 23550 24050
rect 23602 23998 23614 24050
rect 19630 23986 19682 23998
rect 14254 23938 14306 23950
rect 14254 23874 14306 23886
rect 14366 23938 14418 23950
rect 14366 23874 14418 23886
rect 19406 23938 19458 23950
rect 19406 23874 19458 23886
rect 19742 23938 19794 23950
rect 19742 23874 19794 23886
rect 20078 23938 20130 23950
rect 22642 23886 22654 23938
rect 22706 23886 22718 23938
rect 20078 23874 20130 23886
rect 14590 23714 14642 23726
rect 14590 23650 14642 23662
rect 14702 23714 14754 23726
rect 19058 23662 19070 23714
rect 19122 23711 19134 23714
rect 19282 23711 19294 23714
rect 19122 23665 19294 23711
rect 19122 23662 19134 23665
rect 19282 23662 19294 23665
rect 19346 23662 19358 23714
rect 14702 23650 14754 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 19182 23378 19234 23390
rect 27134 23378 27186 23390
rect 17378 23326 17390 23378
rect 17442 23326 17454 23378
rect 19506 23326 19518 23378
rect 19570 23326 19582 23378
rect 21522 23326 21534 23378
rect 21586 23326 21598 23378
rect 19182 23314 19234 23326
rect 27134 23314 27186 23326
rect 20402 23214 20414 23266
rect 20466 23214 20478 23266
rect 14366 23154 14418 23166
rect 4274 23102 4286 23154
rect 4338 23102 4350 23154
rect 14018 23102 14030 23154
rect 14082 23102 14094 23154
rect 14366 23090 14418 23102
rect 14814 23154 14866 23166
rect 14814 23090 14866 23102
rect 14926 23154 14978 23166
rect 14926 23090 14978 23102
rect 15374 23154 15426 23166
rect 17602 23102 17614 23154
rect 17666 23102 17678 23154
rect 19730 23102 19742 23154
rect 19794 23102 19806 23154
rect 20626 23102 20638 23154
rect 20690 23102 20702 23154
rect 21746 23102 21758 23154
rect 21810 23102 21822 23154
rect 27458 23102 27470 23154
rect 27522 23102 27534 23154
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 15374 23090 15426 23102
rect 15150 23042 15202 23054
rect 11218 22990 11230 23042
rect 11282 22990 11294 23042
rect 13346 22990 13358 23042
rect 13410 22990 13422 23042
rect 15150 22978 15202 22990
rect 15262 23042 15314 23054
rect 15262 22978 15314 22990
rect 15822 23042 15874 23054
rect 15822 22978 15874 22990
rect 19070 23042 19122 23054
rect 19070 22978 19122 22990
rect 24446 23042 24498 23054
rect 28242 22990 28254 23042
rect 28306 22990 28318 23042
rect 30370 22990 30382 23042
rect 30434 22990 30446 23042
rect 24446 22978 24498 22990
rect 1934 22930 1986 22942
rect 1934 22866 1986 22878
rect 24558 22930 24610 22942
rect 24558 22866 24610 22878
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 13918 22594 13970 22606
rect 19854 22594 19906 22606
rect 14914 22542 14926 22594
rect 14978 22542 14990 22594
rect 13918 22530 13970 22542
rect 19854 22530 19906 22542
rect 28478 22594 28530 22606
rect 28478 22530 28530 22542
rect 1934 22482 1986 22494
rect 14478 22482 14530 22494
rect 9986 22430 9998 22482
rect 10050 22430 10062 22482
rect 12114 22430 12126 22482
rect 12178 22430 12190 22482
rect 1934 22418 1986 22430
rect 14478 22418 14530 22430
rect 20302 22482 20354 22494
rect 20302 22418 20354 22430
rect 21534 22482 21586 22494
rect 29262 22482 29314 22494
rect 22418 22430 22430 22482
rect 22482 22430 22494 22482
rect 24770 22430 24782 22482
rect 24834 22430 24846 22482
rect 26898 22430 26910 22482
rect 26962 22430 26974 22482
rect 21534 22418 21586 22430
rect 29262 22418 29314 22430
rect 40014 22482 40066 22494
rect 40014 22418 40066 22430
rect 14030 22370 14082 22382
rect 4274 22318 4286 22370
rect 4338 22318 4350 22370
rect 12898 22318 12910 22370
rect 12962 22318 12974 22370
rect 14030 22306 14082 22318
rect 14702 22370 14754 22382
rect 15710 22370 15762 22382
rect 15138 22318 15150 22370
rect 15202 22318 15214 22370
rect 15474 22318 15486 22370
rect 15538 22318 15550 22370
rect 14702 22306 14754 22318
rect 15710 22306 15762 22318
rect 15822 22370 15874 22382
rect 19406 22370 19458 22382
rect 16146 22318 16158 22370
rect 16210 22318 16222 22370
rect 16482 22318 16494 22370
rect 16546 22318 16558 22370
rect 15822 22306 15874 22318
rect 19406 22306 19458 22318
rect 19518 22370 19570 22382
rect 19518 22306 19570 22318
rect 19742 22370 19794 22382
rect 19742 22306 19794 22318
rect 20638 22370 20690 22382
rect 28030 22370 28082 22382
rect 21858 22318 21870 22370
rect 21922 22318 21934 22370
rect 22306 22318 22318 22370
rect 22370 22318 22382 22370
rect 23986 22318 23998 22370
rect 24050 22318 24062 22370
rect 27234 22318 27246 22370
rect 27298 22318 27310 22370
rect 27570 22318 27582 22370
rect 27634 22318 27646 22370
rect 20638 22306 20690 22318
rect 28030 22306 28082 22318
rect 28366 22370 28418 22382
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 28366 22306 28418 22318
rect 13918 22258 13970 22270
rect 13918 22194 13970 22206
rect 14366 22258 14418 22270
rect 20190 22258 20242 22270
rect 16706 22206 16718 22258
rect 16770 22206 16782 22258
rect 17378 22206 17390 22258
rect 17442 22206 17454 22258
rect 14366 22194 14418 22206
rect 20190 22194 20242 22206
rect 20526 22258 20578 22270
rect 20526 22194 20578 22206
rect 22990 22258 23042 22270
rect 22990 22194 23042 22206
rect 23214 22258 23266 22270
rect 23214 22194 23266 22206
rect 23550 22258 23602 22270
rect 23550 22194 23602 22206
rect 29150 22258 29202 22270
rect 29150 22194 29202 22206
rect 15934 22146 15986 22158
rect 23326 22146 23378 22158
rect 17490 22094 17502 22146
rect 17554 22094 17566 22146
rect 15934 22082 15986 22094
rect 23326 22082 23378 22094
rect 27806 22146 27858 22158
rect 27806 22082 27858 22094
rect 27918 22146 27970 22158
rect 27918 22082 27970 22094
rect 28478 22146 28530 22158
rect 28478 22082 28530 22094
rect 29374 22146 29426 22158
rect 29374 22082 29426 22094
rect 29598 22146 29650 22158
rect 29598 22082 29650 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 13134 21810 13186 21822
rect 13134 21746 13186 21758
rect 15710 21810 15762 21822
rect 15710 21746 15762 21758
rect 23774 21810 23826 21822
rect 23774 21746 23826 21758
rect 24334 21810 24386 21822
rect 24334 21746 24386 21758
rect 25230 21810 25282 21822
rect 25230 21746 25282 21758
rect 26238 21810 26290 21822
rect 26238 21746 26290 21758
rect 26798 21810 26850 21822
rect 26798 21746 26850 21758
rect 21534 21698 21586 21710
rect 14914 21646 14926 21698
rect 14978 21646 14990 21698
rect 21534 21634 21586 21646
rect 22766 21698 22818 21710
rect 22766 21634 22818 21646
rect 23662 21698 23714 21710
rect 23662 21634 23714 21646
rect 24110 21698 24162 21710
rect 26014 21698 26066 21710
rect 25554 21646 25566 21698
rect 25618 21646 25630 21698
rect 27906 21646 27918 21698
rect 27970 21646 27982 21698
rect 24110 21634 24162 21646
rect 26014 21634 26066 21646
rect 15262 21586 15314 21598
rect 4274 21534 4286 21586
rect 4338 21534 4350 21586
rect 15262 21522 15314 21534
rect 15822 21586 15874 21598
rect 18622 21586 18674 21598
rect 20078 21586 20130 21598
rect 18162 21534 18174 21586
rect 18226 21534 18238 21586
rect 19506 21534 19518 21586
rect 19570 21534 19582 21586
rect 15822 21522 15874 21534
rect 18622 21522 18674 21534
rect 20078 21522 20130 21534
rect 21310 21586 21362 21598
rect 21310 21522 21362 21534
rect 21646 21586 21698 21598
rect 23438 21586 23490 21598
rect 22978 21534 22990 21586
rect 23042 21534 23054 21586
rect 21646 21522 21698 21534
rect 23438 21522 23490 21534
rect 24334 21586 24386 21598
rect 24334 21522 24386 21534
rect 24670 21586 24722 21598
rect 24670 21522 24722 21534
rect 25902 21586 25954 21598
rect 27122 21534 27134 21586
rect 27186 21534 27198 21586
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 25902 21522 25954 21534
rect 23214 21474 23266 21486
rect 40014 21474 40066 21486
rect 19282 21422 19294 21474
rect 19346 21422 19358 21474
rect 20514 21422 20526 21474
rect 20578 21422 20590 21474
rect 30034 21422 30046 21474
rect 30098 21422 30110 21474
rect 23214 21410 23266 21422
rect 40014 21410 40066 21422
rect 1934 21362 1986 21374
rect 1934 21298 1986 21310
rect 15710 21362 15762 21374
rect 19058 21310 19070 21362
rect 19122 21310 19134 21362
rect 15710 21298 15762 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 17726 21026 17778 21038
rect 17726 20962 17778 20974
rect 19742 21026 19794 21038
rect 19742 20962 19794 20974
rect 18734 20914 18786 20926
rect 17154 20862 17166 20914
rect 17218 20862 17230 20914
rect 18734 20850 18786 20862
rect 19854 20914 19906 20926
rect 27134 20914 27186 20926
rect 23538 20862 23550 20914
rect 23602 20862 23614 20914
rect 19854 20850 19906 20862
rect 27134 20850 27186 20862
rect 15934 20802 15986 20814
rect 29486 20802 29538 20814
rect 16930 20750 16942 20802
rect 16994 20750 17006 20802
rect 17938 20750 17950 20802
rect 18002 20750 18014 20802
rect 19170 20750 19182 20802
rect 19234 20750 19246 20802
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 20626 20750 20638 20802
rect 20690 20750 20702 20802
rect 21298 20750 21310 20802
rect 21362 20750 21374 20802
rect 15934 20738 15986 20750
rect 29486 20738 29538 20750
rect 13470 20690 13522 20702
rect 13470 20626 13522 20638
rect 15598 20690 15650 20702
rect 15598 20626 15650 20638
rect 16158 20690 16210 20702
rect 29150 20690 29202 20702
rect 19394 20638 19406 20690
rect 19458 20638 19470 20690
rect 20402 20638 20414 20690
rect 20466 20638 20478 20690
rect 16158 20626 16210 20638
rect 29150 20626 29202 20638
rect 29262 20690 29314 20702
rect 29262 20626 29314 20638
rect 13582 20578 13634 20590
rect 13582 20514 13634 20526
rect 14142 20578 14194 20590
rect 14142 20514 14194 20526
rect 15710 20578 15762 20590
rect 15710 20514 15762 20526
rect 18622 20578 18674 20590
rect 18622 20514 18674 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 14466 20190 14478 20242
rect 14530 20190 14542 20242
rect 15810 20190 15822 20242
rect 15874 20190 15886 20242
rect 13246 20130 13298 20142
rect 12002 20078 12014 20130
rect 12066 20078 12078 20130
rect 13246 20066 13298 20078
rect 15038 20130 15090 20142
rect 16830 20130 16882 20142
rect 21086 20130 21138 20142
rect 16482 20078 16494 20130
rect 16546 20078 16558 20130
rect 20178 20078 20190 20130
rect 20242 20078 20254 20130
rect 15038 20066 15090 20078
rect 16830 20066 16882 20078
rect 21086 20066 21138 20078
rect 21422 20130 21474 20142
rect 21422 20066 21474 20078
rect 21534 20130 21586 20142
rect 21534 20066 21586 20078
rect 21870 20130 21922 20142
rect 23214 20130 23266 20142
rect 22194 20078 22206 20130
rect 22258 20078 22270 20130
rect 22866 20078 22878 20130
rect 22930 20078 22942 20130
rect 21870 20066 21922 20078
rect 23214 20066 23266 20078
rect 23438 20130 23490 20142
rect 23438 20066 23490 20078
rect 23998 20130 24050 20142
rect 23998 20066 24050 20078
rect 24110 20130 24162 20142
rect 24110 20066 24162 20078
rect 13582 20018 13634 20030
rect 12786 19966 12798 20018
rect 12850 19966 12862 20018
rect 13582 19954 13634 19966
rect 13806 20018 13858 20030
rect 13806 19954 13858 19966
rect 14030 20018 14082 20030
rect 14030 19954 14082 19966
rect 14478 20018 14530 20030
rect 14478 19954 14530 19966
rect 14590 20018 14642 20030
rect 14590 19954 14642 19966
rect 14814 20018 14866 20030
rect 14814 19954 14866 19966
rect 16158 20018 16210 20030
rect 19854 20018 19906 20030
rect 18162 19966 18174 20018
rect 18226 19966 18238 20018
rect 18610 19966 18622 20018
rect 18674 19966 18686 20018
rect 16158 19954 16210 19966
rect 19854 19954 19906 19966
rect 22542 20018 22594 20030
rect 22542 19954 22594 19966
rect 23774 20018 23826 20030
rect 23774 19954 23826 19966
rect 13358 19906 13410 19918
rect 9874 19854 9886 19906
rect 9938 19854 9950 19906
rect 13358 19842 13410 19854
rect 18734 19906 18786 19918
rect 23314 19854 23326 19906
rect 23378 19854 23390 19906
rect 18734 19842 18786 19854
rect 24110 19794 24162 19806
rect 24110 19730 24162 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 23214 19458 23266 19470
rect 23214 19394 23266 19406
rect 1934 19346 1986 19358
rect 40014 19346 40066 19358
rect 9986 19294 9998 19346
rect 10050 19294 10062 19346
rect 12114 19294 12126 19346
rect 12178 19294 12190 19346
rect 1934 19282 1986 19294
rect 40014 19282 40066 19294
rect 13582 19234 13634 19246
rect 4274 19182 4286 19234
rect 4338 19182 4350 19234
rect 12898 19182 12910 19234
rect 12962 19182 12974 19234
rect 13582 19170 13634 19182
rect 15822 19234 15874 19246
rect 22990 19234 23042 19246
rect 21522 19182 21534 19234
rect 21586 19182 21598 19234
rect 15822 19170 15874 19182
rect 22990 19170 23042 19182
rect 27918 19234 27970 19246
rect 27918 19170 27970 19182
rect 29150 19234 29202 19246
rect 37650 19182 37662 19234
rect 37714 19182 37726 19234
rect 29150 19170 29202 19182
rect 13806 19122 13858 19134
rect 13806 19058 13858 19070
rect 13918 19122 13970 19134
rect 29262 19122 29314 19134
rect 21298 19070 21310 19122
rect 21362 19070 21374 19122
rect 13918 19058 13970 19070
rect 29262 19058 29314 19070
rect 14366 19010 14418 19022
rect 14366 18946 14418 18958
rect 15486 19010 15538 19022
rect 15486 18946 15538 18958
rect 15710 19010 15762 19022
rect 15710 18946 15762 18958
rect 17054 19010 17106 19022
rect 27694 19010 27746 19022
rect 23538 18958 23550 19010
rect 23602 18958 23614 19010
rect 17054 18946 17106 18958
rect 27694 18946 27746 18958
rect 27806 19010 27858 19022
rect 27806 18946 27858 18958
rect 28142 19010 28194 19022
rect 28142 18946 28194 18958
rect 29486 19010 29538 19022
rect 29486 18946 29538 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 21646 18674 21698 18686
rect 21646 18610 21698 18622
rect 25678 18674 25730 18686
rect 25678 18610 25730 18622
rect 25902 18674 25954 18686
rect 25902 18610 25954 18622
rect 12898 18510 12910 18562
rect 12962 18510 12974 18562
rect 18274 18510 18286 18562
rect 18338 18510 18350 18562
rect 22530 18510 22542 18562
rect 22594 18510 22606 18562
rect 17950 18450 18002 18462
rect 4274 18398 4286 18450
rect 4338 18398 4350 18450
rect 13122 18398 13134 18450
rect 13186 18398 13198 18450
rect 13906 18398 13918 18450
rect 13970 18398 13982 18450
rect 17602 18398 17614 18450
rect 17666 18398 17678 18450
rect 17950 18386 18002 18398
rect 18622 18450 18674 18462
rect 18622 18386 18674 18398
rect 19070 18450 19122 18462
rect 20862 18450 20914 18462
rect 19506 18398 19518 18450
rect 19570 18398 19582 18450
rect 19070 18386 19122 18398
rect 20862 18386 20914 18398
rect 21086 18450 21138 18462
rect 21758 18450 21810 18462
rect 25454 18450 25506 18462
rect 21410 18398 21422 18450
rect 21474 18398 21486 18450
rect 22306 18398 22318 18450
rect 22370 18398 22382 18450
rect 27010 18398 27022 18450
rect 27074 18398 27086 18450
rect 37874 18398 37886 18450
rect 37938 18398 37950 18450
rect 21086 18386 21138 18398
rect 21758 18386 21810 18398
rect 25454 18386 25506 18398
rect 19966 18338 20018 18350
rect 14690 18286 14702 18338
rect 14754 18286 14766 18338
rect 16818 18286 16830 18338
rect 16882 18286 16894 18338
rect 17714 18286 17726 18338
rect 17778 18286 17790 18338
rect 19966 18274 20018 18286
rect 20638 18338 20690 18350
rect 20638 18274 20690 18286
rect 25790 18338 25842 18350
rect 25790 18274 25842 18286
rect 26686 18338 26738 18350
rect 27794 18286 27806 18338
rect 27858 18286 27870 18338
rect 29922 18286 29934 18338
rect 29986 18286 29998 18338
rect 26686 18274 26738 18286
rect 1934 18226 1986 18238
rect 25230 18226 25282 18238
rect 20290 18174 20302 18226
rect 20354 18174 20366 18226
rect 1934 18162 1986 18174
rect 25230 18162 25282 18174
rect 40014 18226 40066 18238
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 15150 17890 15202 17902
rect 15150 17826 15202 17838
rect 15486 17890 15538 17902
rect 15486 17826 15538 17838
rect 19630 17890 19682 17902
rect 19630 17826 19682 17838
rect 18510 17778 18562 17790
rect 27470 17778 27522 17790
rect 19842 17726 19854 17778
rect 19906 17726 19918 17778
rect 18510 17714 18562 17726
rect 27470 17714 27522 17726
rect 40014 17778 40066 17790
rect 40014 17714 40066 17726
rect 17502 17666 17554 17678
rect 27358 17666 27410 17678
rect 20514 17614 20526 17666
rect 20578 17614 20590 17666
rect 22642 17614 22654 17666
rect 22706 17614 22718 17666
rect 17502 17602 17554 17614
rect 27358 17602 27410 17614
rect 28030 17666 28082 17678
rect 28030 17602 28082 17614
rect 29150 17666 29202 17678
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 29150 17602 29202 17614
rect 18622 17554 18674 17566
rect 29262 17554 29314 17566
rect 19282 17502 19294 17554
rect 19346 17502 19358 17554
rect 26338 17502 26350 17554
rect 26402 17502 26414 17554
rect 18622 17490 18674 17502
rect 29262 17490 29314 17502
rect 15262 17442 15314 17454
rect 17838 17442 17890 17454
rect 18958 17442 19010 17454
rect 17154 17390 17166 17442
rect 17218 17390 17230 17442
rect 18162 17390 18174 17442
rect 18226 17390 18238 17442
rect 15262 17378 15314 17390
rect 17838 17378 17890 17390
rect 18958 17378 19010 17390
rect 19854 17442 19906 17454
rect 27582 17442 27634 17454
rect 20290 17390 20302 17442
rect 20354 17390 20366 17442
rect 19854 17378 19906 17390
rect 27582 17378 27634 17390
rect 29486 17442 29538 17454
rect 29486 17378 29538 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 19070 17106 19122 17118
rect 19070 17042 19122 17054
rect 19518 17106 19570 17118
rect 19518 17042 19570 17054
rect 23214 17106 23266 17118
rect 23214 17042 23266 17054
rect 14926 16994 14978 17006
rect 14926 16930 14978 16942
rect 16606 16994 16658 17006
rect 23102 16994 23154 17006
rect 20402 16942 20414 16994
rect 20466 16942 20478 16994
rect 21634 16942 21646 16994
rect 21698 16942 21710 16994
rect 16606 16930 16658 16942
rect 23102 16930 23154 16942
rect 23438 16994 23490 17006
rect 28018 16942 28030 16994
rect 28082 16942 28094 16994
rect 23438 16930 23490 16942
rect 15262 16882 15314 16894
rect 15262 16818 15314 16830
rect 15486 16882 15538 16894
rect 15486 16818 15538 16830
rect 19182 16882 19234 16894
rect 19182 16818 19234 16830
rect 20078 16882 20130 16894
rect 23550 16882 23602 16894
rect 20626 16830 20638 16882
rect 20690 16830 20702 16882
rect 21410 16830 21422 16882
rect 21474 16830 21486 16882
rect 27234 16830 27246 16882
rect 27298 16830 27310 16882
rect 20078 16818 20130 16830
rect 23550 16818 23602 16830
rect 15038 16770 15090 16782
rect 15038 16706 15090 16718
rect 16494 16770 16546 16782
rect 16494 16706 16546 16718
rect 26910 16770 26962 16782
rect 30146 16718 30158 16770
rect 30210 16718 30222 16770
rect 26910 16706 26962 16718
rect 16382 16658 16434 16670
rect 16382 16594 16434 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 16830 16210 16882 16222
rect 14242 16158 14254 16210
rect 14306 16158 14318 16210
rect 16370 16158 16382 16210
rect 16434 16158 16446 16210
rect 23986 16158 23998 16210
rect 24050 16158 24062 16210
rect 26114 16158 26126 16210
rect 26178 16158 26190 16210
rect 16830 16146 16882 16158
rect 19966 16098 20018 16110
rect 23214 16098 23266 16110
rect 27358 16098 27410 16110
rect 13570 16046 13582 16098
rect 13634 16046 13646 16098
rect 20514 16046 20526 16098
rect 20578 16046 20590 16098
rect 26898 16046 26910 16098
rect 26962 16046 26974 16098
rect 19966 16034 20018 16046
rect 23214 16034 23266 16046
rect 27358 16034 27410 16046
rect 22878 15986 22930 15998
rect 22878 15922 22930 15934
rect 23438 15986 23490 15998
rect 23438 15922 23490 15934
rect 20078 15874 20130 15886
rect 20078 15810 20130 15822
rect 20190 15874 20242 15886
rect 20190 15810 20242 15822
rect 22990 15874 23042 15886
rect 22990 15810 23042 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 22878 15538 22930 15550
rect 22878 15474 22930 15486
rect 23662 15426 23714 15438
rect 17378 15374 17390 15426
rect 17442 15374 17454 15426
rect 23426 15374 23438 15426
rect 23490 15374 23502 15426
rect 23662 15362 23714 15374
rect 23998 15426 24050 15438
rect 23998 15362 24050 15374
rect 16482 15262 16494 15314
rect 16546 15262 16558 15314
rect 17602 15262 17614 15314
rect 17666 15262 17678 15314
rect 23090 15262 23102 15314
rect 23154 15262 23166 15314
rect 24322 15262 24334 15314
rect 24386 15262 24398 15314
rect 23214 15202 23266 15214
rect 23214 15138 23266 15150
rect 24110 15202 24162 15214
rect 24110 15138 24162 15150
rect 16494 15090 16546 15102
rect 16494 15026 16546 15038
rect 16830 15090 16882 15102
rect 16830 15026 16882 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 15598 14754 15650 14766
rect 15598 14690 15650 14702
rect 15822 14754 15874 14766
rect 15822 14690 15874 14702
rect 17826 14590 17838 14642
rect 17890 14590 17902 14642
rect 19954 14590 19966 14642
rect 20018 14590 20030 14642
rect 22866 14590 22878 14642
rect 22930 14590 22942 14642
rect 24994 14590 25006 14642
rect 25058 14590 25070 14642
rect 22318 14530 22370 14542
rect 16034 14478 16046 14530
rect 16098 14478 16110 14530
rect 20738 14478 20750 14530
rect 20802 14478 20814 14530
rect 22318 14466 22370 14478
rect 22654 14530 22706 14542
rect 26238 14530 26290 14542
rect 25666 14478 25678 14530
rect 25730 14478 25742 14530
rect 22654 14466 22706 14478
rect 26238 14466 26290 14478
rect 15486 14418 15538 14430
rect 15486 14354 15538 14366
rect 16942 14418 16994 14430
rect 16942 14354 16994 14366
rect 17166 14418 17218 14430
rect 17166 14354 17218 14366
rect 17054 14306 17106 14318
rect 17054 14242 17106 14254
rect 21422 14306 21474 14318
rect 21422 14242 21474 14254
rect 22430 14306 22482 14318
rect 22430 14242 22482 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 18286 13970 18338 13982
rect 18286 13906 18338 13918
rect 18398 13970 18450 13982
rect 18398 13906 18450 13918
rect 14690 13806 14702 13858
rect 14754 13806 14766 13858
rect 22530 13806 22542 13858
rect 22594 13806 22606 13858
rect 18510 13746 18562 13758
rect 14018 13694 14030 13746
rect 14082 13694 14094 13746
rect 18834 13694 18846 13746
rect 18898 13694 18910 13746
rect 21746 13694 21758 13746
rect 21810 13694 21822 13746
rect 18510 13682 18562 13694
rect 17502 13634 17554 13646
rect 25342 13634 25394 13646
rect 16818 13582 16830 13634
rect 16882 13582 16894 13634
rect 24658 13582 24670 13634
rect 24722 13582 24734 13634
rect 17502 13570 17554 13582
rect 25342 13570 25394 13582
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 19294 13074 19346 13086
rect 25006 13074 25058 13086
rect 16594 13022 16606 13074
rect 16658 13022 16670 13074
rect 18722 13022 18734 13074
rect 18786 13022 18798 13074
rect 24434 13022 24446 13074
rect 24498 13022 24510 13074
rect 19294 13010 19346 13022
rect 25006 13010 25058 13022
rect 15922 12910 15934 12962
rect 15986 12910 15998 12962
rect 21522 12910 21534 12962
rect 21586 12910 21598 12962
rect 22306 12798 22318 12850
rect 22370 12798 22382 12850
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 19058 4286 19070 4338
rect 19122 4286 19134 4338
rect 25554 4286 25566 4338
rect 25618 4286 25630 4338
rect 20078 4114 20130 4126
rect 20078 4050 20130 4062
rect 26238 4114 26290 4126
rect 26238 4050 26290 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 17042 3502 17054 3554
rect 17106 3502 17118 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 18062 3330 18114 3342
rect 18062 3266 18114 3278
rect 35982 3330 36034 3342
rect 35982 3266 36034 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 22094 38222 22146 38274
rect 25566 38222 25618 38274
rect 14814 38110 14866 38162
rect 18846 38110 18898 38162
rect 16382 37998 16434 38050
rect 18062 37998 18114 38050
rect 21086 37998 21138 38050
rect 24558 37998 24610 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 18398 37438 18450 37490
rect 21422 37438 21474 37490
rect 26798 37438 26850 37490
rect 17390 37214 17442 37266
rect 20414 37214 20466 37266
rect 25790 37214 25842 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 16718 36654 16770 36706
rect 15710 36430 15762 36482
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 16158 28030 16210 28082
rect 13246 27806 13298 27858
rect 17726 27806 17778 27858
rect 13918 27694 13970 27746
rect 16830 27694 16882 27746
rect 18510 27694 18562 27746
rect 20638 27694 20690 27746
rect 21198 27694 21250 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 20302 27134 20354 27186
rect 20750 27134 20802 27186
rect 15486 27022 15538 27074
rect 16606 27022 16658 27074
rect 17390 27022 17442 27074
rect 22990 27022 23042 27074
rect 23326 27022 23378 27074
rect 14814 26910 14866 26962
rect 14926 26910 14978 26962
rect 15710 26910 15762 26962
rect 16382 26910 16434 26962
rect 18174 26910 18226 26962
rect 15150 26798 15202 26850
rect 23102 26798 23154 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 16382 26462 16434 26514
rect 18958 26462 19010 26514
rect 19854 26462 19906 26514
rect 16046 26350 16098 26402
rect 16158 26350 16210 26402
rect 19742 26350 19794 26402
rect 20414 26350 20466 26402
rect 20974 26350 21026 26402
rect 18846 26238 18898 26290
rect 19070 26238 19122 26290
rect 19518 26238 19570 26290
rect 20078 26238 20130 26290
rect 20302 26238 20354 26290
rect 20862 26238 20914 26290
rect 21310 26238 21362 26290
rect 37662 26238 37714 26290
rect 22094 26126 22146 26178
rect 24222 26126 24274 26178
rect 24670 26126 24722 26178
rect 25790 26126 25842 26178
rect 20414 26014 20466 26066
rect 40014 26014 40066 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 21870 25678 21922 25730
rect 1934 25566 1986 25618
rect 18734 25566 18786 25618
rect 22206 25566 22258 25618
rect 25566 25566 25618 25618
rect 26686 25566 26738 25618
rect 27582 25566 27634 25618
rect 4286 25454 4338 25506
rect 15822 25454 15874 25506
rect 20078 25454 20130 25506
rect 21758 25454 21810 25506
rect 22094 25454 22146 25506
rect 22654 25454 22706 25506
rect 16606 25342 16658 25394
rect 20190 25342 20242 25394
rect 20414 25342 20466 25394
rect 21422 25342 21474 25394
rect 22318 25342 22370 25394
rect 23438 25342 23490 25394
rect 26238 25342 26290 25394
rect 26350 25342 26402 25394
rect 19182 25230 19234 25282
rect 25902 25230 25954 25282
rect 26126 25230 26178 25282
rect 27470 25230 27522 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 15038 24894 15090 24946
rect 17614 24894 17666 24946
rect 18510 24894 18562 24946
rect 18622 24894 18674 24946
rect 23438 24894 23490 24946
rect 24558 24894 24610 24946
rect 25342 24894 25394 24946
rect 26462 24782 26514 24834
rect 14030 24670 14082 24722
rect 18846 24670 18898 24722
rect 19070 24670 19122 24722
rect 22654 24670 22706 24722
rect 22878 24670 22930 24722
rect 23438 24670 23490 24722
rect 24446 24670 24498 24722
rect 25678 24670 25730 24722
rect 11118 24558 11170 24610
rect 13246 24558 13298 24610
rect 14590 24558 14642 24610
rect 17726 24558 17778 24610
rect 18734 24558 18786 24610
rect 28590 24558 28642 24610
rect 14478 24446 14530 24498
rect 23214 24446 23266 24498
rect 24334 24446 24386 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 14478 23998 14530 24050
rect 19630 23998 19682 24050
rect 23550 23998 23602 24050
rect 14254 23886 14306 23938
rect 14366 23886 14418 23938
rect 19406 23886 19458 23938
rect 19742 23886 19794 23938
rect 20078 23886 20130 23938
rect 22654 23886 22706 23938
rect 14590 23662 14642 23714
rect 14702 23662 14754 23714
rect 19070 23662 19122 23714
rect 19294 23662 19346 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 17390 23326 17442 23378
rect 19182 23326 19234 23378
rect 19518 23326 19570 23378
rect 21534 23326 21586 23378
rect 27134 23326 27186 23378
rect 20414 23214 20466 23266
rect 4286 23102 4338 23154
rect 14030 23102 14082 23154
rect 14366 23102 14418 23154
rect 14814 23102 14866 23154
rect 14926 23102 14978 23154
rect 15374 23102 15426 23154
rect 17614 23102 17666 23154
rect 19742 23102 19794 23154
rect 20638 23102 20690 23154
rect 21758 23102 21810 23154
rect 27470 23102 27522 23154
rect 37662 23102 37714 23154
rect 11230 22990 11282 23042
rect 13358 22990 13410 23042
rect 15150 22990 15202 23042
rect 15262 22990 15314 23042
rect 15822 22990 15874 23042
rect 19070 22990 19122 23042
rect 24446 22990 24498 23042
rect 28254 22990 28306 23042
rect 30382 22990 30434 23042
rect 1934 22878 1986 22930
rect 24558 22878 24610 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 13918 22542 13970 22594
rect 14926 22542 14978 22594
rect 19854 22542 19906 22594
rect 28478 22542 28530 22594
rect 1934 22430 1986 22482
rect 9998 22430 10050 22482
rect 12126 22430 12178 22482
rect 14478 22430 14530 22482
rect 20302 22430 20354 22482
rect 21534 22430 21586 22482
rect 22430 22430 22482 22482
rect 24782 22430 24834 22482
rect 26910 22430 26962 22482
rect 29262 22430 29314 22482
rect 40014 22430 40066 22482
rect 4286 22318 4338 22370
rect 12910 22318 12962 22370
rect 14030 22318 14082 22370
rect 14702 22318 14754 22370
rect 15150 22318 15202 22370
rect 15486 22318 15538 22370
rect 15710 22318 15762 22370
rect 15822 22318 15874 22370
rect 16158 22318 16210 22370
rect 16494 22318 16546 22370
rect 19406 22318 19458 22370
rect 19518 22318 19570 22370
rect 19742 22318 19794 22370
rect 20638 22318 20690 22370
rect 21870 22318 21922 22370
rect 22318 22318 22370 22370
rect 23998 22318 24050 22370
rect 27246 22318 27298 22370
rect 27582 22318 27634 22370
rect 28030 22318 28082 22370
rect 28366 22318 28418 22370
rect 37662 22318 37714 22370
rect 13918 22206 13970 22258
rect 14366 22206 14418 22258
rect 16718 22206 16770 22258
rect 17390 22206 17442 22258
rect 20190 22206 20242 22258
rect 20526 22206 20578 22258
rect 22990 22206 23042 22258
rect 23214 22206 23266 22258
rect 23550 22206 23602 22258
rect 29150 22206 29202 22258
rect 15934 22094 15986 22146
rect 17502 22094 17554 22146
rect 23326 22094 23378 22146
rect 27806 22094 27858 22146
rect 27918 22094 27970 22146
rect 28478 22094 28530 22146
rect 29374 22094 29426 22146
rect 29598 22094 29650 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 13134 21758 13186 21810
rect 15710 21758 15762 21810
rect 23774 21758 23826 21810
rect 24334 21758 24386 21810
rect 25230 21758 25282 21810
rect 26238 21758 26290 21810
rect 26798 21758 26850 21810
rect 14926 21646 14978 21698
rect 21534 21646 21586 21698
rect 22766 21646 22818 21698
rect 23662 21646 23714 21698
rect 24110 21646 24162 21698
rect 25566 21646 25618 21698
rect 26014 21646 26066 21698
rect 27918 21646 27970 21698
rect 4286 21534 4338 21586
rect 15262 21534 15314 21586
rect 15822 21534 15874 21586
rect 18174 21534 18226 21586
rect 18622 21534 18674 21586
rect 19518 21534 19570 21586
rect 20078 21534 20130 21586
rect 21310 21534 21362 21586
rect 21646 21534 21698 21586
rect 22990 21534 23042 21586
rect 23438 21534 23490 21586
rect 24334 21534 24386 21586
rect 24670 21534 24722 21586
rect 25902 21534 25954 21586
rect 27134 21534 27186 21586
rect 37662 21534 37714 21586
rect 19294 21422 19346 21474
rect 20526 21422 20578 21474
rect 23214 21422 23266 21474
rect 30046 21422 30098 21474
rect 40014 21422 40066 21474
rect 1934 21310 1986 21362
rect 15710 21310 15762 21362
rect 19070 21310 19122 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 17726 20974 17778 21026
rect 19742 20974 19794 21026
rect 17166 20862 17218 20914
rect 18734 20862 18786 20914
rect 19854 20862 19906 20914
rect 23550 20862 23602 20914
rect 27134 20862 27186 20914
rect 15934 20750 15986 20802
rect 16942 20750 16994 20802
rect 17950 20750 18002 20802
rect 19182 20750 19234 20802
rect 20078 20750 20130 20802
rect 20638 20750 20690 20802
rect 21310 20750 21362 20802
rect 29486 20750 29538 20802
rect 13470 20638 13522 20690
rect 15598 20638 15650 20690
rect 16158 20638 16210 20690
rect 19406 20638 19458 20690
rect 20414 20638 20466 20690
rect 29150 20638 29202 20690
rect 29262 20638 29314 20690
rect 13582 20526 13634 20578
rect 14142 20526 14194 20578
rect 15710 20526 15762 20578
rect 18622 20526 18674 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 14478 20190 14530 20242
rect 15822 20190 15874 20242
rect 12014 20078 12066 20130
rect 13246 20078 13298 20130
rect 15038 20078 15090 20130
rect 16494 20078 16546 20130
rect 16830 20078 16882 20130
rect 20190 20078 20242 20130
rect 21086 20078 21138 20130
rect 21422 20078 21474 20130
rect 21534 20078 21586 20130
rect 21870 20078 21922 20130
rect 22206 20078 22258 20130
rect 22878 20078 22930 20130
rect 23214 20078 23266 20130
rect 23438 20078 23490 20130
rect 23998 20078 24050 20130
rect 24110 20078 24162 20130
rect 12798 19966 12850 20018
rect 13582 19966 13634 20018
rect 13806 19966 13858 20018
rect 14030 19966 14082 20018
rect 14478 19966 14530 20018
rect 14590 19966 14642 20018
rect 14814 19966 14866 20018
rect 16158 19966 16210 20018
rect 18174 19966 18226 20018
rect 18622 19966 18674 20018
rect 19854 19966 19906 20018
rect 22542 19966 22594 20018
rect 23774 19966 23826 20018
rect 9886 19854 9938 19906
rect 13358 19854 13410 19906
rect 18734 19854 18786 19906
rect 23326 19854 23378 19906
rect 24110 19742 24162 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 23214 19406 23266 19458
rect 1934 19294 1986 19346
rect 9998 19294 10050 19346
rect 12126 19294 12178 19346
rect 40014 19294 40066 19346
rect 4286 19182 4338 19234
rect 12910 19182 12962 19234
rect 13582 19182 13634 19234
rect 15822 19182 15874 19234
rect 21534 19182 21586 19234
rect 22990 19182 23042 19234
rect 27918 19182 27970 19234
rect 29150 19182 29202 19234
rect 37662 19182 37714 19234
rect 13806 19070 13858 19122
rect 13918 19070 13970 19122
rect 21310 19070 21362 19122
rect 29262 19070 29314 19122
rect 14366 18958 14418 19010
rect 15486 18958 15538 19010
rect 15710 18958 15762 19010
rect 17054 18958 17106 19010
rect 23550 18958 23602 19010
rect 27694 18958 27746 19010
rect 27806 18958 27858 19010
rect 28142 18958 28194 19010
rect 29486 18958 29538 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 21646 18622 21698 18674
rect 25678 18622 25730 18674
rect 25902 18622 25954 18674
rect 12910 18510 12962 18562
rect 18286 18510 18338 18562
rect 22542 18510 22594 18562
rect 4286 18398 4338 18450
rect 13134 18398 13186 18450
rect 13918 18398 13970 18450
rect 17614 18398 17666 18450
rect 17950 18398 18002 18450
rect 18622 18398 18674 18450
rect 19070 18398 19122 18450
rect 19518 18398 19570 18450
rect 20862 18398 20914 18450
rect 21086 18398 21138 18450
rect 21422 18398 21474 18450
rect 21758 18398 21810 18450
rect 22318 18398 22370 18450
rect 25454 18398 25506 18450
rect 27022 18398 27074 18450
rect 37886 18398 37938 18450
rect 14702 18286 14754 18338
rect 16830 18286 16882 18338
rect 17726 18286 17778 18338
rect 19966 18286 20018 18338
rect 20638 18286 20690 18338
rect 25790 18286 25842 18338
rect 26686 18286 26738 18338
rect 27806 18286 27858 18338
rect 29934 18286 29986 18338
rect 1934 18174 1986 18226
rect 20302 18174 20354 18226
rect 25230 18174 25282 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 15150 17838 15202 17890
rect 15486 17838 15538 17890
rect 19630 17838 19682 17890
rect 18510 17726 18562 17778
rect 19854 17726 19906 17778
rect 27470 17726 27522 17778
rect 40014 17726 40066 17778
rect 17502 17614 17554 17666
rect 20526 17614 20578 17666
rect 22654 17614 22706 17666
rect 27358 17614 27410 17666
rect 28030 17614 28082 17666
rect 29150 17614 29202 17666
rect 37662 17614 37714 17666
rect 18622 17502 18674 17554
rect 19294 17502 19346 17554
rect 26350 17502 26402 17554
rect 29262 17502 29314 17554
rect 15262 17390 15314 17442
rect 17166 17390 17218 17442
rect 17838 17390 17890 17442
rect 18174 17390 18226 17442
rect 18958 17390 19010 17442
rect 19854 17390 19906 17442
rect 20302 17390 20354 17442
rect 27582 17390 27634 17442
rect 29486 17390 29538 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 19070 17054 19122 17106
rect 19518 17054 19570 17106
rect 23214 17054 23266 17106
rect 14926 16942 14978 16994
rect 16606 16942 16658 16994
rect 20414 16942 20466 16994
rect 21646 16942 21698 16994
rect 23102 16942 23154 16994
rect 23438 16942 23490 16994
rect 28030 16942 28082 16994
rect 15262 16830 15314 16882
rect 15486 16830 15538 16882
rect 19182 16830 19234 16882
rect 20078 16830 20130 16882
rect 20638 16830 20690 16882
rect 21422 16830 21474 16882
rect 23550 16830 23602 16882
rect 27246 16830 27298 16882
rect 15038 16718 15090 16770
rect 16494 16718 16546 16770
rect 26910 16718 26962 16770
rect 30158 16718 30210 16770
rect 16382 16606 16434 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 14254 16158 14306 16210
rect 16382 16158 16434 16210
rect 16830 16158 16882 16210
rect 23998 16158 24050 16210
rect 26126 16158 26178 16210
rect 13582 16046 13634 16098
rect 19966 16046 20018 16098
rect 20526 16046 20578 16098
rect 23214 16046 23266 16098
rect 26910 16046 26962 16098
rect 27358 16046 27410 16098
rect 22878 15934 22930 15986
rect 23438 15934 23490 15986
rect 20078 15822 20130 15874
rect 20190 15822 20242 15874
rect 22990 15822 23042 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 22878 15486 22930 15538
rect 17390 15374 17442 15426
rect 23438 15374 23490 15426
rect 23662 15374 23714 15426
rect 23998 15374 24050 15426
rect 16494 15262 16546 15314
rect 17614 15262 17666 15314
rect 23102 15262 23154 15314
rect 24334 15262 24386 15314
rect 23214 15150 23266 15202
rect 24110 15150 24162 15202
rect 16494 15038 16546 15090
rect 16830 15038 16882 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 15598 14702 15650 14754
rect 15822 14702 15874 14754
rect 17838 14590 17890 14642
rect 19966 14590 20018 14642
rect 22878 14590 22930 14642
rect 25006 14590 25058 14642
rect 16046 14478 16098 14530
rect 20750 14478 20802 14530
rect 22318 14478 22370 14530
rect 22654 14478 22706 14530
rect 25678 14478 25730 14530
rect 26238 14478 26290 14530
rect 15486 14366 15538 14418
rect 16942 14366 16994 14418
rect 17166 14366 17218 14418
rect 17054 14254 17106 14306
rect 21422 14254 21474 14306
rect 22430 14254 22482 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 18286 13918 18338 13970
rect 18398 13918 18450 13970
rect 14702 13806 14754 13858
rect 22542 13806 22594 13858
rect 14030 13694 14082 13746
rect 18510 13694 18562 13746
rect 18846 13694 18898 13746
rect 21758 13694 21810 13746
rect 16830 13582 16882 13634
rect 17502 13582 17554 13634
rect 24670 13582 24722 13634
rect 25342 13582 25394 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 16606 13022 16658 13074
rect 18734 13022 18786 13074
rect 19294 13022 19346 13074
rect 24446 13022 24498 13074
rect 25006 13022 25058 13074
rect 15934 12910 15986 12962
rect 21534 12910 21586 12962
rect 22318 12798 22370 12850
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 19070 4286 19122 4338
rect 25566 4286 25618 4338
rect 20078 4062 20130 4114
rect 26238 4062 26290 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 25566 3614 25618 3666
rect 17054 3502 17106 3554
rect 24558 3502 24610 3554
rect 18062 3278 18114 3330
rect 35982 3278 36034 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 14784 41200 14896 42000
rect 15456 41200 15568 42000
rect 16128 41200 16240 42000
rect 18816 41200 18928 42000
rect 20160 41200 20272 42000
rect 20832 41200 20944 42000
rect 24192 41200 24304 42000
rect 25536 41200 25648 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 14812 38162 14868 41200
rect 14812 38110 14814 38162
rect 14866 38110 14868 38162
rect 14812 38098 14868 38110
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 15484 36708 15540 41200
rect 16156 37492 16212 41200
rect 18844 38162 18900 41200
rect 18844 38110 18846 38162
rect 18898 38110 18900 38162
rect 18844 38098 18900 38110
rect 16156 37426 16212 37436
rect 16380 38050 16436 38062
rect 16380 37998 16382 38050
rect 16434 37998 16436 38050
rect 15484 36642 15540 36652
rect 15708 36482 15764 36494
rect 15708 36430 15710 36482
rect 15762 36430 15764 36482
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 13244 27858 13300 27870
rect 13244 27806 13246 27858
rect 13298 27806 13300 27858
rect 4172 27636 4228 27646
rect 1932 25618 1988 25630
rect 1932 25566 1934 25618
rect 1986 25566 1988 25618
rect 1932 24948 1988 25566
rect 1932 24882 1988 24892
rect 1932 22932 1988 22942
rect 1932 22838 1988 22876
rect 1932 22484 1988 22494
rect 1932 22390 1988 22428
rect 1932 21362 1988 21374
rect 1932 21310 1934 21362
rect 1986 21310 1988 21362
rect 1932 20916 1988 21310
rect 4172 21028 4228 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4284 25506 4340 25518
rect 4284 25454 4286 25506
rect 4338 25454 4340 25506
rect 4284 24612 4340 25454
rect 13244 25284 13300 27806
rect 13916 27746 13972 27758
rect 13916 27694 13918 27746
rect 13970 27694 13972 27746
rect 13916 26516 13972 27694
rect 14924 27076 14980 27086
rect 13916 26450 13972 26460
rect 14812 26962 14868 26974
rect 14812 26910 14814 26962
rect 14866 26910 14868 26962
rect 13244 25218 13300 25228
rect 14028 25284 14084 25294
rect 14028 24722 14084 25228
rect 14028 24670 14030 24722
rect 14082 24670 14084 24722
rect 4284 24546 4340 24556
rect 11116 24612 11172 24622
rect 11116 24518 11172 24556
rect 13244 24610 13300 24622
rect 13244 24558 13246 24610
rect 13298 24558 13300 24610
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 13244 24052 13300 24558
rect 13244 23986 13300 23996
rect 4284 23156 4340 23166
rect 4284 23062 4340 23100
rect 9996 23156 10052 23166
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 9996 22482 10052 23100
rect 14028 23154 14084 24670
rect 14588 24612 14644 24622
rect 14588 24518 14644 24556
rect 14476 24500 14532 24510
rect 14252 24498 14532 24500
rect 14252 24446 14478 24498
rect 14530 24446 14532 24498
rect 14252 24444 14532 24446
rect 14252 23938 14308 24444
rect 14476 24434 14532 24444
rect 14476 24052 14532 24062
rect 14476 23958 14532 23996
rect 14252 23886 14254 23938
rect 14306 23886 14308 23938
rect 14252 23874 14308 23886
rect 14364 23940 14420 23950
rect 14364 23846 14420 23884
rect 14812 23940 14868 26910
rect 14924 26962 14980 27020
rect 15484 27076 15540 27086
rect 15484 26982 15540 27020
rect 14924 26910 14926 26962
rect 14978 26910 14980 26962
rect 14924 26898 14980 26910
rect 15708 26962 15764 36430
rect 16156 28084 16212 28094
rect 16156 27990 16212 28028
rect 15708 26910 15710 26962
rect 15762 26910 15764 26962
rect 15708 26898 15764 26910
rect 16380 26962 16436 37998
rect 18060 38052 18116 38062
rect 18060 37958 18116 37996
rect 18732 38052 18788 38062
rect 18396 37492 18452 37502
rect 18396 37398 18452 37436
rect 17388 37266 17444 37278
rect 17388 37214 17390 37266
rect 17442 37214 17444 37266
rect 16716 36708 16772 36718
rect 16716 36614 16772 36652
rect 16604 28084 16660 28094
rect 16604 27076 16660 28028
rect 17388 28084 17444 37214
rect 17388 28018 17444 28028
rect 17724 27858 17780 27870
rect 17724 27806 17726 27858
rect 17778 27806 17780 27858
rect 16604 26982 16660 27020
rect 16828 27746 16884 27758
rect 16828 27694 16830 27746
rect 16882 27694 16884 27746
rect 16828 27076 16884 27694
rect 17388 27076 17444 27086
rect 17724 27076 17780 27806
rect 16828 27074 17780 27076
rect 16828 27022 17390 27074
rect 17442 27022 17780 27074
rect 16828 27020 17780 27022
rect 18508 27746 18564 27758
rect 18508 27694 18510 27746
rect 18562 27694 18564 27746
rect 16380 26910 16382 26962
rect 16434 26910 16436 26962
rect 16380 26898 16436 26910
rect 15148 26850 15204 26862
rect 15148 26798 15150 26850
rect 15202 26798 15204 26850
rect 15148 26404 15204 26798
rect 16380 26516 16436 26526
rect 16380 26422 16436 26460
rect 15148 26338 15204 26348
rect 16044 26404 16100 26414
rect 16044 26310 16100 26348
rect 16156 26402 16212 26414
rect 16156 26350 16158 26402
rect 16210 26350 16212 26402
rect 15820 25506 15876 25518
rect 15820 25454 15822 25506
rect 15874 25454 15876 25506
rect 15036 25284 15092 25294
rect 15036 24946 15092 25228
rect 15820 25284 15876 25454
rect 16156 25396 16212 26350
rect 16156 25330 16212 25340
rect 16604 25394 16660 25406
rect 16604 25342 16606 25394
rect 16658 25342 16660 25394
rect 15820 25218 15876 25228
rect 15036 24894 15038 24946
rect 15090 24894 15092 24946
rect 15036 24882 15092 24894
rect 16604 24948 16660 25342
rect 16828 25284 16884 27020
rect 17388 27010 17444 27020
rect 18172 26962 18228 26974
rect 18172 26910 18174 26962
rect 18226 26910 18228 26962
rect 18172 26516 18228 26910
rect 18172 26450 18228 26460
rect 18508 26180 18564 27694
rect 18508 26114 18564 26124
rect 18732 25618 18788 37996
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20188 37492 20244 41200
rect 20860 38276 20916 41200
rect 20860 38210 20916 38220
rect 22092 38276 22148 38286
rect 22092 38182 22148 38220
rect 24220 38276 24276 41200
rect 25564 38612 25620 41200
rect 25564 38546 25620 38556
rect 26796 38612 26852 38622
rect 24220 38210 24276 38220
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 20188 37426 20244 37436
rect 21084 38050 21140 38062
rect 21084 37998 21086 38050
rect 21138 37998 21140 38050
rect 20412 37266 20468 37278
rect 20412 37214 20414 37266
rect 20466 37214 20468 37266
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20412 31948 20468 37214
rect 21084 31948 21140 37998
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 21420 37492 21476 37502
rect 21420 37398 21476 37436
rect 20300 31892 20468 31948
rect 20636 31892 21140 31948
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20300 27188 20356 31892
rect 20636 27746 20692 31892
rect 21196 27748 21252 27758
rect 20636 27694 20638 27746
rect 20690 27694 20692 27746
rect 20300 27186 20580 27188
rect 20300 27134 20302 27186
rect 20354 27134 20580 27186
rect 20300 27132 20580 27134
rect 20300 27122 20356 27132
rect 20188 26740 20244 26750
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 18956 26516 19012 26526
rect 19852 26516 19908 26526
rect 20188 26516 20244 26684
rect 18956 26422 19012 26460
rect 19404 26460 19684 26516
rect 18732 25566 18734 25618
rect 18786 25566 18788 25618
rect 16828 25218 16884 25228
rect 17500 25396 17556 25406
rect 16604 24882 16660 24892
rect 14812 23874 14868 23884
rect 17388 24836 17444 24846
rect 17388 23940 17444 24780
rect 14588 23714 14644 23726
rect 14588 23662 14590 23714
rect 14642 23662 14644 23714
rect 14588 23380 14644 23662
rect 14700 23714 14756 23726
rect 14700 23662 14702 23714
rect 14754 23662 14756 23714
rect 14700 23604 14756 23662
rect 14700 23538 14756 23548
rect 16492 23492 16548 23502
rect 14588 23324 15092 23380
rect 14364 23156 14420 23166
rect 14028 23102 14030 23154
rect 14082 23102 14084 23154
rect 11228 23042 11284 23054
rect 11228 22990 11230 23042
rect 11282 22990 11284 23042
rect 11228 22708 11284 22990
rect 11228 22642 11284 22652
rect 12908 23044 12964 23054
rect 9996 22430 9998 22482
rect 10050 22430 10052 22482
rect 4284 22372 4340 22382
rect 4284 22278 4340 22316
rect 9996 22260 10052 22430
rect 12124 22596 12180 22606
rect 12124 22482 12180 22540
rect 12124 22430 12126 22482
rect 12178 22430 12180 22482
rect 12124 22418 12180 22430
rect 9996 22194 10052 22204
rect 12908 22370 12964 22988
rect 13356 23042 13412 23054
rect 13356 22990 13358 23042
rect 13410 22990 13412 23042
rect 13356 22484 13412 22990
rect 14028 23044 14084 23102
rect 14028 22978 14084 22988
rect 14140 23154 14420 23156
rect 14140 23102 14366 23154
rect 14418 23102 14420 23154
rect 14140 23100 14420 23102
rect 13916 22596 13972 22606
rect 14140 22596 14196 23100
rect 14364 23090 14420 23100
rect 14812 23154 14868 23166
rect 14812 23102 14814 23154
rect 14866 23102 14868 23154
rect 13916 22594 14196 22596
rect 13916 22542 13918 22594
rect 13970 22542 14196 22594
rect 13916 22540 14196 22542
rect 14700 22932 14756 22942
rect 13916 22530 13972 22540
rect 13356 22418 13412 22428
rect 14476 22484 14532 22494
rect 14476 22390 14532 22428
rect 12908 22318 12910 22370
rect 12962 22318 12964 22370
rect 12908 21812 12964 22318
rect 14028 22372 14084 22382
rect 14028 22278 14084 22316
rect 14700 22370 14756 22876
rect 14700 22318 14702 22370
rect 14754 22318 14756 22370
rect 14700 22306 14756 22318
rect 13916 22260 13972 22270
rect 13916 22166 13972 22204
rect 14364 22258 14420 22270
rect 14364 22206 14366 22258
rect 14418 22206 14420 22258
rect 13132 21812 13188 21822
rect 12908 21810 13188 21812
rect 12908 21758 13134 21810
rect 13186 21758 13188 21810
rect 12908 21756 13188 21758
rect 13132 21746 13188 21756
rect 14364 21700 14420 22206
rect 14812 21924 14868 23102
rect 14924 23156 14980 23166
rect 14924 22594 14980 23100
rect 14924 22542 14926 22594
rect 14978 22542 14980 22594
rect 14924 22530 14980 22542
rect 15036 23044 15092 23324
rect 15372 23154 15428 23166
rect 15372 23102 15374 23154
rect 15426 23102 15428 23154
rect 15148 23044 15204 23054
rect 15036 23042 15204 23044
rect 15036 22990 15150 23042
rect 15202 22990 15204 23042
rect 15036 22988 15204 22990
rect 14812 21858 14868 21868
rect 14924 21700 14980 21710
rect 15036 21700 15092 22988
rect 15148 22978 15204 22988
rect 15260 23042 15316 23054
rect 15260 22990 15262 23042
rect 15314 22990 15316 23042
rect 15260 22596 15316 22990
rect 15372 22932 15428 23102
rect 15820 23044 15876 23054
rect 15820 22950 15876 22988
rect 15372 22866 15428 22876
rect 15260 22530 15316 22540
rect 15484 22708 15540 22718
rect 15148 22372 15204 22382
rect 15148 22278 15204 22316
rect 15484 22370 15540 22652
rect 15484 22318 15486 22370
rect 15538 22318 15540 22370
rect 15484 22306 15540 22318
rect 15708 22596 15764 22606
rect 15708 22370 15764 22540
rect 15708 22318 15710 22370
rect 15762 22318 15764 22370
rect 15708 22306 15764 22318
rect 15820 22372 15876 22382
rect 15820 22278 15876 22316
rect 16156 22370 16212 22382
rect 16156 22318 16158 22370
rect 16210 22318 16212 22370
rect 15932 22148 15988 22158
rect 15932 22146 16100 22148
rect 15932 22094 15934 22146
rect 15986 22094 16100 22146
rect 15932 22092 16100 22094
rect 15932 22082 15988 22092
rect 15708 21924 15764 21934
rect 15708 21812 15764 21868
rect 15708 21810 15988 21812
rect 15708 21758 15710 21810
rect 15762 21758 15988 21810
rect 15708 21756 15988 21758
rect 15708 21746 15764 21756
rect 14364 21698 15092 21700
rect 14364 21646 14926 21698
rect 14978 21646 15092 21698
rect 14364 21644 15092 21646
rect 4284 21588 4340 21598
rect 4284 21494 4340 21532
rect 9884 21588 9940 21598
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4172 20962 4228 20972
rect 1932 20850 1988 20860
rect 9884 20692 9940 21532
rect 9884 19906 9940 20636
rect 13244 21364 13300 21374
rect 12012 20244 12068 20254
rect 12012 20130 12068 20188
rect 12012 20078 12014 20130
rect 12066 20078 12068 20130
rect 12012 20066 12068 20078
rect 13244 20130 13300 21308
rect 13468 20692 13524 20702
rect 13468 20598 13524 20636
rect 13580 20578 13636 20590
rect 13580 20526 13582 20578
rect 13634 20526 13636 20578
rect 13580 20188 13636 20526
rect 14140 20578 14196 20590
rect 14140 20526 14142 20578
rect 14194 20526 14196 20578
rect 14140 20188 14196 20526
rect 14588 20580 14644 20590
rect 14476 20244 14532 20282
rect 13580 20132 14084 20188
rect 14140 20132 14308 20188
rect 14476 20178 14532 20188
rect 13244 20078 13246 20130
rect 13298 20078 13300 20130
rect 13244 20066 13300 20078
rect 12796 20020 12852 20030
rect 12796 20018 12964 20020
rect 12796 19966 12798 20018
rect 12850 19966 12964 20018
rect 12796 19964 12964 19966
rect 12796 19954 12852 19964
rect 9884 19854 9886 19906
rect 9938 19854 9940 19906
rect 9884 19842 9940 19854
rect 12124 19908 12180 19918
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 1932 19346 1988 19358
rect 1932 19294 1934 19346
rect 1986 19294 1988 19346
rect 1932 18900 1988 19294
rect 9996 19346 10052 19358
rect 9996 19294 9998 19346
rect 10050 19294 10052 19346
rect 4284 19236 4340 19246
rect 4284 19142 4340 19180
rect 9996 19236 10052 19294
rect 12124 19346 12180 19852
rect 12124 19294 12126 19346
rect 12178 19294 12180 19346
rect 12124 19282 12180 19294
rect 9996 19170 10052 19180
rect 12908 19234 12964 19964
rect 13580 20018 13636 20030
rect 13580 19966 13582 20018
rect 13634 19966 13636 20018
rect 13356 19908 13412 19918
rect 13356 19814 13412 19852
rect 12908 19182 12910 19234
rect 12962 19182 12964 19234
rect 12908 19012 12964 19182
rect 12908 18946 12964 18956
rect 13132 19236 13188 19246
rect 1932 18834 1988 18844
rect 12908 18562 12964 18574
rect 12908 18510 12910 18562
rect 12962 18510 12964 18562
rect 4284 18452 4340 18462
rect 4284 18358 4340 18396
rect 12908 18452 12964 18510
rect 12908 18386 12964 18396
rect 13132 18450 13188 19180
rect 13580 19234 13636 19966
rect 13804 20018 13860 20030
rect 13804 19966 13806 20018
rect 13858 19966 13860 20018
rect 13804 19684 13860 19966
rect 14028 20018 14084 20132
rect 14028 19966 14030 20018
rect 14082 19966 14084 20018
rect 14028 19954 14084 19966
rect 13804 19618 13860 19628
rect 13580 19182 13582 19234
rect 13634 19182 13636 19234
rect 13580 19170 13636 19182
rect 13804 19236 13860 19246
rect 13804 19122 13860 19180
rect 13804 19070 13806 19122
rect 13858 19070 13860 19122
rect 13804 19058 13860 19070
rect 13916 19122 13972 19134
rect 13916 19070 13918 19122
rect 13970 19070 13972 19122
rect 13916 18788 13972 19070
rect 14252 19012 14308 20132
rect 14476 20018 14532 20030
rect 14476 19966 14478 20018
rect 14530 19966 14532 20018
rect 14364 19012 14420 19022
rect 14252 18956 14364 19012
rect 13916 18722 13972 18732
rect 13132 18398 13134 18450
rect 13186 18398 13188 18450
rect 13132 18386 13188 18398
rect 13916 18452 13972 18462
rect 14364 18452 14420 18956
rect 14476 18788 14532 19966
rect 14588 20018 14644 20524
rect 14588 19966 14590 20018
rect 14642 19966 14644 20018
rect 14588 19954 14644 19966
rect 14812 20020 14868 20030
rect 14924 20020 14980 21644
rect 15260 21588 15316 21598
rect 15260 21494 15316 21532
rect 15820 21586 15876 21598
rect 15820 21534 15822 21586
rect 15874 21534 15876 21586
rect 15708 21364 15764 21374
rect 15708 21270 15764 21308
rect 15820 21252 15876 21534
rect 15820 21186 15876 21196
rect 15036 21140 15092 21150
rect 15036 20130 15092 21084
rect 15036 20078 15038 20130
rect 15090 20078 15092 20130
rect 15036 20066 15092 20078
rect 15596 21028 15652 21038
rect 15596 20690 15652 20972
rect 15932 20804 15988 21756
rect 15596 20638 15598 20690
rect 15650 20638 15652 20690
rect 14812 20018 14980 20020
rect 14812 19966 14814 20018
rect 14866 19966 14980 20018
rect 14812 19964 14980 19966
rect 14812 19954 14868 19964
rect 15484 19012 15540 19022
rect 15484 18918 15540 18956
rect 14476 18722 14532 18732
rect 15148 18788 15204 18798
rect 15204 18732 15316 18788
rect 15148 18722 15204 18732
rect 13916 18450 14420 18452
rect 13916 18398 13918 18450
rect 13970 18398 14420 18450
rect 13916 18396 14420 18398
rect 1932 18228 1988 18238
rect 1932 18134 1988 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 13580 16100 13636 16110
rect 13916 16100 13972 18396
rect 14700 18340 14756 18350
rect 14700 18338 15204 18340
rect 14700 18286 14702 18338
rect 14754 18286 15204 18338
rect 14700 18284 15204 18286
rect 14700 18274 14756 18284
rect 15148 17890 15204 18284
rect 15148 17838 15150 17890
rect 15202 17838 15204 17890
rect 15148 17826 15204 17838
rect 15260 17668 15316 18732
rect 15484 17892 15540 17902
rect 15596 17892 15652 20638
rect 15820 20802 15988 20804
rect 15820 20750 15934 20802
rect 15986 20750 15988 20802
rect 15820 20748 15988 20750
rect 15708 20580 15764 20590
rect 15708 20486 15764 20524
rect 15820 20242 15876 20748
rect 15932 20738 15988 20748
rect 16044 21588 16100 22092
rect 15820 20190 15822 20242
rect 15874 20190 15876 20242
rect 15820 19234 15876 20190
rect 16044 19908 16100 21532
rect 16156 21252 16212 22318
rect 16156 21186 16212 21196
rect 16492 22370 16548 23436
rect 17388 23378 17444 23884
rect 17388 23326 17390 23378
rect 17442 23326 17444 23378
rect 17388 23314 17444 23326
rect 16492 22318 16494 22370
rect 16546 22318 16548 22370
rect 16492 21028 16548 22318
rect 16716 22258 16772 22270
rect 16716 22206 16718 22258
rect 16770 22206 16772 22258
rect 16716 21924 16772 22206
rect 16716 21858 16772 21868
rect 17388 22260 17444 22270
rect 16492 20962 16548 20972
rect 16940 21140 16996 21150
rect 16940 20802 16996 21084
rect 16940 20750 16942 20802
rect 16994 20750 16996 20802
rect 16940 20738 16996 20750
rect 17164 20914 17220 20926
rect 17164 20862 17166 20914
rect 17218 20862 17220 20914
rect 16156 20692 16212 20702
rect 16156 20690 16324 20692
rect 16156 20638 16158 20690
rect 16210 20638 16324 20690
rect 16156 20636 16324 20638
rect 16156 20626 16212 20636
rect 16268 20132 16324 20636
rect 16492 20132 16548 20142
rect 16268 20130 16548 20132
rect 16268 20078 16494 20130
rect 16546 20078 16548 20130
rect 16268 20076 16548 20078
rect 16156 20020 16212 20030
rect 16156 19926 16212 19964
rect 16044 19842 16100 19852
rect 15820 19182 15822 19234
rect 15874 19182 15876 19234
rect 15820 19170 15876 19182
rect 15932 19684 15988 19694
rect 15708 19012 15764 19022
rect 15708 18918 15764 18956
rect 15484 17890 15652 17892
rect 15484 17838 15486 17890
rect 15538 17838 15652 17890
rect 15484 17836 15652 17838
rect 15484 17826 15540 17836
rect 15036 17612 15316 17668
rect 14924 16996 14980 17006
rect 15036 16996 15092 17612
rect 14924 16994 15092 16996
rect 14924 16942 14926 16994
rect 14978 16942 15092 16994
rect 14924 16940 15092 16942
rect 15260 17442 15316 17454
rect 15260 17390 15262 17442
rect 15314 17390 15316 17442
rect 14924 16930 14980 16940
rect 15260 16882 15316 17390
rect 15260 16830 15262 16882
rect 15314 16830 15316 16882
rect 15036 16770 15092 16782
rect 15036 16718 15038 16770
rect 15090 16718 15092 16770
rect 15036 16324 15092 16718
rect 15260 16660 15316 16830
rect 15260 16594 15316 16604
rect 15484 16882 15540 16894
rect 15484 16830 15486 16882
rect 15538 16830 15540 16882
rect 15484 16772 15540 16830
rect 14252 16268 15092 16324
rect 14252 16210 14308 16268
rect 14252 16158 14254 16210
rect 14306 16158 14308 16210
rect 14252 16146 14308 16158
rect 13580 16098 13972 16100
rect 13580 16046 13582 16098
rect 13634 16046 13972 16098
rect 13580 16044 13972 16046
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 13580 13748 13636 16044
rect 15484 14756 15540 16716
rect 15596 14756 15652 14766
rect 15484 14754 15652 14756
rect 15484 14702 15598 14754
rect 15650 14702 15652 14754
rect 15484 14700 15652 14702
rect 15596 14532 15652 14700
rect 15820 14756 15876 14766
rect 15932 14756 15988 19628
rect 16492 19124 16548 20076
rect 16828 20132 16884 20142
rect 16828 20038 16884 20076
rect 16492 19058 16548 19068
rect 17052 19012 17108 19022
rect 16940 19010 17108 19012
rect 16940 18958 17054 19010
rect 17106 18958 17108 19010
rect 16940 18956 17108 18958
rect 16828 18340 16884 18350
rect 16828 18246 16884 18284
rect 16716 17444 16772 17454
rect 16604 16996 16660 17006
rect 16604 16902 16660 16940
rect 16492 16772 16548 16782
rect 16492 16678 16548 16716
rect 16380 16660 16436 16670
rect 16380 16566 16436 16604
rect 16380 16212 16436 16222
rect 16716 16212 16772 17388
rect 16380 16210 16772 16212
rect 16380 16158 16382 16210
rect 16434 16158 16772 16210
rect 16380 16156 16772 16158
rect 16828 16212 16884 16222
rect 16940 16212 16996 18956
rect 17052 18946 17108 18956
rect 17164 19012 17220 20862
rect 17164 17442 17220 18956
rect 17164 17390 17166 17442
rect 17218 17390 17220 17442
rect 17164 17332 17220 17390
rect 17388 17444 17444 22204
rect 17500 22146 17556 25340
rect 17612 24948 17668 24958
rect 17612 24854 17668 24892
rect 18508 24948 18564 24958
rect 18508 24854 18564 24892
rect 18620 24948 18676 24958
rect 18732 24948 18788 25566
rect 18844 26290 18900 26302
rect 18844 26238 18846 26290
rect 18898 26238 18900 26290
rect 18844 25508 18900 26238
rect 19068 26292 19124 26302
rect 19068 26198 19124 26236
rect 18844 25442 18900 25452
rect 19180 25284 19236 25294
rect 19180 25190 19236 25228
rect 18620 24946 18788 24948
rect 18620 24894 18622 24946
rect 18674 24894 18788 24946
rect 18620 24892 18788 24894
rect 19404 24948 19460 26460
rect 19628 26404 19684 26460
rect 19852 26514 20244 26516
rect 19852 26462 19854 26514
rect 19906 26462 20244 26514
rect 19852 26460 20244 26462
rect 20524 26516 20580 27132
rect 20636 26740 20692 27694
rect 20748 27746 21364 27748
rect 20748 27694 21198 27746
rect 21250 27694 21364 27746
rect 20748 27692 21364 27694
rect 20748 27186 20804 27692
rect 21196 27682 21252 27692
rect 20748 27134 20750 27186
rect 20802 27134 20804 27186
rect 20748 27122 20804 27134
rect 20636 26674 20692 26684
rect 20524 26460 21028 26516
rect 19852 26450 19908 26460
rect 19740 26404 19796 26414
rect 19628 26402 19796 26404
rect 19628 26350 19742 26402
rect 19794 26350 19796 26402
rect 19628 26348 19796 26350
rect 19740 26338 19796 26348
rect 20412 26404 20468 26414
rect 20412 26402 20580 26404
rect 20412 26350 20414 26402
rect 20466 26350 20580 26402
rect 20412 26348 20580 26350
rect 20412 26338 20468 26348
rect 19516 26292 19572 26302
rect 20076 26292 20132 26302
rect 20300 26292 20356 26302
rect 19516 26290 19684 26292
rect 19516 26238 19518 26290
rect 19570 26238 19684 26290
rect 19516 26236 19684 26238
rect 19516 26226 19572 26236
rect 18620 24882 18676 24892
rect 19404 24882 19460 24892
rect 18844 24722 18900 24734
rect 18844 24670 18846 24722
rect 18898 24670 18900 24722
rect 17724 24612 17780 24622
rect 17724 24518 17780 24556
rect 18732 24612 18788 24622
rect 18732 24518 18788 24556
rect 18844 23940 18900 24670
rect 18844 23874 18900 23884
rect 19068 24722 19124 24734
rect 19068 24670 19070 24722
rect 19122 24670 19124 24722
rect 18732 23828 18788 23838
rect 18508 23772 18732 23828
rect 17500 22094 17502 22146
rect 17554 22094 17556 22146
rect 17500 22082 17556 22094
rect 17612 23154 17668 23166
rect 17612 23102 17614 23154
rect 17666 23102 17668 23154
rect 17612 20132 17668 23102
rect 17724 22596 17780 22606
rect 17724 21026 17780 22540
rect 17724 20974 17726 21026
rect 17778 20974 17780 21026
rect 17724 20962 17780 20974
rect 18172 21586 18228 21598
rect 18172 21534 18174 21586
rect 18226 21534 18228 21586
rect 18172 20916 18228 21534
rect 18172 20850 18228 20860
rect 17948 20804 18004 20814
rect 17948 20802 18116 20804
rect 17948 20750 17950 20802
rect 18002 20750 18116 20802
rect 17948 20748 18116 20750
rect 17948 20738 18004 20748
rect 17668 20076 17780 20132
rect 17612 20066 17668 20076
rect 17612 18452 17668 18462
rect 17500 18450 17668 18452
rect 17500 18398 17614 18450
rect 17666 18398 17668 18450
rect 17500 18396 17668 18398
rect 17500 17780 17556 18396
rect 17612 18386 17668 18396
rect 17724 18338 17780 20076
rect 18060 20020 18116 20748
rect 18060 18564 18116 19964
rect 18172 20018 18228 20030
rect 18172 19966 18174 20018
rect 18226 19966 18228 20018
rect 18172 19012 18228 19966
rect 18172 18946 18228 18956
rect 18508 19684 18564 23772
rect 18732 23762 18788 23772
rect 19068 23714 19124 24670
rect 19628 24050 19684 26236
rect 20076 26290 20356 26292
rect 20076 26238 20078 26290
rect 20130 26238 20302 26290
rect 20354 26238 20356 26290
rect 20076 26236 20356 26238
rect 20076 26226 20132 26236
rect 20300 26226 20356 26236
rect 20412 26180 20468 26190
rect 20412 26066 20468 26124
rect 20412 26014 20414 26066
rect 20466 26014 20468 26066
rect 20412 26002 20468 26014
rect 20076 25508 20132 25518
rect 20076 25414 20132 25452
rect 20188 25396 20244 25406
rect 20188 25302 20244 25340
rect 20412 25396 20468 25406
rect 20412 25302 20468 25340
rect 20524 25172 20580 26348
rect 20972 26402 21028 26460
rect 20972 26350 20974 26402
rect 21026 26350 21028 26402
rect 20972 26338 21028 26350
rect 20860 26292 20916 26302
rect 20860 26198 20916 26236
rect 21308 26290 21364 27692
rect 22988 27076 23044 27086
rect 23324 27076 23380 27086
rect 22988 27074 23268 27076
rect 22988 27022 22990 27074
rect 23042 27022 23268 27074
rect 22988 27020 23268 27022
rect 22988 27010 23044 27020
rect 23100 26852 23156 26862
rect 21308 26238 21310 26290
rect 21362 26238 21364 26290
rect 21308 25284 21364 26238
rect 21980 26850 23156 26852
rect 21980 26798 23102 26850
rect 23154 26798 23156 26850
rect 21980 26796 23156 26798
rect 21868 25732 21924 25742
rect 21980 25732 22036 26796
rect 23100 26786 23156 26796
rect 22092 26180 22148 26190
rect 22092 26178 22260 26180
rect 22092 26126 22094 26178
rect 22146 26126 22260 26178
rect 22092 26124 22260 26126
rect 22092 26114 22148 26124
rect 21868 25730 22036 25732
rect 21868 25678 21870 25730
rect 21922 25678 22036 25730
rect 21868 25676 22036 25678
rect 21868 25666 21924 25676
rect 22204 25618 22260 26124
rect 22204 25566 22206 25618
rect 22258 25566 22260 25618
rect 22204 25554 22260 25566
rect 21420 25508 21476 25518
rect 21420 25396 21476 25452
rect 21756 25506 21812 25518
rect 21756 25454 21758 25506
rect 21810 25454 21812 25506
rect 21420 25394 21700 25396
rect 21420 25342 21422 25394
rect 21474 25342 21700 25394
rect 21420 25340 21700 25342
rect 21420 25330 21476 25340
rect 21308 25218 21364 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20524 25106 20580 25116
rect 19836 25050 20100 25060
rect 19628 23998 19630 24050
rect 19682 23998 19684 24050
rect 19628 23986 19684 23998
rect 19404 23940 19460 23950
rect 19068 23662 19070 23714
rect 19122 23662 19124 23714
rect 19068 23650 19124 23662
rect 19180 23938 19460 23940
rect 19180 23886 19406 23938
rect 19458 23886 19460 23938
rect 19180 23884 19460 23886
rect 19180 23378 19236 23884
rect 19404 23874 19460 23884
rect 19516 23940 19572 23950
rect 19180 23326 19182 23378
rect 19234 23326 19236 23378
rect 19180 23314 19236 23326
rect 19292 23716 19348 23726
rect 19292 23714 19460 23716
rect 19292 23662 19294 23714
rect 19346 23662 19460 23714
rect 19292 23660 19460 23662
rect 19068 23044 19124 23054
rect 19292 23044 19348 23660
rect 19404 23380 19460 23660
rect 19516 23604 19572 23884
rect 19740 23938 19796 23950
rect 19740 23886 19742 23938
rect 19794 23886 19796 23938
rect 19740 23828 19796 23886
rect 20076 23940 20132 23950
rect 20076 23846 20132 23884
rect 19740 23762 19796 23772
rect 19516 23548 19684 23604
rect 19516 23380 19572 23390
rect 19404 23378 19572 23380
rect 19404 23326 19518 23378
rect 19570 23326 19572 23378
rect 19404 23324 19572 23326
rect 19516 23314 19572 23324
rect 19068 22950 19124 22988
rect 19180 22988 19348 23044
rect 19180 21812 19236 22988
rect 19180 21746 19236 21756
rect 19292 22820 19348 22830
rect 18620 21588 18676 21598
rect 19292 21588 19348 22764
rect 19628 22596 19684 23548
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 21532 23380 21588 23390
rect 21532 23286 21588 23324
rect 20412 23266 20468 23278
rect 20412 23214 20414 23266
rect 20466 23214 20468 23266
rect 19740 23154 19796 23166
rect 19740 23102 19742 23154
rect 19794 23102 19796 23154
rect 19740 22820 19796 23102
rect 19740 22754 19796 22764
rect 20300 23044 20356 23054
rect 19852 22596 19908 22606
rect 19628 22594 19908 22596
rect 19628 22542 19854 22594
rect 19906 22542 19908 22594
rect 19628 22540 19908 22542
rect 19852 22530 19908 22540
rect 20300 22482 20356 22988
rect 20412 22932 20468 23214
rect 20412 22866 20468 22876
rect 20636 23154 20692 23166
rect 20636 23102 20638 23154
rect 20690 23102 20692 23154
rect 20300 22430 20302 22482
rect 20354 22430 20356 22482
rect 20300 22418 20356 22430
rect 18620 21586 19348 21588
rect 18620 21534 18622 21586
rect 18674 21534 19348 21586
rect 18620 21532 19348 21534
rect 18620 21522 18676 21532
rect 18620 21140 18676 21150
rect 18620 20578 18676 21084
rect 18732 20914 18788 21532
rect 19292 21474 19348 21532
rect 19292 21422 19294 21474
rect 19346 21422 19348 21474
rect 19292 21410 19348 21422
rect 19404 22370 19460 22382
rect 19404 22318 19406 22370
rect 19458 22318 19460 22370
rect 19404 21700 19460 22318
rect 19516 22370 19572 22382
rect 19516 22318 19518 22370
rect 19570 22318 19572 22370
rect 19516 22260 19572 22318
rect 19516 22194 19572 22204
rect 19740 22370 19796 22382
rect 19740 22318 19742 22370
rect 19794 22318 19796 22370
rect 19740 22148 19796 22318
rect 20636 22370 20692 23102
rect 21532 22484 21588 22494
rect 20636 22318 20638 22370
rect 20690 22318 20692 22370
rect 19740 22082 19796 22092
rect 20188 22258 20244 22270
rect 20188 22206 20190 22258
rect 20242 22206 20244 22258
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20188 21924 20244 22206
rect 20524 22258 20580 22270
rect 20524 22206 20526 22258
rect 20578 22206 20580 22258
rect 20524 22148 20580 22206
rect 20524 22082 20580 22092
rect 20188 21700 20244 21868
rect 20188 21644 20468 21700
rect 19068 21364 19124 21374
rect 18956 21362 19124 21364
rect 18956 21310 19070 21362
rect 19122 21310 19124 21362
rect 18956 21308 19124 21310
rect 18956 21028 19012 21308
rect 19068 21298 19124 21308
rect 19404 21140 19460 21644
rect 19516 21588 19572 21598
rect 20076 21588 20132 21598
rect 19516 21586 20244 21588
rect 19516 21534 19518 21586
rect 19570 21534 20078 21586
rect 20130 21534 20244 21586
rect 19516 21532 20244 21534
rect 19516 21522 19572 21532
rect 20076 21522 20132 21532
rect 18956 20962 19012 20972
rect 19292 21084 19460 21140
rect 19740 21364 19796 21374
rect 18732 20862 18734 20914
rect 18786 20862 18788 20914
rect 18732 20850 18788 20862
rect 19180 20916 19236 20926
rect 18620 20526 18622 20578
rect 18674 20526 18676 20578
rect 18620 20514 18676 20526
rect 19180 20802 19236 20860
rect 19180 20750 19182 20802
rect 19234 20750 19236 20802
rect 18620 20020 18676 20030
rect 18620 19926 18676 19964
rect 19068 20020 19124 20030
rect 18732 19908 18788 19918
rect 18732 19814 18788 19852
rect 18284 18564 18340 18574
rect 18060 18562 18340 18564
rect 18060 18510 18286 18562
rect 18338 18510 18340 18562
rect 18060 18508 18340 18510
rect 17948 18452 18004 18462
rect 17948 18358 18004 18396
rect 17724 18286 17726 18338
rect 17778 18286 17780 18338
rect 17724 18274 17780 18286
rect 18284 18228 18340 18508
rect 18284 18162 18340 18172
rect 18508 18116 18564 19628
rect 19068 18676 19124 19964
rect 18844 18620 19124 18676
rect 18620 18452 18676 18462
rect 18620 18358 18676 18396
rect 18508 18050 18564 18060
rect 17500 17666 17556 17724
rect 18508 17780 18564 17790
rect 18508 17686 18564 17724
rect 17500 17614 17502 17666
rect 17554 17614 17556 17666
rect 17500 17602 17556 17614
rect 18620 17554 18676 17566
rect 18620 17502 18622 17554
rect 18674 17502 18676 17554
rect 17836 17444 17892 17454
rect 17388 17388 17668 17444
rect 17164 17276 17556 17332
rect 16828 16210 16996 16212
rect 16828 16158 16830 16210
rect 16882 16158 16996 16210
rect 16828 16156 16996 16158
rect 16380 16146 16436 16156
rect 16492 15316 16548 15326
rect 16828 15316 16884 16156
rect 17388 15426 17444 15438
rect 17388 15374 17390 15426
rect 17442 15374 17444 15426
rect 16492 15222 16548 15260
rect 16716 15260 16884 15316
rect 16940 15316 16996 15326
rect 16492 15092 16548 15102
rect 15820 14754 15988 14756
rect 15820 14702 15822 14754
rect 15874 14702 15988 14754
rect 15820 14700 15988 14702
rect 16044 15090 16548 15092
rect 16044 15038 16494 15090
rect 16546 15038 16548 15090
rect 16044 15036 16548 15038
rect 15820 14690 15876 14700
rect 15596 14466 15652 14476
rect 16044 14530 16100 15036
rect 16492 15026 16548 15036
rect 16044 14478 16046 14530
rect 16098 14478 16100 14530
rect 16044 14466 16100 14478
rect 14700 14420 14756 14430
rect 14700 13858 14756 14364
rect 15484 14420 15540 14430
rect 15484 14326 15540 14364
rect 14700 13806 14702 13858
rect 14754 13806 14756 13858
rect 14700 13794 14756 13806
rect 16604 14308 16660 14318
rect 14028 13748 14084 13758
rect 13580 13746 14084 13748
rect 13580 13694 14030 13746
rect 14082 13694 14084 13746
rect 13580 13692 14084 13694
rect 14028 13524 14084 13692
rect 14028 13458 14084 13468
rect 15932 13524 15988 13534
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 15932 12962 15988 13468
rect 16604 13074 16660 14252
rect 16716 13524 16772 15260
rect 16828 15092 16884 15102
rect 16828 14998 16884 15036
rect 16940 14756 16996 15260
rect 17388 15316 17444 15374
rect 17500 15316 17556 17276
rect 17612 16996 17668 17388
rect 17836 17350 17892 17388
rect 18172 17442 18228 17454
rect 18172 17390 18174 17442
rect 18226 17390 18228 17442
rect 17612 16930 17668 16940
rect 18172 16996 18228 17390
rect 18620 17444 18676 17502
rect 18844 17444 18900 18620
rect 18956 18452 19012 18462
rect 18956 17668 19012 18396
rect 19068 18450 19124 18620
rect 19068 18398 19070 18450
rect 19122 18398 19124 18450
rect 19068 18386 19124 18398
rect 19180 18340 19236 20750
rect 19180 18274 19236 18284
rect 18956 17612 19124 17668
rect 18956 17444 19012 17454
rect 18844 17442 19012 17444
rect 18844 17390 18958 17442
rect 19010 17390 19012 17442
rect 18844 17388 19012 17390
rect 18620 17378 18676 17388
rect 18172 16930 18228 16940
rect 17836 16884 17892 16894
rect 17612 15316 17668 15326
rect 17500 15314 17668 15316
rect 17500 15262 17614 15314
rect 17666 15262 17668 15314
rect 17500 15260 17668 15262
rect 17388 15250 17444 15260
rect 17612 15250 17668 15260
rect 16716 13458 16772 13468
rect 16828 14700 16996 14756
rect 16828 13634 16884 14700
rect 17836 14642 17892 16828
rect 18956 16772 19012 17388
rect 19068 17106 19124 17612
rect 19068 17054 19070 17106
rect 19122 17054 19124 17106
rect 19068 17042 19124 17054
rect 19292 17554 19348 21084
rect 19740 21028 19796 21308
rect 19404 21026 19796 21028
rect 19404 20974 19742 21026
rect 19794 20974 19796 21026
rect 19404 20972 19796 20974
rect 19404 20690 19460 20972
rect 19740 20962 19796 20972
rect 19852 21252 19908 21262
rect 19852 20914 19908 21196
rect 19852 20862 19854 20914
rect 19906 20862 19908 20914
rect 19852 20850 19908 20862
rect 20188 20916 20244 21532
rect 20412 21140 20468 21644
rect 20524 21476 20580 21486
rect 20636 21476 20692 22318
rect 21308 22482 21588 22484
rect 21308 22430 21534 22482
rect 21586 22430 21588 22482
rect 21308 22428 21588 22430
rect 20524 21474 20692 21476
rect 20524 21422 20526 21474
rect 20578 21422 20692 21474
rect 20524 21420 20692 21422
rect 20972 22148 21028 22158
rect 20524 21364 20580 21420
rect 20524 21298 20580 21308
rect 20412 21084 20804 21140
rect 20188 20860 20692 20916
rect 19404 20638 19406 20690
rect 19458 20638 19460 20690
rect 19404 20626 19460 20638
rect 20076 20802 20132 20814
rect 20076 20750 20078 20802
rect 20130 20750 20132 20802
rect 20076 20580 20132 20750
rect 20636 20802 20692 20860
rect 20636 20750 20638 20802
rect 20690 20750 20692 20802
rect 20412 20692 20468 20702
rect 20412 20598 20468 20636
rect 20636 20580 20692 20750
rect 20076 20524 20356 20580
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20130 20244 20142
rect 20188 20078 20190 20130
rect 20242 20078 20244 20130
rect 19852 20020 19908 20030
rect 19852 19926 19908 19964
rect 20188 19908 20244 20078
rect 20300 20132 20356 20524
rect 20636 20514 20692 20524
rect 20300 20066 20356 20076
rect 20748 19908 20804 21084
rect 20972 20692 21028 22092
rect 21308 21588 21364 22428
rect 21532 22418 21588 22428
rect 21644 22260 21700 25340
rect 21756 25172 21812 25454
rect 21756 23604 21812 25116
rect 22092 25506 22148 25518
rect 22092 25454 22094 25506
rect 22146 25454 22148 25506
rect 22092 24724 22148 25454
rect 22652 25506 22708 25518
rect 22652 25454 22654 25506
rect 22706 25454 22708 25506
rect 22316 25394 22372 25406
rect 22316 25342 22318 25394
rect 22370 25342 22372 25394
rect 22316 24948 22372 25342
rect 22652 25284 22708 25454
rect 22652 25218 22708 25228
rect 22316 24892 22820 24948
rect 22652 24724 22708 24734
rect 22092 24722 22708 24724
rect 22092 24670 22654 24722
rect 22706 24670 22708 24722
rect 22092 24668 22708 24670
rect 22764 24724 22820 24892
rect 22876 24724 22932 24734
rect 23212 24724 23268 27020
rect 23324 26982 23380 27020
rect 24220 27076 24276 27086
rect 24220 26178 24276 27020
rect 24556 27076 24612 37998
rect 26796 37490 26852 38556
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 26796 37438 26798 37490
rect 26850 37438 26852 37490
rect 26796 37426 26852 37438
rect 25788 37266 25844 37278
rect 25788 37214 25790 37266
rect 25842 37214 25844 37266
rect 25788 31948 25844 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 24556 27010 24612 27020
rect 25564 31892 25844 31948
rect 24220 26126 24222 26178
rect 24274 26126 24276 26178
rect 24220 26114 24276 26126
rect 24668 26178 24724 26190
rect 24668 26126 24670 26178
rect 24722 26126 24724 26178
rect 23436 25394 23492 25406
rect 23436 25342 23438 25394
rect 23490 25342 23492 25394
rect 23436 24946 23492 25342
rect 23436 24894 23438 24946
rect 23490 24894 23492 24946
rect 23436 24882 23492 24894
rect 23548 25284 23604 25294
rect 22764 24722 22932 24724
rect 22764 24670 22878 24722
rect 22930 24670 22932 24722
rect 22764 24668 22932 24670
rect 22428 24500 22484 24510
rect 21756 23548 22036 23604
rect 21532 22204 21700 22260
rect 21756 23154 21812 23166
rect 21756 23102 21758 23154
rect 21810 23102 21812 23154
rect 21532 21698 21588 22204
rect 21532 21646 21534 21698
rect 21586 21646 21588 21698
rect 21532 21634 21588 21646
rect 21644 21924 21700 21934
rect 21308 21586 21476 21588
rect 21308 21534 21310 21586
rect 21362 21534 21476 21586
rect 21308 21532 21476 21534
rect 21308 21522 21364 21532
rect 21308 20804 21364 20814
rect 20972 20626 21028 20636
rect 21084 20748 21308 20804
rect 21420 20804 21476 21532
rect 21644 21586 21700 21868
rect 21644 21534 21646 21586
rect 21698 21534 21700 21586
rect 21644 21522 21700 21534
rect 21756 21588 21812 23102
rect 21868 22820 21924 22830
rect 21868 22370 21924 22764
rect 21868 22318 21870 22370
rect 21922 22318 21924 22370
rect 21868 22306 21924 22318
rect 21980 21588 22036 23548
rect 22428 22482 22484 24444
rect 22540 23380 22596 24668
rect 22652 24658 22708 24668
rect 22540 23314 22596 23324
rect 22652 23938 22708 23950
rect 22652 23886 22654 23938
rect 22706 23886 22708 23938
rect 22428 22430 22430 22482
rect 22482 22430 22484 22482
rect 22428 22418 22484 22430
rect 22316 22370 22372 22382
rect 22316 22318 22318 22370
rect 22370 22318 22372 22370
rect 22316 22260 22372 22318
rect 22316 21924 22372 22204
rect 22316 21858 22372 21868
rect 22092 21588 22148 21598
rect 21756 21532 21924 21588
rect 21980 21532 22092 21588
rect 21868 21364 21924 21532
rect 22092 21522 22148 21532
rect 21868 21308 22036 21364
rect 21420 20748 21700 20804
rect 21084 20130 21140 20748
rect 21308 20710 21364 20748
rect 21420 20580 21476 20590
rect 21420 20132 21476 20524
rect 21084 20078 21086 20130
rect 21138 20078 21140 20130
rect 21084 20066 21140 20078
rect 21308 20130 21476 20132
rect 21308 20078 21422 20130
rect 21474 20078 21476 20130
rect 21308 20076 21476 20078
rect 20188 19852 20804 19908
rect 21308 19122 21364 20076
rect 21420 20066 21476 20076
rect 21532 20132 21588 20142
rect 21532 20038 21588 20076
rect 21308 19070 21310 19122
rect 21362 19070 21364 19122
rect 21308 19058 21364 19070
rect 21532 19234 21588 19246
rect 21532 19182 21534 19234
rect 21586 19182 21588 19234
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19852 18676 19908 18686
rect 21532 18676 21588 19182
rect 19516 18564 19572 18574
rect 19516 18450 19572 18508
rect 19516 18398 19518 18450
rect 19570 18398 19572 18450
rect 19516 17668 19572 18398
rect 19628 18452 19684 18462
rect 19628 17890 19684 18396
rect 19628 17838 19630 17890
rect 19682 17838 19684 17890
rect 19628 17826 19684 17838
rect 19852 17778 19908 18620
rect 20860 18620 21588 18676
rect 20860 18450 20916 18620
rect 20860 18398 20862 18450
rect 20914 18398 20916 18450
rect 20860 18386 20916 18398
rect 21084 18450 21140 18462
rect 21084 18398 21086 18450
rect 21138 18398 21140 18450
rect 19964 18338 20020 18350
rect 19964 18286 19966 18338
rect 20018 18286 20020 18338
rect 19964 18116 20020 18286
rect 20636 18340 20692 18350
rect 20636 18246 20692 18284
rect 20300 18228 20356 18238
rect 20300 18226 20580 18228
rect 20300 18174 20302 18226
rect 20354 18174 20580 18226
rect 20300 18172 20580 18174
rect 20300 18162 20356 18172
rect 19964 18050 20020 18060
rect 19852 17726 19854 17778
rect 19906 17726 19908 17778
rect 19852 17714 19908 17726
rect 20524 18004 20580 18172
rect 21084 18004 21140 18398
rect 20524 17948 21140 18004
rect 21420 18450 21476 18462
rect 21420 18398 21422 18450
rect 21474 18398 21476 18450
rect 21420 18228 21476 18398
rect 19516 17612 19684 17668
rect 19292 17502 19294 17554
rect 19346 17502 19348 17554
rect 19180 16884 19236 16894
rect 19180 16790 19236 16828
rect 18956 16706 19012 16716
rect 17836 14590 17838 14642
rect 17890 14590 17892 14642
rect 17836 14578 17892 14590
rect 18284 15316 18340 15326
rect 16940 14532 16996 14542
rect 16940 14418 16996 14476
rect 16940 14366 16942 14418
rect 16994 14366 16996 14418
rect 16940 14354 16996 14366
rect 17164 14420 17220 14430
rect 17164 14326 17220 14364
rect 17052 14308 17108 14318
rect 17052 14214 17108 14252
rect 18284 13970 18340 15260
rect 18844 15092 18900 15102
rect 18284 13918 18286 13970
rect 18338 13918 18340 13970
rect 18284 13906 18340 13918
rect 18396 14420 18452 14430
rect 18396 13970 18452 14364
rect 18396 13918 18398 13970
rect 18450 13918 18452 13970
rect 18396 13906 18452 13918
rect 18508 13746 18564 13758
rect 18508 13694 18510 13746
rect 18562 13694 18564 13746
rect 16828 13582 16830 13634
rect 16882 13582 16884 13634
rect 16604 13022 16606 13074
rect 16658 13022 16660 13074
rect 16604 13010 16660 13022
rect 15932 12910 15934 12962
rect 15986 12910 15988 12962
rect 15932 12898 15988 12910
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 16828 8428 16884 13582
rect 17500 13634 17556 13646
rect 17500 13582 17502 13634
rect 17554 13582 17556 13634
rect 17500 13524 17556 13582
rect 17500 13458 17556 13468
rect 18508 13076 18564 13694
rect 18844 13746 18900 15036
rect 19292 15092 19348 17502
rect 19516 17444 19572 17454
rect 19516 17106 19572 17388
rect 19516 17054 19518 17106
rect 19570 17054 19572 17106
rect 19516 17042 19572 17054
rect 19628 17108 19684 17612
rect 20524 17666 20580 17948
rect 20524 17614 20526 17666
rect 20578 17614 20580 17666
rect 20524 17602 20580 17614
rect 19852 17444 19908 17482
rect 19852 17378 19908 17388
rect 20300 17442 20356 17454
rect 20300 17390 20302 17442
rect 20354 17390 20356 17442
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 17052 20132 17108
rect 20076 16882 20132 17052
rect 20076 16830 20078 16882
rect 20130 16830 20132 16882
rect 20076 16818 20132 16830
rect 20300 16660 20356 17390
rect 20524 17444 20580 17454
rect 20412 16994 20468 17006
rect 20412 16942 20414 16994
rect 20466 16942 20468 16994
rect 20412 16772 20468 16942
rect 20412 16706 20468 16716
rect 20300 16212 20356 16604
rect 19964 16156 20356 16212
rect 19964 16098 20020 16156
rect 19964 16046 19966 16098
rect 20018 16046 20020 16098
rect 19964 16034 20020 16046
rect 20076 16044 20356 16100
rect 20076 15874 20132 16044
rect 20076 15822 20078 15874
rect 20130 15822 20132 15874
rect 20076 15810 20132 15822
rect 20188 15876 20244 15886
rect 20188 15782 20244 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20300 15148 20356 16044
rect 20524 16098 20580 17388
rect 20636 16884 20692 16894
rect 20636 16790 20692 16828
rect 21420 16882 21476 18172
rect 21420 16830 21422 16882
rect 21474 16830 21476 16882
rect 21420 16818 21476 16830
rect 20524 16046 20526 16098
rect 20578 16046 20580 16098
rect 20524 16034 20580 16046
rect 21532 15204 21588 18620
rect 21644 18674 21700 20748
rect 21868 20132 21924 20142
rect 21868 20038 21924 20076
rect 21980 19908 22036 21308
rect 22652 21140 22708 23886
rect 22876 22932 22932 24668
rect 23100 24668 23268 24724
rect 23436 24724 23492 24734
rect 23100 24500 23156 24668
rect 23436 24630 23492 24668
rect 23100 24434 23156 24444
rect 23212 24500 23268 24510
rect 23212 24498 23380 24500
rect 23212 24446 23214 24498
rect 23266 24446 23380 24498
rect 23212 24444 23380 24446
rect 23212 24434 23268 24444
rect 22876 22866 22932 22876
rect 22988 22260 23044 22270
rect 22988 22166 23044 22204
rect 23212 22258 23268 22270
rect 23212 22206 23214 22258
rect 23266 22206 23268 22258
rect 23212 22148 23268 22206
rect 23212 22082 23268 22092
rect 23324 22146 23380 24444
rect 23548 24052 23604 25228
rect 24668 25284 24724 26126
rect 25564 25618 25620 31892
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 27580 26292 27636 26302
rect 25788 26180 25844 26190
rect 25564 25566 25566 25618
rect 25618 25566 25620 25618
rect 24668 25218 24724 25228
rect 25340 25284 25396 25294
rect 24556 25172 24612 25182
rect 24556 24946 24612 25116
rect 24556 24894 24558 24946
rect 24610 24894 24612 24946
rect 24556 24882 24612 24894
rect 25340 24948 25396 25228
rect 25564 25172 25620 25566
rect 25564 25106 25620 25116
rect 25676 26178 25844 26180
rect 25676 26126 25790 26178
rect 25842 26126 25844 26178
rect 25676 26124 25844 26126
rect 25676 24948 25732 26124
rect 25788 26114 25844 26124
rect 26684 25620 26740 25630
rect 26460 25618 26740 25620
rect 26460 25566 26686 25618
rect 26738 25566 26740 25618
rect 26460 25564 26740 25566
rect 26236 25396 26292 25406
rect 26236 25302 26292 25340
rect 26348 25394 26404 25406
rect 26348 25342 26350 25394
rect 26402 25342 26404 25394
rect 25340 24946 25732 24948
rect 25340 24894 25342 24946
rect 25394 24894 25732 24946
rect 25340 24892 25732 24894
rect 25340 24882 25396 24892
rect 24444 24724 24500 24734
rect 24444 24630 24500 24668
rect 25676 24722 25732 24892
rect 25676 24670 25678 24722
rect 25730 24670 25732 24722
rect 24332 24500 24388 24510
rect 24332 24406 24388 24444
rect 23548 24050 24052 24052
rect 23548 23998 23550 24050
rect 23602 23998 24052 24050
rect 23548 23996 24052 23998
rect 23548 23986 23604 23996
rect 23996 22370 24052 23996
rect 25676 23604 25732 24670
rect 25900 25282 25956 25294
rect 25900 25230 25902 25282
rect 25954 25230 25956 25282
rect 25900 24500 25956 25230
rect 26124 25284 26180 25294
rect 26124 25190 26180 25228
rect 25900 24434 25956 24444
rect 25676 23538 25732 23548
rect 24444 23044 24500 23054
rect 23996 22318 23998 22370
rect 24050 22318 24052 22370
rect 23996 22306 24052 22318
rect 24108 23042 24500 23044
rect 24108 22990 24446 23042
rect 24498 22990 24500 23042
rect 24108 22988 24500 22990
rect 23324 22094 23326 22146
rect 23378 22094 23380 22146
rect 22764 21980 23156 22036
rect 22764 21698 22820 21980
rect 23100 21924 23156 21980
rect 23324 21924 23380 22094
rect 23100 21868 23380 21924
rect 23548 22258 23604 22270
rect 23548 22206 23550 22258
rect 23602 22206 23604 22258
rect 23212 21700 23268 21868
rect 22764 21646 22766 21698
rect 22818 21646 22820 21698
rect 22764 21634 22820 21646
rect 23100 21644 23268 21700
rect 23436 21700 23492 21710
rect 22204 20132 22260 20142
rect 22204 20038 22260 20076
rect 22540 20020 22596 20030
rect 22428 20018 22596 20020
rect 22428 19966 22542 20018
rect 22594 19966 22596 20018
rect 22428 19964 22596 19966
rect 22428 19908 22484 19964
rect 22540 19954 22596 19964
rect 21980 19852 22484 19908
rect 21644 18622 21646 18674
rect 21698 18622 21700 18674
rect 21644 18564 21700 18622
rect 22428 18676 22484 19852
rect 22428 18610 22484 18620
rect 21644 18498 21700 18508
rect 22540 18562 22596 18574
rect 22540 18510 22542 18562
rect 22594 18510 22596 18562
rect 21756 18452 21812 18462
rect 21756 18358 21812 18396
rect 22316 18452 22372 18462
rect 22316 18358 22372 18396
rect 22540 18340 22596 18510
rect 22540 17444 22596 18284
rect 22652 17666 22708 21084
rect 22988 21588 23044 21598
rect 22876 20132 22932 20142
rect 22876 20038 22932 20076
rect 22652 17614 22654 17666
rect 22706 17614 22708 17666
rect 22652 17602 22708 17614
rect 22764 20020 22820 20030
rect 22540 17378 22596 17388
rect 21644 16994 21700 17006
rect 21644 16942 21646 16994
rect 21698 16942 21700 16994
rect 21644 16772 21700 16942
rect 21644 15876 21700 16716
rect 22764 16660 22820 19964
rect 22988 19908 23044 21532
rect 22876 19852 23044 19908
rect 22876 18340 22932 19852
rect 23100 19460 23156 21644
rect 23324 21588 23380 21598
rect 23212 21532 23324 21588
rect 23212 21474 23268 21532
rect 23324 21522 23380 21532
rect 23436 21586 23492 21644
rect 23436 21534 23438 21586
rect 23490 21534 23492 21586
rect 23436 21522 23492 21534
rect 23212 21422 23214 21474
rect 23266 21422 23268 21474
rect 23212 21410 23268 21422
rect 23324 21364 23380 21374
rect 23212 20130 23268 20142
rect 23212 20078 23214 20130
rect 23266 20078 23268 20130
rect 23212 20020 23268 20078
rect 23324 20132 23380 21308
rect 23548 21364 23604 22206
rect 24108 22148 24164 22988
rect 24444 22978 24500 22988
rect 24556 22932 24612 22942
rect 24556 22930 24836 22932
rect 24556 22878 24558 22930
rect 24610 22878 24836 22930
rect 24556 22876 24836 22878
rect 24556 22866 24612 22876
rect 24780 22482 24836 22876
rect 24780 22430 24782 22482
rect 24834 22430 24836 22482
rect 24780 22418 24836 22430
rect 23772 22092 24164 22148
rect 24332 22372 24388 22382
rect 23772 21810 23828 22092
rect 23772 21758 23774 21810
rect 23826 21758 23828 21810
rect 23772 21746 23828 21758
rect 23884 21756 24164 21812
rect 23660 21700 23716 21710
rect 23660 21606 23716 21644
rect 23548 21298 23604 21308
rect 23436 21140 23492 21150
rect 23492 21084 23604 21140
rect 23436 21074 23492 21084
rect 23548 20914 23604 21084
rect 23548 20862 23550 20914
rect 23602 20862 23604 20914
rect 23548 20850 23604 20862
rect 23436 20132 23492 20142
rect 23324 20130 23492 20132
rect 23324 20078 23438 20130
rect 23490 20078 23492 20130
rect 23324 20076 23492 20078
rect 23436 20066 23492 20076
rect 23212 19954 23268 19964
rect 23772 20020 23828 20030
rect 23884 20020 23940 21756
rect 24108 21698 24164 21756
rect 24332 21810 24388 22316
rect 26348 22260 26404 25342
rect 26460 24834 26516 25564
rect 26684 25554 26740 25564
rect 27580 25618 27636 26236
rect 27580 25566 27582 25618
rect 27634 25566 27636 25618
rect 27580 25554 27636 25566
rect 28588 26292 28644 26302
rect 27468 25284 27524 25294
rect 27468 25190 27524 25228
rect 26460 24782 26462 24834
rect 26514 24782 26516 24834
rect 26460 24770 26516 24782
rect 28588 24610 28644 26236
rect 37660 26292 37716 26302
rect 37660 26198 37716 26236
rect 40012 26066 40068 26078
rect 40012 26014 40014 26066
rect 40066 26014 40068 26066
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 40012 25620 40068 26014
rect 40012 25554 40068 25564
rect 28588 24558 28590 24610
rect 28642 24558 28644 24610
rect 28588 24546 28644 24558
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 27132 23492 27188 23502
rect 27132 23380 27188 23436
rect 27132 23378 27524 23380
rect 27132 23326 27134 23378
rect 27186 23326 27524 23378
rect 27132 23324 27524 23326
rect 25564 22148 25620 22158
rect 24332 21758 24334 21810
rect 24386 21758 24388 21810
rect 24332 21746 24388 21758
rect 25228 21812 25284 21822
rect 25228 21718 25284 21756
rect 24108 21646 24110 21698
rect 24162 21646 24164 21698
rect 24108 21634 24164 21646
rect 25564 21698 25620 22092
rect 26236 21812 26292 21822
rect 26348 21812 26404 22204
rect 26908 22484 26964 22494
rect 26908 22036 26964 22428
rect 26908 21970 26964 21980
rect 26236 21810 26404 21812
rect 26236 21758 26238 21810
rect 26290 21758 26404 21810
rect 26236 21756 26404 21758
rect 26796 21812 26852 21822
rect 27132 21812 27188 23324
rect 27468 23154 27524 23324
rect 27468 23102 27470 23154
rect 27522 23102 27524 23154
rect 27468 23090 27524 23102
rect 37660 23154 37716 23166
rect 37660 23102 37662 23154
rect 37714 23102 37716 23154
rect 28252 23044 28308 23054
rect 28252 22950 28308 22988
rect 29260 23044 29316 23054
rect 28028 22596 28084 22606
rect 27244 22372 27300 22382
rect 27244 22278 27300 22316
rect 27580 22372 27636 22382
rect 27580 22278 27636 22316
rect 28028 22372 28084 22540
rect 28476 22594 28532 22606
rect 28476 22542 28478 22594
rect 28530 22542 28532 22594
rect 28364 22372 28420 22382
rect 28028 22370 28420 22372
rect 28028 22318 28030 22370
rect 28082 22318 28366 22370
rect 28418 22318 28420 22370
rect 28028 22316 28420 22318
rect 28028 22306 28084 22316
rect 28364 22306 28420 22316
rect 28476 22372 28532 22542
rect 29260 22482 29316 22988
rect 29260 22430 29262 22482
rect 29314 22430 29316 22482
rect 29260 22418 29316 22430
rect 30380 23042 30436 23054
rect 30380 22990 30382 23042
rect 30434 22990 30436 23042
rect 28700 22372 28756 22382
rect 28476 22306 28532 22316
rect 28588 22316 28700 22372
rect 27804 22148 27860 22158
rect 27804 22054 27860 22092
rect 27916 22146 27972 22158
rect 27916 22094 27918 22146
rect 27970 22094 27972 22146
rect 26796 21810 27188 21812
rect 26796 21758 26798 21810
rect 26850 21758 27188 21810
rect 26796 21756 27188 21758
rect 26236 21746 26292 21756
rect 26796 21746 26852 21756
rect 25564 21646 25566 21698
rect 25618 21646 25620 21698
rect 23996 21588 24052 21598
rect 23996 20132 24052 21532
rect 24332 21586 24388 21598
rect 24332 21534 24334 21586
rect 24386 21534 24388 21586
rect 24332 21476 24388 21534
rect 24668 21588 24724 21598
rect 24668 21494 24724 21532
rect 24332 21410 24388 21420
rect 23996 20038 24052 20076
rect 24108 21364 24164 21374
rect 24108 20130 24164 21308
rect 24108 20078 24110 20130
rect 24162 20078 24164 20130
rect 24108 20066 24164 20078
rect 23772 20018 23940 20020
rect 23772 19966 23774 20018
rect 23826 19966 23940 20018
rect 23772 19964 23940 19966
rect 23324 19906 23380 19918
rect 23324 19854 23326 19906
rect 23378 19854 23380 19906
rect 23212 19460 23268 19470
rect 23100 19458 23268 19460
rect 23100 19406 23214 19458
rect 23266 19406 23268 19458
rect 23100 19404 23268 19406
rect 23212 19394 23268 19404
rect 22988 19234 23044 19246
rect 22988 19182 22990 19234
rect 23042 19182 23044 19234
rect 22988 18452 23044 19182
rect 22988 18386 23044 18396
rect 22876 18274 22932 18284
rect 23212 18228 23268 18238
rect 23212 17106 23268 18172
rect 23212 17054 23214 17106
rect 23266 17054 23268 17106
rect 23212 17042 23268 17054
rect 23100 16996 23156 17006
rect 23100 16902 23156 16940
rect 22764 16594 22820 16604
rect 23212 16100 23268 16110
rect 23324 16100 23380 19854
rect 23772 19908 23828 19964
rect 23772 19842 23828 19852
rect 24108 19796 24164 19806
rect 24108 19702 24164 19740
rect 25564 19236 25620 21646
rect 26012 21698 26068 21710
rect 26012 21646 26014 21698
rect 26066 21646 26068 21698
rect 25900 21588 25956 21598
rect 25900 21494 25956 21532
rect 26012 21476 26068 21646
rect 26012 21410 26068 21420
rect 27132 21586 27188 21756
rect 27916 21698 27972 22094
rect 28476 22148 28532 22158
rect 28588 22148 28644 22316
rect 28700 22306 28756 22316
rect 30044 22372 30100 22382
rect 29148 22260 29204 22270
rect 29148 22166 29204 22204
rect 28476 22146 28644 22148
rect 28476 22094 28478 22146
rect 28530 22094 28644 22146
rect 28476 22092 28644 22094
rect 29372 22148 29428 22158
rect 28476 22082 28532 22092
rect 29372 22054 29428 22092
rect 29596 22146 29652 22158
rect 29596 22094 29598 22146
rect 29650 22094 29652 22146
rect 27916 21646 27918 21698
rect 27970 21646 27972 21698
rect 27916 21634 27972 21646
rect 27132 21534 27134 21586
rect 27186 21534 27188 21586
rect 27132 20914 27188 21534
rect 27132 20862 27134 20914
rect 27186 20862 27188 20914
rect 27132 20850 27188 20862
rect 29484 20804 29540 20814
rect 29596 20804 29652 22094
rect 30044 21474 30100 22316
rect 30044 21422 30046 21474
rect 30098 21422 30100 21474
rect 30044 21410 30100 21422
rect 30380 21588 30436 22990
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 37660 22596 37716 23102
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 37660 22530 37716 22540
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 37660 22372 37716 22382
rect 37660 22278 37716 22316
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 29484 20802 29652 20804
rect 29484 20750 29486 20802
rect 29538 20750 29652 20802
rect 29484 20748 29652 20750
rect 29484 20738 29540 20748
rect 29148 20690 29204 20702
rect 29148 20638 29150 20690
rect 29202 20638 29204 20690
rect 25900 19796 25956 19806
rect 25676 19236 25732 19246
rect 25564 19180 25676 19236
rect 23548 19010 23604 19022
rect 23548 18958 23550 19010
rect 23602 18958 23604 19010
rect 23548 18452 23604 18958
rect 25676 18674 25732 19180
rect 25676 18622 25678 18674
rect 25730 18622 25732 18674
rect 25676 18610 25732 18622
rect 25900 19012 25956 19740
rect 27916 19236 27972 19246
rect 27916 19142 27972 19180
rect 29148 19234 29204 20638
rect 29260 20692 29316 20702
rect 29260 20598 29316 20636
rect 30380 20692 30436 21532
rect 37660 21588 37716 21598
rect 37660 21494 37716 21532
rect 40012 21588 40068 21598
rect 40012 21474 40068 21532
rect 40012 21422 40014 21474
rect 40066 21422 40068 21474
rect 40012 21410 40068 21422
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 30380 20626 30436 20636
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 40012 19346 40068 19358
rect 40012 19294 40014 19346
rect 40066 19294 40068 19346
rect 29148 19182 29150 19234
rect 29202 19182 29204 19234
rect 29036 19124 29092 19134
rect 29148 19124 29204 19182
rect 37660 19236 37716 19246
rect 37660 19142 37716 19180
rect 29092 19068 29204 19124
rect 29036 19058 29092 19068
rect 25900 18674 25956 18956
rect 25900 18622 25902 18674
rect 25954 18622 25956 18674
rect 25900 18610 25956 18622
rect 27356 19012 27412 19022
rect 23548 18386 23604 18396
rect 25452 18452 25508 18462
rect 25452 18358 25508 18396
rect 27020 18450 27076 18462
rect 27020 18398 27022 18450
rect 27074 18398 27076 18450
rect 25788 18338 25844 18350
rect 25788 18286 25790 18338
rect 25842 18286 25844 18338
rect 25228 18228 25284 18238
rect 25228 18134 25284 18172
rect 23436 17668 23492 17678
rect 23436 16994 23492 17612
rect 23436 16942 23438 16994
rect 23490 16942 23492 16994
rect 23436 16930 23492 16942
rect 23996 17668 24052 17678
rect 23548 16882 23604 16894
rect 23548 16830 23550 16882
rect 23602 16830 23604 16882
rect 23548 16772 23604 16830
rect 23604 16716 23716 16772
rect 23548 16706 23604 16716
rect 23436 16660 23492 16670
rect 23436 16212 23492 16604
rect 23436 16156 23604 16212
rect 23212 16098 23380 16100
rect 23212 16046 23214 16098
rect 23266 16046 23380 16098
rect 23212 16044 23380 16046
rect 23212 16034 23268 16044
rect 22876 15988 22932 15998
rect 23436 15988 23492 15998
rect 21644 15810 21700 15820
rect 22652 15986 22932 15988
rect 22652 15934 22878 15986
rect 22930 15934 22932 15986
rect 22652 15932 22932 15934
rect 21644 15204 21700 15214
rect 21532 15148 21644 15204
rect 19292 15026 19348 15036
rect 19964 15092 20356 15148
rect 21644 15138 21700 15148
rect 22316 15092 22372 15102
rect 19964 14642 20020 15092
rect 19964 14590 19966 14642
rect 20018 14590 20020 14642
rect 19964 14578 20020 14590
rect 20748 14532 20804 14542
rect 20748 14438 20804 14476
rect 21420 14532 21476 14542
rect 21420 14306 21476 14476
rect 22316 14530 22372 15036
rect 22316 14478 22318 14530
rect 22370 14478 22372 14530
rect 22316 14466 22372 14478
rect 22652 14530 22708 15932
rect 22876 15922 22932 15932
rect 23324 15986 23492 15988
rect 23324 15934 23438 15986
rect 23490 15934 23492 15986
rect 23324 15932 23492 15934
rect 22988 15874 23044 15886
rect 22988 15822 22990 15874
rect 23042 15822 23044 15874
rect 22876 15540 22932 15550
rect 22652 14478 22654 14530
rect 22706 14478 22708 14530
rect 22652 14466 22708 14478
rect 22764 15538 22932 15540
rect 22764 15486 22878 15538
rect 22930 15486 22932 15538
rect 22764 15484 22932 15486
rect 21420 14254 21422 14306
rect 21474 14254 21476 14306
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 18844 13694 18846 13746
rect 18898 13694 18900 13746
rect 18844 13682 18900 13694
rect 19292 13524 19348 13534
rect 18732 13076 18788 13086
rect 18508 13074 18788 13076
rect 18508 13022 18734 13074
rect 18786 13022 18788 13074
rect 18508 13020 18788 13022
rect 18732 8428 18788 13020
rect 19292 13076 19348 13468
rect 21420 13076 21476 14254
rect 22428 14306 22484 14318
rect 22428 14254 22430 14306
rect 22482 14254 22484 14306
rect 21756 13746 21812 13758
rect 21756 13694 21758 13746
rect 21810 13694 21812 13746
rect 21756 13524 21812 13694
rect 21532 13076 21588 13086
rect 21756 13076 21812 13468
rect 21420 13020 21532 13076
rect 21588 13020 21812 13076
rect 22428 13076 22484 14254
rect 22540 13860 22596 13870
rect 22764 13860 22820 15484
rect 22876 15474 22932 15484
rect 22876 15092 22932 15102
rect 22876 14642 22932 15036
rect 22876 14590 22878 14642
rect 22930 14590 22932 14642
rect 22876 14578 22932 14590
rect 22540 13858 22820 13860
rect 22540 13806 22542 13858
rect 22594 13806 22820 13858
rect 22540 13804 22820 13806
rect 22540 13794 22596 13804
rect 19292 12982 19348 13020
rect 21532 12962 21588 13020
rect 22428 13010 22484 13020
rect 21532 12910 21534 12962
rect 21586 12910 21588 12962
rect 21532 12898 21588 12910
rect 22316 12852 22372 12862
rect 22988 12852 23044 15822
rect 23324 15428 23380 15932
rect 23436 15922 23492 15932
rect 23100 15372 23380 15428
rect 23436 15428 23492 15438
rect 23548 15428 23604 16156
rect 23436 15426 23548 15428
rect 23436 15374 23438 15426
rect 23490 15374 23548 15426
rect 23436 15372 23548 15374
rect 23100 15316 23156 15372
rect 23436 15362 23492 15372
rect 23548 15334 23604 15372
rect 23660 15428 23716 16716
rect 23996 16210 24052 17612
rect 23996 16158 23998 16210
rect 24050 16158 24052 16210
rect 23996 16146 24052 16158
rect 25788 16212 25844 18286
rect 26684 18340 26740 18350
rect 27020 18340 27076 18398
rect 26684 18338 27076 18340
rect 26684 18286 26686 18338
rect 26738 18286 27076 18338
rect 26684 18284 27076 18286
rect 26684 18274 26740 18284
rect 26348 17556 26404 17566
rect 26796 17556 26852 18284
rect 27356 17666 27412 18956
rect 27692 19012 27748 19022
rect 27692 18918 27748 18956
rect 27804 19010 27860 19022
rect 27804 18958 27806 19010
rect 27858 18958 27860 19010
rect 27804 18564 27860 18958
rect 28140 19012 28196 19022
rect 28140 18918 28196 18956
rect 27804 18508 27972 18564
rect 27804 18340 27860 18350
rect 27468 18338 27860 18340
rect 27468 18286 27806 18338
rect 27858 18286 27860 18338
rect 27468 18284 27860 18286
rect 27468 17778 27524 18284
rect 27804 18274 27860 18284
rect 27468 17726 27470 17778
rect 27522 17726 27524 17778
rect 27468 17714 27524 17726
rect 27356 17614 27358 17666
rect 27410 17614 27412 17666
rect 27356 17602 27412 17614
rect 26908 17556 26964 17566
rect 26796 17500 26908 17556
rect 26348 17462 26404 17500
rect 26908 16770 26964 17500
rect 27580 17442 27636 17454
rect 27580 17390 27582 17442
rect 27634 17390 27636 17442
rect 26908 16718 26910 16770
rect 26962 16718 26964 16770
rect 26124 16212 26180 16222
rect 25788 16210 26180 16212
rect 25788 16158 26126 16210
rect 26178 16158 26180 16210
rect 25788 16156 26180 16158
rect 26124 16146 26180 16156
rect 26908 16100 26964 16718
rect 27244 16882 27300 16894
rect 27244 16830 27246 16882
rect 27298 16830 27300 16882
rect 27244 16100 27300 16830
rect 27356 16100 27412 16110
rect 26796 16098 27412 16100
rect 26796 16046 26910 16098
rect 26962 16046 27358 16098
rect 27410 16046 27412 16098
rect 26796 16044 27412 16046
rect 23996 15428 24052 15438
rect 23660 15426 24052 15428
rect 23660 15374 23662 15426
rect 23714 15374 23998 15426
rect 24050 15374 24052 15426
rect 23660 15372 24052 15374
rect 23660 15362 23716 15372
rect 23996 15362 24052 15372
rect 25004 15428 25060 15438
rect 23100 15222 23156 15260
rect 24332 15314 24388 15326
rect 24332 15262 24334 15314
rect 24386 15262 24388 15314
rect 23212 15204 23268 15242
rect 23212 15138 23268 15148
rect 24108 15204 24164 15242
rect 24108 15138 24164 15148
rect 24332 13636 24388 15262
rect 25004 14642 25060 15372
rect 25004 14590 25006 14642
rect 25058 14590 25060 14642
rect 25004 14578 25060 14590
rect 25676 14532 25732 14542
rect 26236 14532 26292 14542
rect 26796 14532 26852 16044
rect 26908 16034 26964 16044
rect 27356 16034 27412 16044
rect 27580 15428 27636 17390
rect 27916 16996 27972 18508
rect 28028 17666 28084 17678
rect 28028 17614 28030 17666
rect 28082 17614 28084 17666
rect 28028 17444 28084 17614
rect 29148 17666 29204 19068
rect 29260 19124 29316 19134
rect 29260 19030 29316 19068
rect 30156 19124 30212 19134
rect 29484 19012 29540 19022
rect 29484 18918 29540 18956
rect 29148 17614 29150 17666
rect 29202 17614 29204 17666
rect 29148 17602 29204 17614
rect 29932 18338 29988 18350
rect 29932 18286 29934 18338
rect 29986 18286 29988 18338
rect 29260 17556 29316 17566
rect 29260 17462 29316 17500
rect 29932 17556 29988 18286
rect 29932 17490 29988 17500
rect 28028 17378 28084 17388
rect 29484 17444 29540 17454
rect 29484 17350 29540 17388
rect 28028 16996 28084 17006
rect 27916 16994 28084 16996
rect 27916 16942 28030 16994
rect 28082 16942 28084 16994
rect 27916 16940 28084 16942
rect 28028 16930 28084 16940
rect 30156 16770 30212 19068
rect 40012 18900 40068 19294
rect 40012 18834 40068 18844
rect 37884 18450 37940 18462
rect 37884 18398 37886 18450
rect 37938 18398 37940 18450
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 37660 17668 37716 17678
rect 37660 17574 37716 17612
rect 37884 17556 37940 18398
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 37884 17490 37940 17500
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 40012 17556 40068 17726
rect 40012 17490 40068 17500
rect 30156 16718 30158 16770
rect 30210 16718 30212 16770
rect 30156 16706 30212 16718
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 27580 15362 27636 15372
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 25676 14530 26852 14532
rect 25676 14478 25678 14530
rect 25730 14478 26238 14530
rect 26290 14478 26852 14530
rect 25676 14476 26852 14478
rect 24668 13636 24724 13646
rect 24332 13580 24668 13636
rect 24668 13542 24724 13580
rect 25340 13636 25396 13646
rect 25676 13636 25732 14476
rect 26236 14466 26292 14476
rect 25340 13634 25732 13636
rect 25340 13582 25342 13634
rect 25394 13582 25732 13634
rect 25340 13580 25732 13582
rect 25788 13636 25844 13646
rect 25004 13524 25060 13534
rect 25340 13524 25396 13580
rect 25060 13468 25396 13524
rect 24444 13076 24500 13086
rect 24500 13020 24612 13076
rect 24444 12982 24500 13020
rect 22316 12850 23044 12852
rect 22316 12798 22318 12850
rect 22370 12798 23044 12850
rect 22316 12796 23044 12798
rect 22316 12786 22372 12796
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 16828 8372 17108 8428
rect 18732 8372 19124 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 17052 3554 17108 8372
rect 19068 4338 19124 8372
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19068 4286 19070 4338
rect 19122 4286 19124 4338
rect 19068 4274 19124 4286
rect 17052 3502 17054 3554
rect 17106 3502 17108 3554
rect 17052 3490 17108 3502
rect 18844 4116 18900 4126
rect 16828 3444 16884 3454
rect 16828 800 16884 3388
rect 18060 3444 18116 3454
rect 18060 3330 18116 3388
rect 18060 3278 18062 3330
rect 18114 3278 18116 3330
rect 18060 3266 18116 3278
rect 18844 800 18900 4060
rect 20076 4116 20132 4126
rect 20076 4022 20132 4060
rect 24220 4116 24276 4126
rect 23548 3668 23604 3678
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 23548 800 23604 3612
rect 24220 800 24276 4060
rect 24556 3554 24612 13020
rect 25004 13074 25060 13468
rect 25004 13022 25006 13074
rect 25058 13022 25060 13074
rect 25004 13010 25060 13022
rect 25788 8428 25844 13580
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 25564 8372 25844 8428
rect 25564 4338 25620 8372
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 25564 4286 25566 4338
rect 25618 4286 25620 4338
rect 25564 4274 25620 4286
rect 26236 4116 26292 4126
rect 26236 4022 26292 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 35980 3332 36036 3342
rect 35644 3330 36036 3332
rect 35644 3278 35982 3330
rect 36034 3278 36036 3330
rect 35644 3276 36036 3278
rect 35644 800 35700 3276
rect 35980 3266 36036 3276
rect 16800 0 16912 800
rect 18816 0 18928 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 35616 0 35728 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 16156 37436 16212 37492
rect 15484 36652 15540 36708
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4172 27580 4228 27636
rect 1932 24892 1988 24948
rect 1932 22930 1988 22932
rect 1932 22878 1934 22930
rect 1934 22878 1986 22930
rect 1986 22878 1988 22930
rect 1932 22876 1988 22878
rect 1932 22482 1988 22484
rect 1932 22430 1934 22482
rect 1934 22430 1986 22482
rect 1986 22430 1988 22482
rect 1932 22428 1988 22430
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 14924 27020 14980 27076
rect 13916 26460 13972 26516
rect 13244 25228 13300 25284
rect 14028 25228 14084 25284
rect 4284 24556 4340 24612
rect 11116 24610 11172 24612
rect 11116 24558 11118 24610
rect 11118 24558 11170 24610
rect 11170 24558 11172 24610
rect 11116 24556 11172 24558
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 13244 23996 13300 24052
rect 4284 23154 4340 23156
rect 4284 23102 4286 23154
rect 4286 23102 4338 23154
rect 4338 23102 4340 23154
rect 4284 23100 4340 23102
rect 9996 23100 10052 23156
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 14588 24610 14644 24612
rect 14588 24558 14590 24610
rect 14590 24558 14642 24610
rect 14642 24558 14644 24610
rect 14588 24556 14644 24558
rect 14476 24050 14532 24052
rect 14476 23998 14478 24050
rect 14478 23998 14530 24050
rect 14530 23998 14532 24050
rect 14476 23996 14532 23998
rect 14364 23938 14420 23940
rect 14364 23886 14366 23938
rect 14366 23886 14418 23938
rect 14418 23886 14420 23938
rect 14364 23884 14420 23886
rect 15484 27074 15540 27076
rect 15484 27022 15486 27074
rect 15486 27022 15538 27074
rect 15538 27022 15540 27074
rect 15484 27020 15540 27022
rect 16156 28082 16212 28084
rect 16156 28030 16158 28082
rect 16158 28030 16210 28082
rect 16210 28030 16212 28082
rect 16156 28028 16212 28030
rect 18060 38050 18116 38052
rect 18060 37998 18062 38050
rect 18062 37998 18114 38050
rect 18114 37998 18116 38050
rect 18060 37996 18116 37998
rect 18732 37996 18788 38052
rect 18396 37490 18452 37492
rect 18396 37438 18398 37490
rect 18398 37438 18450 37490
rect 18450 37438 18452 37490
rect 18396 37436 18452 37438
rect 16716 36706 16772 36708
rect 16716 36654 16718 36706
rect 16718 36654 16770 36706
rect 16770 36654 16772 36706
rect 16716 36652 16772 36654
rect 16604 28028 16660 28084
rect 17388 28028 17444 28084
rect 16604 27074 16660 27076
rect 16604 27022 16606 27074
rect 16606 27022 16658 27074
rect 16658 27022 16660 27074
rect 16604 27020 16660 27022
rect 16380 26514 16436 26516
rect 16380 26462 16382 26514
rect 16382 26462 16434 26514
rect 16434 26462 16436 26514
rect 16380 26460 16436 26462
rect 15148 26348 15204 26404
rect 16044 26402 16100 26404
rect 16044 26350 16046 26402
rect 16046 26350 16098 26402
rect 16098 26350 16100 26402
rect 16044 26348 16100 26350
rect 15036 25228 15092 25284
rect 16156 25340 16212 25396
rect 15820 25228 15876 25284
rect 18172 26460 18228 26516
rect 18508 26124 18564 26180
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20860 38220 20916 38276
rect 22092 38274 22148 38276
rect 22092 38222 22094 38274
rect 22094 38222 22146 38274
rect 22146 38222 22148 38274
rect 22092 38220 22148 38222
rect 25564 38556 25620 38612
rect 26796 38556 26852 38612
rect 24220 38220 24276 38276
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 20188 37436 20244 37492
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 21420 37490 21476 37492
rect 21420 37438 21422 37490
rect 21422 37438 21474 37490
rect 21474 37438 21476 37490
rect 21420 37436 21476 37438
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20188 26684 20244 26740
rect 18956 26514 19012 26516
rect 18956 26462 18958 26514
rect 18958 26462 19010 26514
rect 19010 26462 19012 26514
rect 18956 26460 19012 26462
rect 16828 25228 16884 25284
rect 17500 25340 17556 25396
rect 16604 24892 16660 24948
rect 14812 23884 14868 23940
rect 17388 24780 17444 24836
rect 17388 23884 17444 23940
rect 14700 23548 14756 23604
rect 16492 23436 16548 23492
rect 11228 22652 11284 22708
rect 12908 22988 12964 23044
rect 4284 22370 4340 22372
rect 4284 22318 4286 22370
rect 4286 22318 4338 22370
rect 4338 22318 4340 22370
rect 4284 22316 4340 22318
rect 12124 22540 12180 22596
rect 9996 22204 10052 22260
rect 14028 22988 14084 23044
rect 14700 22876 14756 22932
rect 13356 22428 13412 22484
rect 14476 22482 14532 22484
rect 14476 22430 14478 22482
rect 14478 22430 14530 22482
rect 14530 22430 14532 22482
rect 14476 22428 14532 22430
rect 14028 22370 14084 22372
rect 14028 22318 14030 22370
rect 14030 22318 14082 22370
rect 14082 22318 14084 22370
rect 14028 22316 14084 22318
rect 13916 22258 13972 22260
rect 13916 22206 13918 22258
rect 13918 22206 13970 22258
rect 13970 22206 13972 22258
rect 13916 22204 13972 22206
rect 14924 23154 14980 23156
rect 14924 23102 14926 23154
rect 14926 23102 14978 23154
rect 14978 23102 14980 23154
rect 14924 23100 14980 23102
rect 14812 21868 14868 21924
rect 15820 23042 15876 23044
rect 15820 22990 15822 23042
rect 15822 22990 15874 23042
rect 15874 22990 15876 23042
rect 15820 22988 15876 22990
rect 15372 22876 15428 22932
rect 15260 22540 15316 22596
rect 15484 22652 15540 22708
rect 15148 22370 15204 22372
rect 15148 22318 15150 22370
rect 15150 22318 15202 22370
rect 15202 22318 15204 22370
rect 15148 22316 15204 22318
rect 15708 22540 15764 22596
rect 15820 22370 15876 22372
rect 15820 22318 15822 22370
rect 15822 22318 15874 22370
rect 15874 22318 15876 22370
rect 15820 22316 15876 22318
rect 15708 21868 15764 21924
rect 4284 21586 4340 21588
rect 4284 21534 4286 21586
rect 4286 21534 4338 21586
rect 4338 21534 4340 21586
rect 4284 21532 4340 21534
rect 9884 21532 9940 21588
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4172 20972 4228 21028
rect 1932 20860 1988 20916
rect 9884 20636 9940 20692
rect 13244 21308 13300 21364
rect 12012 20188 12068 20244
rect 13468 20690 13524 20692
rect 13468 20638 13470 20690
rect 13470 20638 13522 20690
rect 13522 20638 13524 20690
rect 13468 20636 13524 20638
rect 14588 20524 14644 20580
rect 14476 20242 14532 20244
rect 14476 20190 14478 20242
rect 14478 20190 14530 20242
rect 14530 20190 14532 20242
rect 14476 20188 14532 20190
rect 12124 19852 12180 19908
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4284 19234 4340 19236
rect 4284 19182 4286 19234
rect 4286 19182 4338 19234
rect 4338 19182 4340 19234
rect 4284 19180 4340 19182
rect 9996 19180 10052 19236
rect 13356 19906 13412 19908
rect 13356 19854 13358 19906
rect 13358 19854 13410 19906
rect 13410 19854 13412 19906
rect 13356 19852 13412 19854
rect 12908 18956 12964 19012
rect 13132 19180 13188 19236
rect 1932 18844 1988 18900
rect 4284 18450 4340 18452
rect 4284 18398 4286 18450
rect 4286 18398 4338 18450
rect 4338 18398 4340 18450
rect 4284 18396 4340 18398
rect 12908 18396 12964 18452
rect 13804 19628 13860 19684
rect 13804 19180 13860 19236
rect 14364 19010 14420 19012
rect 14364 18958 14366 19010
rect 14366 18958 14418 19010
rect 14418 18958 14420 19010
rect 14364 18956 14420 18958
rect 13916 18732 13972 18788
rect 15260 21586 15316 21588
rect 15260 21534 15262 21586
rect 15262 21534 15314 21586
rect 15314 21534 15316 21586
rect 15260 21532 15316 21534
rect 15708 21362 15764 21364
rect 15708 21310 15710 21362
rect 15710 21310 15762 21362
rect 15762 21310 15764 21362
rect 15708 21308 15764 21310
rect 15820 21196 15876 21252
rect 15036 21084 15092 21140
rect 15596 20972 15652 21028
rect 15484 19010 15540 19012
rect 15484 18958 15486 19010
rect 15486 18958 15538 19010
rect 15538 18958 15540 19010
rect 15484 18956 15540 18958
rect 14476 18732 14532 18788
rect 15148 18732 15204 18788
rect 1932 18226 1988 18228
rect 1932 18174 1934 18226
rect 1934 18174 1986 18226
rect 1986 18174 1988 18226
rect 1932 18172 1988 18174
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 15708 20578 15764 20580
rect 15708 20526 15710 20578
rect 15710 20526 15762 20578
rect 15762 20526 15764 20578
rect 15708 20524 15764 20526
rect 16044 21532 16100 21588
rect 16156 21196 16212 21252
rect 16716 21868 16772 21924
rect 17388 22258 17444 22260
rect 17388 22206 17390 22258
rect 17390 22206 17442 22258
rect 17442 22206 17444 22258
rect 17388 22204 17444 22206
rect 16492 20972 16548 21028
rect 16940 21084 16996 21140
rect 16156 20018 16212 20020
rect 16156 19966 16158 20018
rect 16158 19966 16210 20018
rect 16210 19966 16212 20018
rect 16156 19964 16212 19966
rect 16044 19852 16100 19908
rect 15932 19628 15988 19684
rect 15708 19010 15764 19012
rect 15708 18958 15710 19010
rect 15710 18958 15762 19010
rect 15762 18958 15764 19010
rect 15708 18956 15764 18958
rect 15260 16604 15316 16660
rect 15484 16716 15540 16772
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 16828 20130 16884 20132
rect 16828 20078 16830 20130
rect 16830 20078 16882 20130
rect 16882 20078 16884 20130
rect 16828 20076 16884 20078
rect 16492 19068 16548 19124
rect 16828 18338 16884 18340
rect 16828 18286 16830 18338
rect 16830 18286 16882 18338
rect 16882 18286 16884 18338
rect 16828 18284 16884 18286
rect 16716 17388 16772 17444
rect 16604 16994 16660 16996
rect 16604 16942 16606 16994
rect 16606 16942 16658 16994
rect 16658 16942 16660 16994
rect 16604 16940 16660 16942
rect 16492 16770 16548 16772
rect 16492 16718 16494 16770
rect 16494 16718 16546 16770
rect 16546 16718 16548 16770
rect 16492 16716 16548 16718
rect 16380 16658 16436 16660
rect 16380 16606 16382 16658
rect 16382 16606 16434 16658
rect 16434 16606 16436 16658
rect 16380 16604 16436 16606
rect 17164 18956 17220 19012
rect 17612 24946 17668 24948
rect 17612 24894 17614 24946
rect 17614 24894 17666 24946
rect 17666 24894 17668 24946
rect 17612 24892 17668 24894
rect 18508 24946 18564 24948
rect 18508 24894 18510 24946
rect 18510 24894 18562 24946
rect 18562 24894 18564 24946
rect 18508 24892 18564 24894
rect 19068 26290 19124 26292
rect 19068 26238 19070 26290
rect 19070 26238 19122 26290
rect 19122 26238 19124 26290
rect 19068 26236 19124 26238
rect 18844 25452 18900 25508
rect 19180 25282 19236 25284
rect 19180 25230 19182 25282
rect 19182 25230 19234 25282
rect 19234 25230 19236 25282
rect 19180 25228 19236 25230
rect 20636 26684 20692 26740
rect 19404 24892 19460 24948
rect 17724 24610 17780 24612
rect 17724 24558 17726 24610
rect 17726 24558 17778 24610
rect 17778 24558 17780 24610
rect 17724 24556 17780 24558
rect 18732 24610 18788 24612
rect 18732 24558 18734 24610
rect 18734 24558 18786 24610
rect 18786 24558 18788 24610
rect 18732 24556 18788 24558
rect 18844 23884 18900 23940
rect 18732 23772 18788 23828
rect 17724 22540 17780 22596
rect 18172 20860 18228 20916
rect 17612 20076 17668 20132
rect 18060 19964 18116 20020
rect 18172 18956 18228 19012
rect 20412 26124 20468 26180
rect 20076 25506 20132 25508
rect 20076 25454 20078 25506
rect 20078 25454 20130 25506
rect 20130 25454 20132 25506
rect 20076 25452 20132 25454
rect 20188 25394 20244 25396
rect 20188 25342 20190 25394
rect 20190 25342 20242 25394
rect 20242 25342 20244 25394
rect 20188 25340 20244 25342
rect 20412 25394 20468 25396
rect 20412 25342 20414 25394
rect 20414 25342 20466 25394
rect 20466 25342 20468 25394
rect 20412 25340 20468 25342
rect 20860 26290 20916 26292
rect 20860 26238 20862 26290
rect 20862 26238 20914 26290
rect 20914 26238 20916 26290
rect 20860 26236 20916 26238
rect 21420 25452 21476 25508
rect 21308 25228 21364 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20524 25116 20580 25172
rect 20044 25060 20100 25062
rect 19516 23884 19572 23940
rect 20076 23938 20132 23940
rect 20076 23886 20078 23938
rect 20078 23886 20130 23938
rect 20130 23886 20132 23938
rect 20076 23884 20132 23886
rect 19740 23772 19796 23828
rect 19068 23042 19124 23044
rect 19068 22990 19070 23042
rect 19070 22990 19122 23042
rect 19122 22990 19124 23042
rect 19068 22988 19124 22990
rect 19180 21756 19236 21812
rect 19292 22764 19348 22820
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 21532 23378 21588 23380
rect 21532 23326 21534 23378
rect 21534 23326 21586 23378
rect 21586 23326 21588 23378
rect 21532 23324 21588 23326
rect 19740 22764 19796 22820
rect 20300 22988 20356 23044
rect 20412 22876 20468 22932
rect 18620 21084 18676 21140
rect 19516 22204 19572 22260
rect 19740 22092 19796 22148
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20524 22092 20580 22148
rect 19404 21644 19460 21700
rect 20188 21868 20244 21924
rect 18956 20972 19012 21028
rect 19740 21308 19796 21364
rect 19180 20860 19236 20916
rect 18620 20018 18676 20020
rect 18620 19966 18622 20018
rect 18622 19966 18674 20018
rect 18674 19966 18676 20018
rect 18620 19964 18676 19966
rect 19068 19964 19124 20020
rect 18732 19906 18788 19908
rect 18732 19854 18734 19906
rect 18734 19854 18786 19906
rect 18786 19854 18788 19906
rect 18732 19852 18788 19854
rect 18508 19628 18564 19684
rect 17948 18450 18004 18452
rect 17948 18398 17950 18450
rect 17950 18398 18002 18450
rect 18002 18398 18004 18450
rect 17948 18396 18004 18398
rect 18284 18172 18340 18228
rect 18620 18450 18676 18452
rect 18620 18398 18622 18450
rect 18622 18398 18674 18450
rect 18674 18398 18676 18450
rect 18620 18396 18676 18398
rect 18508 18060 18564 18116
rect 17500 17724 17556 17780
rect 18508 17778 18564 17780
rect 18508 17726 18510 17778
rect 18510 17726 18562 17778
rect 18562 17726 18564 17778
rect 18508 17724 18564 17726
rect 16492 15314 16548 15316
rect 16492 15262 16494 15314
rect 16494 15262 16546 15314
rect 16546 15262 16548 15314
rect 16492 15260 16548 15262
rect 16940 15260 16996 15316
rect 15596 14476 15652 14532
rect 14700 14364 14756 14420
rect 15484 14418 15540 14420
rect 15484 14366 15486 14418
rect 15486 14366 15538 14418
rect 15538 14366 15540 14418
rect 15484 14364 15540 14366
rect 16604 14252 16660 14308
rect 14028 13468 14084 13524
rect 15932 13468 15988 13524
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 16828 15090 16884 15092
rect 16828 15038 16830 15090
rect 16830 15038 16882 15090
rect 16882 15038 16884 15090
rect 16828 15036 16884 15038
rect 17388 15260 17444 15316
rect 17836 17442 17892 17444
rect 17836 17390 17838 17442
rect 17838 17390 17890 17442
rect 17890 17390 17892 17442
rect 17836 17388 17892 17390
rect 17612 16940 17668 16996
rect 18620 17388 18676 17444
rect 18956 18396 19012 18452
rect 19180 18284 19236 18340
rect 18172 16940 18228 16996
rect 17836 16828 17892 16884
rect 16716 13468 16772 13524
rect 19852 21196 19908 21252
rect 20972 22092 21028 22148
rect 20524 21308 20580 21364
rect 20412 20690 20468 20692
rect 20412 20638 20414 20690
rect 20414 20638 20466 20690
rect 20466 20638 20468 20690
rect 20412 20636 20468 20638
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19852 20018 19908 20020
rect 19852 19966 19854 20018
rect 19854 19966 19906 20018
rect 19906 19966 19908 20018
rect 19852 19964 19908 19966
rect 20636 20524 20692 20580
rect 20300 20076 20356 20132
rect 21756 25116 21812 25172
rect 22652 25228 22708 25284
rect 23324 27074 23380 27076
rect 23324 27022 23326 27074
rect 23326 27022 23378 27074
rect 23378 27022 23380 27074
rect 23324 27020 23380 27022
rect 24220 27020 24276 27076
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 24556 27020 24612 27076
rect 23548 25228 23604 25284
rect 22428 24444 22484 24500
rect 21644 21868 21700 21924
rect 20972 20636 21028 20692
rect 21308 20802 21364 20804
rect 21308 20750 21310 20802
rect 21310 20750 21362 20802
rect 21362 20750 21364 20802
rect 21308 20748 21364 20750
rect 21868 22764 21924 22820
rect 22540 23324 22596 23380
rect 22316 22204 22372 22260
rect 22316 21868 22372 21924
rect 22092 21532 22148 21588
rect 21420 20524 21476 20580
rect 21532 20130 21588 20132
rect 21532 20078 21534 20130
rect 21534 20078 21586 20130
rect 21586 20078 21588 20130
rect 21532 20076 21588 20078
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19852 18620 19908 18676
rect 19516 18508 19572 18564
rect 19628 18396 19684 18452
rect 20636 18338 20692 18340
rect 20636 18286 20638 18338
rect 20638 18286 20690 18338
rect 20690 18286 20692 18338
rect 20636 18284 20692 18286
rect 19964 18060 20020 18116
rect 21420 18172 21476 18228
rect 19180 16882 19236 16884
rect 19180 16830 19182 16882
rect 19182 16830 19234 16882
rect 19234 16830 19236 16882
rect 19180 16828 19236 16830
rect 18956 16716 19012 16772
rect 18284 15260 18340 15316
rect 16940 14476 16996 14532
rect 17164 14418 17220 14420
rect 17164 14366 17166 14418
rect 17166 14366 17218 14418
rect 17218 14366 17220 14418
rect 17164 14364 17220 14366
rect 17052 14306 17108 14308
rect 17052 14254 17054 14306
rect 17054 14254 17106 14306
rect 17106 14254 17108 14306
rect 17052 14252 17108 14254
rect 18844 15036 18900 15092
rect 18396 14364 18452 14420
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 17500 13468 17556 13524
rect 19516 17388 19572 17444
rect 19852 17442 19908 17444
rect 19852 17390 19854 17442
rect 19854 17390 19906 17442
rect 19906 17390 19908 17442
rect 19852 17388 19908 17390
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20524 17388 20580 17444
rect 20412 16716 20468 16772
rect 20300 16604 20356 16660
rect 20188 15874 20244 15876
rect 20188 15822 20190 15874
rect 20190 15822 20242 15874
rect 20242 15822 20244 15874
rect 20188 15820 20244 15822
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20636 16882 20692 16884
rect 20636 16830 20638 16882
rect 20638 16830 20690 16882
rect 20690 16830 20692 16882
rect 20636 16828 20692 16830
rect 21868 20130 21924 20132
rect 21868 20078 21870 20130
rect 21870 20078 21922 20130
rect 21922 20078 21924 20130
rect 21868 20076 21924 20078
rect 23436 24722 23492 24724
rect 23436 24670 23438 24722
rect 23438 24670 23490 24722
rect 23490 24670 23492 24722
rect 23436 24668 23492 24670
rect 23100 24444 23156 24500
rect 22876 22876 22932 22932
rect 22988 22258 23044 22260
rect 22988 22206 22990 22258
rect 22990 22206 23042 22258
rect 23042 22206 23044 22258
rect 22988 22204 23044 22206
rect 23212 22092 23268 22148
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 27580 26236 27636 26292
rect 24668 25228 24724 25284
rect 25340 25228 25396 25284
rect 24556 25116 24612 25172
rect 25564 25116 25620 25172
rect 26236 25394 26292 25396
rect 26236 25342 26238 25394
rect 26238 25342 26290 25394
rect 26290 25342 26292 25394
rect 26236 25340 26292 25342
rect 24444 24722 24500 24724
rect 24444 24670 24446 24722
rect 24446 24670 24498 24722
rect 24498 24670 24500 24722
rect 24444 24668 24500 24670
rect 24332 24498 24388 24500
rect 24332 24446 24334 24498
rect 24334 24446 24386 24498
rect 24386 24446 24388 24498
rect 24332 24444 24388 24446
rect 26124 25282 26180 25284
rect 26124 25230 26126 25282
rect 26126 25230 26178 25282
rect 26178 25230 26180 25282
rect 26124 25228 26180 25230
rect 25900 24444 25956 24500
rect 25676 23548 25732 23604
rect 23436 21644 23492 21700
rect 22652 21084 22708 21140
rect 22204 20130 22260 20132
rect 22204 20078 22206 20130
rect 22206 20078 22258 20130
rect 22258 20078 22260 20130
rect 22204 20076 22260 20078
rect 22428 18620 22484 18676
rect 21644 18508 21700 18564
rect 21756 18450 21812 18452
rect 21756 18398 21758 18450
rect 21758 18398 21810 18450
rect 21810 18398 21812 18450
rect 21756 18396 21812 18398
rect 22316 18450 22372 18452
rect 22316 18398 22318 18450
rect 22318 18398 22370 18450
rect 22370 18398 22372 18450
rect 22316 18396 22372 18398
rect 22540 18284 22596 18340
rect 22988 21586 23044 21588
rect 22988 21534 22990 21586
rect 22990 21534 23042 21586
rect 23042 21534 23044 21586
rect 22988 21532 23044 21534
rect 22876 20130 22932 20132
rect 22876 20078 22878 20130
rect 22878 20078 22930 20130
rect 22930 20078 22932 20130
rect 22876 20076 22932 20078
rect 22764 19964 22820 20020
rect 22540 17388 22596 17444
rect 21644 16716 21700 16772
rect 23324 21532 23380 21588
rect 23324 21308 23380 21364
rect 24332 22316 24388 22372
rect 23660 21698 23716 21700
rect 23660 21646 23662 21698
rect 23662 21646 23714 21698
rect 23714 21646 23716 21698
rect 23660 21644 23716 21646
rect 23548 21308 23604 21364
rect 23436 21084 23492 21140
rect 23212 19964 23268 20020
rect 28588 26236 28644 26292
rect 27468 25282 27524 25284
rect 27468 25230 27470 25282
rect 27470 25230 27522 25282
rect 27522 25230 27524 25282
rect 27468 25228 27524 25230
rect 37660 26290 37716 26292
rect 37660 26238 37662 26290
rect 37662 26238 37714 26290
rect 37714 26238 37716 26290
rect 37660 26236 37716 26238
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 40012 25564 40068 25620
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 27132 23436 27188 23492
rect 26348 22204 26404 22260
rect 25564 22092 25620 22148
rect 25228 21810 25284 21812
rect 25228 21758 25230 21810
rect 25230 21758 25282 21810
rect 25282 21758 25284 21810
rect 25228 21756 25284 21758
rect 26908 22482 26964 22484
rect 26908 22430 26910 22482
rect 26910 22430 26962 22482
rect 26962 22430 26964 22482
rect 26908 22428 26964 22430
rect 26908 21980 26964 22036
rect 28252 23042 28308 23044
rect 28252 22990 28254 23042
rect 28254 22990 28306 23042
rect 28306 22990 28308 23042
rect 28252 22988 28308 22990
rect 29260 22988 29316 23044
rect 28028 22540 28084 22596
rect 27244 22370 27300 22372
rect 27244 22318 27246 22370
rect 27246 22318 27298 22370
rect 27298 22318 27300 22370
rect 27244 22316 27300 22318
rect 27580 22370 27636 22372
rect 27580 22318 27582 22370
rect 27582 22318 27634 22370
rect 27634 22318 27636 22370
rect 27580 22316 27636 22318
rect 28476 22316 28532 22372
rect 28700 22316 28756 22372
rect 27804 22146 27860 22148
rect 27804 22094 27806 22146
rect 27806 22094 27858 22146
rect 27858 22094 27860 22146
rect 27804 22092 27860 22094
rect 23996 21532 24052 21588
rect 24668 21586 24724 21588
rect 24668 21534 24670 21586
rect 24670 21534 24722 21586
rect 24722 21534 24724 21586
rect 24668 21532 24724 21534
rect 24332 21420 24388 21476
rect 23996 20130 24052 20132
rect 23996 20078 23998 20130
rect 23998 20078 24050 20130
rect 24050 20078 24052 20130
rect 23996 20076 24052 20078
rect 24108 21308 24164 21364
rect 22988 18396 23044 18452
rect 22876 18284 22932 18340
rect 23212 18172 23268 18228
rect 23100 16994 23156 16996
rect 23100 16942 23102 16994
rect 23102 16942 23154 16994
rect 23154 16942 23156 16994
rect 23100 16940 23156 16942
rect 22764 16604 22820 16660
rect 23772 19852 23828 19908
rect 24108 19794 24164 19796
rect 24108 19742 24110 19794
rect 24110 19742 24162 19794
rect 24162 19742 24164 19794
rect 24108 19740 24164 19742
rect 25900 21586 25956 21588
rect 25900 21534 25902 21586
rect 25902 21534 25954 21586
rect 25954 21534 25956 21586
rect 25900 21532 25956 21534
rect 26012 21420 26068 21476
rect 30044 22316 30100 22372
rect 29148 22258 29204 22260
rect 29148 22206 29150 22258
rect 29150 22206 29202 22258
rect 29202 22206 29204 22258
rect 29148 22204 29204 22206
rect 29372 22146 29428 22148
rect 29372 22094 29374 22146
rect 29374 22094 29426 22146
rect 29426 22094 29428 22146
rect 29372 22092 29428 22094
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 37660 22540 37716 22596
rect 37660 22370 37716 22372
rect 37660 22318 37662 22370
rect 37662 22318 37714 22370
rect 37714 22318 37716 22370
rect 37660 22316 37716 22318
rect 40012 22204 40068 22260
rect 30380 21532 30436 21588
rect 25900 19740 25956 19796
rect 25676 19180 25732 19236
rect 27916 19234 27972 19236
rect 27916 19182 27918 19234
rect 27918 19182 27970 19234
rect 27970 19182 27972 19234
rect 27916 19180 27972 19182
rect 29260 20690 29316 20692
rect 29260 20638 29262 20690
rect 29262 20638 29314 20690
rect 29314 20638 29316 20690
rect 29260 20636 29316 20638
rect 37660 21586 37716 21588
rect 37660 21534 37662 21586
rect 37662 21534 37714 21586
rect 37714 21534 37716 21586
rect 37660 21532 37716 21534
rect 40012 21532 40068 21588
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 30380 20636 30436 20692
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 37660 19234 37716 19236
rect 37660 19182 37662 19234
rect 37662 19182 37714 19234
rect 37714 19182 37716 19234
rect 37660 19180 37716 19182
rect 29036 19068 29092 19124
rect 25900 18956 25956 19012
rect 27356 18956 27412 19012
rect 23548 18396 23604 18452
rect 25452 18450 25508 18452
rect 25452 18398 25454 18450
rect 25454 18398 25506 18450
rect 25506 18398 25508 18450
rect 25452 18396 25508 18398
rect 25228 18226 25284 18228
rect 25228 18174 25230 18226
rect 25230 18174 25282 18226
rect 25282 18174 25284 18226
rect 25228 18172 25284 18174
rect 23436 17612 23492 17668
rect 23996 17612 24052 17668
rect 23548 16716 23604 16772
rect 23436 16604 23492 16660
rect 21644 15820 21700 15876
rect 21644 15148 21700 15204
rect 19292 15036 19348 15092
rect 22316 15036 22372 15092
rect 20748 14530 20804 14532
rect 20748 14478 20750 14530
rect 20750 14478 20802 14530
rect 20802 14478 20804 14530
rect 20748 14476 20804 14478
rect 21420 14476 21476 14532
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19292 13468 19348 13524
rect 19292 13074 19348 13076
rect 19292 13022 19294 13074
rect 19294 13022 19346 13074
rect 19346 13022 19348 13074
rect 19292 13020 19348 13022
rect 21756 13468 21812 13524
rect 21532 13020 21588 13076
rect 22876 15036 22932 15092
rect 22428 13020 22484 13076
rect 23548 15372 23604 15428
rect 26348 17554 26404 17556
rect 26348 17502 26350 17554
rect 26350 17502 26402 17554
rect 26402 17502 26404 17554
rect 26348 17500 26404 17502
rect 27692 19010 27748 19012
rect 27692 18958 27694 19010
rect 27694 18958 27746 19010
rect 27746 18958 27748 19010
rect 27692 18956 27748 18958
rect 28140 19010 28196 19012
rect 28140 18958 28142 19010
rect 28142 18958 28194 19010
rect 28194 18958 28196 19010
rect 28140 18956 28196 18958
rect 26908 17500 26964 17556
rect 25004 15372 25060 15428
rect 23100 15314 23156 15316
rect 23100 15262 23102 15314
rect 23102 15262 23154 15314
rect 23154 15262 23156 15314
rect 23100 15260 23156 15262
rect 23212 15202 23268 15204
rect 23212 15150 23214 15202
rect 23214 15150 23266 15202
rect 23266 15150 23268 15202
rect 23212 15148 23268 15150
rect 24108 15202 24164 15204
rect 24108 15150 24110 15202
rect 24110 15150 24162 15202
rect 24162 15150 24164 15202
rect 24108 15148 24164 15150
rect 29260 19122 29316 19124
rect 29260 19070 29262 19122
rect 29262 19070 29314 19122
rect 29314 19070 29316 19122
rect 29260 19068 29316 19070
rect 30156 19068 30212 19124
rect 29484 19010 29540 19012
rect 29484 18958 29486 19010
rect 29486 18958 29538 19010
rect 29538 18958 29540 19010
rect 29484 18956 29540 18958
rect 29260 17554 29316 17556
rect 29260 17502 29262 17554
rect 29262 17502 29314 17554
rect 29314 17502 29316 17554
rect 29260 17500 29316 17502
rect 29932 17500 29988 17556
rect 28028 17388 28084 17444
rect 29484 17442 29540 17444
rect 29484 17390 29486 17442
rect 29486 17390 29538 17442
rect 29538 17390 29540 17442
rect 29484 17388 29540 17390
rect 40012 18844 40068 18900
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 37660 17666 37716 17668
rect 37660 17614 37662 17666
rect 37662 17614 37714 17666
rect 37714 17614 37716 17666
rect 37660 17612 37716 17614
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 37884 17500 37940 17556
rect 40012 17500 40068 17556
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 27580 15372 27636 15428
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 24668 13634 24724 13636
rect 24668 13582 24670 13634
rect 24670 13582 24722 13634
rect 24722 13582 24724 13634
rect 24668 13580 24724 13582
rect 25788 13580 25844 13636
rect 25004 13468 25060 13524
rect 24444 13074 24500 13076
rect 24444 13022 24446 13074
rect 24446 13022 24498 13074
rect 24498 13022 24500 13074
rect 24444 13020 24500 13022
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 18844 4060 18900 4116
rect 16828 3388 16884 3444
rect 18060 3388 18116 3444
rect 20076 4114 20132 4116
rect 20076 4062 20078 4114
rect 20078 4062 20130 4114
rect 20130 4062 20132 4114
rect 20076 4060 20132 4062
rect 24220 4060 24276 4116
rect 23548 3612 23604 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 26236 4114 26292 4116
rect 26236 4062 26238 4114
rect 26238 4062 26290 4114
rect 26290 4062 26292 4114
rect 26236 4060 26292 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
<< metal3 >>
rect 25554 38556 25564 38612
rect 25620 38556 26796 38612
rect 26852 38556 26862 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 20850 38220 20860 38276
rect 20916 38220 22092 38276
rect 22148 38220 22158 38276
rect 24210 38220 24220 38276
rect 24276 38220 25564 38276
rect 25620 38220 25630 38276
rect 18050 37996 18060 38052
rect 18116 37996 18732 38052
rect 18788 37996 18798 38052
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 16146 37436 16156 37492
rect 16212 37436 18396 37492
rect 18452 37436 18462 37492
rect 20178 37436 20188 37492
rect 20244 37436 21420 37492
rect 21476 37436 21486 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 15474 36652 15484 36708
rect 15540 36652 16716 36708
rect 16772 36652 16782 36708
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 16146 28028 16156 28084
rect 16212 28028 16604 28084
rect 16660 28028 17388 28084
rect 17444 28028 17454 28084
rect 0 27636 800 27664
rect 0 27580 4172 27636
rect 4228 27580 4238 27636
rect 0 27552 800 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 14914 27020 14924 27076
rect 14980 27020 15484 27076
rect 15540 27020 16604 27076
rect 16660 27020 16670 27076
rect 23314 27020 23324 27076
rect 23380 27020 24220 27076
rect 24276 27020 24556 27076
rect 24612 27020 24622 27076
rect 20178 26684 20188 26740
rect 20244 26684 20636 26740
rect 20692 26684 20702 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 13906 26460 13916 26516
rect 13972 26460 16380 26516
rect 16436 26460 16446 26516
rect 18162 26460 18172 26516
rect 18228 26460 18956 26516
rect 19012 26460 19022 26516
rect 15138 26348 15148 26404
rect 15204 26348 16044 26404
rect 16100 26348 16110 26404
rect 19058 26236 19068 26292
rect 19124 26236 20860 26292
rect 20916 26236 20926 26292
rect 27570 26236 27580 26292
rect 27636 26236 28588 26292
rect 28644 26236 37660 26292
rect 37716 26236 37726 26292
rect 18498 26124 18508 26180
rect 18564 26124 20412 26180
rect 20468 26124 20478 26180
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 41200 25620 42000 25648
rect 40002 25564 40012 25620
rect 40068 25564 42000 25620
rect 41200 25536 42000 25564
rect 18834 25452 18844 25508
rect 18900 25452 20076 25508
rect 20132 25452 21420 25508
rect 21476 25452 21486 25508
rect 16146 25340 16156 25396
rect 16212 25340 17500 25396
rect 17556 25340 20188 25396
rect 20244 25340 20254 25396
rect 20402 25340 20412 25396
rect 20468 25340 26236 25396
rect 26292 25340 26302 25396
rect 13234 25228 13244 25284
rect 13300 25228 14028 25284
rect 14084 25228 15036 25284
rect 15092 25228 15820 25284
rect 15876 25228 16828 25284
rect 16884 25228 19180 25284
rect 19236 25228 21308 25284
rect 21364 25228 22652 25284
rect 22708 25228 23548 25284
rect 23604 25228 24668 25284
rect 24724 25228 25340 25284
rect 25396 25228 25406 25284
rect 26114 25228 26124 25284
rect 26180 25228 27468 25284
rect 27524 25228 27534 25284
rect 20514 25116 20524 25172
rect 20580 25116 21756 25172
rect 21812 25116 21822 25172
rect 24546 25116 24556 25172
rect 24612 25116 25564 25172
rect 25620 25116 25630 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 0 24948 800 24976
rect 0 24892 1932 24948
rect 1988 24892 1998 24948
rect 16594 24892 16604 24948
rect 16660 24892 17612 24948
rect 17668 24892 17678 24948
rect 18498 24892 18508 24948
rect 18564 24892 19404 24948
rect 19460 24892 19470 24948
rect 0 24864 800 24892
rect 18508 24836 18564 24892
rect 17378 24780 17388 24836
rect 17444 24780 18564 24836
rect 23426 24668 23436 24724
rect 23492 24668 24444 24724
rect 24500 24668 24510 24724
rect 4274 24556 4284 24612
rect 4340 24556 11116 24612
rect 11172 24556 14588 24612
rect 14644 24556 14654 24612
rect 17714 24556 17724 24612
rect 17780 24556 18732 24612
rect 18788 24556 18798 24612
rect 22418 24444 22428 24500
rect 22484 24444 23100 24500
rect 23156 24444 24332 24500
rect 24388 24444 25900 24500
rect 25956 24444 25966 24500
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 13234 23996 13244 24052
rect 13300 23996 14476 24052
rect 14532 23996 14542 24052
rect 14354 23884 14364 23940
rect 14420 23884 14812 23940
rect 14868 23884 17388 23940
rect 17444 23884 17454 23940
rect 18834 23884 18844 23940
rect 18900 23884 19516 23940
rect 19572 23884 20076 23940
rect 20132 23884 20142 23940
rect 18722 23772 18732 23828
rect 18788 23772 19740 23828
rect 19796 23772 19806 23828
rect 14690 23548 14700 23604
rect 14756 23548 14766 23604
rect 25666 23548 25676 23604
rect 25732 23548 26908 23604
rect 14700 23492 14756 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 26852 23492 26908 23548
rect 14700 23436 16492 23492
rect 16548 23436 16558 23492
rect 26852 23436 27132 23492
rect 27188 23436 27198 23492
rect 14924 23324 21532 23380
rect 21588 23324 22540 23380
rect 22596 23324 22606 23380
rect 14924 23156 14980 23324
rect 4274 23100 4284 23156
rect 4340 23100 9996 23156
rect 10052 23100 10062 23156
rect 14914 23100 14924 23156
rect 14980 23100 14990 23156
rect 12898 22988 12908 23044
rect 12964 22988 14028 23044
rect 14084 22988 15820 23044
rect 15876 22988 15886 23044
rect 19058 22988 19068 23044
rect 19124 22988 20300 23044
rect 20356 22988 20366 23044
rect 28242 22988 28252 23044
rect 28308 22988 29260 23044
rect 29316 22988 29326 23044
rect 0 22932 800 22960
rect 41200 22932 42000 22960
rect 0 22876 1932 22932
rect 1988 22876 1998 22932
rect 14690 22876 14700 22932
rect 14756 22876 15372 22932
rect 15428 22876 20412 22932
rect 20468 22876 22876 22932
rect 22932 22876 22942 22932
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 0 22848 800 22876
rect 41200 22848 42000 22876
rect 19282 22764 19292 22820
rect 19348 22764 19740 22820
rect 19796 22764 21868 22820
rect 21924 22764 21934 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 8372 22652 11228 22708
rect 11284 22652 15484 22708
rect 15540 22652 15550 22708
rect 1922 22428 1932 22484
rect 1988 22428 1998 22484
rect 0 22260 800 22288
rect 1932 22260 1988 22428
rect 8372 22372 8428 22652
rect 12114 22540 12124 22596
rect 12180 22540 15260 22596
rect 15316 22540 15326 22596
rect 15698 22540 15708 22596
rect 15764 22540 17724 22596
rect 17780 22540 28028 22596
rect 28084 22540 28094 22596
rect 31892 22540 37660 22596
rect 37716 22540 37726 22596
rect 15708 22484 15764 22540
rect 31892 22484 31948 22540
rect 13346 22428 13356 22484
rect 13412 22428 14476 22484
rect 14532 22428 14542 22484
rect 14924 22428 15764 22484
rect 26898 22428 26908 22484
rect 26964 22428 31948 22484
rect 14924 22372 14980 22428
rect 4274 22316 4284 22372
rect 4340 22316 8428 22372
rect 14018 22316 14028 22372
rect 14084 22316 14980 22372
rect 15138 22316 15148 22372
rect 15204 22316 15820 22372
rect 15876 22316 15886 22372
rect 24322 22316 24332 22372
rect 24388 22316 27244 22372
rect 27300 22316 27310 22372
rect 27570 22316 27580 22372
rect 27636 22316 28476 22372
rect 28532 22316 28542 22372
rect 28690 22316 28700 22372
rect 28756 22316 30044 22372
rect 30100 22316 37660 22372
rect 37716 22316 37726 22372
rect 41200 22260 42000 22288
rect 0 22204 1988 22260
rect 9986 22204 9996 22260
rect 10052 22204 13916 22260
rect 13972 22204 13982 22260
rect 17378 22204 17388 22260
rect 17444 22204 19516 22260
rect 19572 22204 19582 22260
rect 22306 22204 22316 22260
rect 22372 22204 22988 22260
rect 23044 22204 23054 22260
rect 26338 22204 26348 22260
rect 26404 22204 29148 22260
rect 29204 22204 29214 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 0 22176 800 22204
rect 41200 22176 42000 22204
rect 19730 22092 19740 22148
rect 19796 22092 20524 22148
rect 20580 22092 20972 22148
rect 21028 22092 23212 22148
rect 23268 22092 23278 22148
rect 25554 22092 25564 22148
rect 25620 22092 27804 22148
rect 27860 22092 29372 22148
rect 29428 22092 29438 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 14802 21868 14812 21924
rect 14868 21868 14878 21924
rect 15698 21868 15708 21924
rect 15764 21868 16716 21924
rect 16772 21868 16782 21924
rect 20178 21868 20188 21924
rect 20244 21868 21644 21924
rect 21700 21868 22316 21924
rect 22372 21868 22382 21924
rect 4274 21532 4284 21588
rect 4340 21532 9884 21588
rect 9940 21532 9950 21588
rect 14812 21364 14868 21868
rect 23212 21812 23268 22092
rect 26898 21980 26908 22036
rect 26964 21980 26974 22036
rect 26908 21812 26964 21980
rect 19170 21756 19180 21812
rect 19236 21756 19246 21812
rect 23212 21756 25228 21812
rect 25284 21756 25294 21812
rect 26852 21756 26964 21812
rect 15250 21532 15260 21588
rect 15316 21532 16044 21588
rect 16100 21532 16110 21588
rect 19180 21476 19236 21756
rect 26852 21700 26908 21756
rect 19394 21644 19404 21700
rect 19460 21644 23436 21700
rect 23492 21644 23502 21700
rect 23650 21644 23660 21700
rect 23716 21644 26908 21700
rect 41200 21588 42000 21616
rect 22082 21532 22092 21588
rect 22148 21532 22988 21588
rect 23044 21532 23054 21588
rect 23314 21532 23324 21588
rect 23380 21532 23996 21588
rect 24052 21532 24668 21588
rect 24724 21532 25900 21588
rect 25956 21532 25966 21588
rect 30370 21532 30380 21588
rect 30436 21532 37660 21588
rect 37716 21532 37726 21588
rect 40002 21532 40012 21588
rect 40068 21532 42000 21588
rect 41200 21504 42000 21532
rect 19180 21420 24332 21476
rect 24388 21420 26012 21476
rect 26068 21420 26078 21476
rect 23324 21364 23380 21420
rect 13234 21308 13244 21364
rect 13300 21308 15708 21364
rect 15764 21308 15774 21364
rect 19730 21308 19740 21364
rect 19796 21308 20524 21364
rect 20580 21308 20590 21364
rect 23314 21308 23324 21364
rect 23380 21308 23390 21364
rect 23538 21308 23548 21364
rect 23604 21308 24108 21364
rect 24164 21308 24174 21364
rect 23548 21252 23604 21308
rect 15810 21196 15820 21252
rect 15876 21196 16156 21252
rect 16212 21196 19852 21252
rect 19908 21196 19918 21252
rect 20076 21196 23604 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 20076 21140 20132 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 15026 21084 15036 21140
rect 15092 21084 16940 21140
rect 16996 21084 18620 21140
rect 18676 21084 20132 21140
rect 22642 21084 22652 21140
rect 22708 21084 23436 21140
rect 23492 21084 23502 21140
rect 4162 20972 4172 21028
rect 4228 20972 8428 21028
rect 15586 20972 15596 21028
rect 15652 20972 16492 21028
rect 16548 20972 18956 21028
rect 19012 20972 19022 21028
rect 0 20916 800 20944
rect 0 20860 1932 20916
rect 1988 20860 1998 20916
rect 0 20832 800 20860
rect 8372 20804 8428 20972
rect 18162 20860 18172 20916
rect 18228 20860 19180 20916
rect 19236 20860 19246 20916
rect 8372 20748 21308 20804
rect 21364 20748 21374 20804
rect 9874 20636 9884 20692
rect 9940 20636 13468 20692
rect 13524 20636 13534 20692
rect 20402 20636 20412 20692
rect 20468 20636 20972 20692
rect 21028 20636 21038 20692
rect 29250 20636 29260 20692
rect 29316 20636 30380 20692
rect 30436 20636 30446 20692
rect 14578 20524 14588 20580
rect 14644 20524 15708 20580
rect 15764 20524 15774 20580
rect 20626 20524 20636 20580
rect 20692 20524 21420 20580
rect 21476 20524 21486 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 12002 20188 12012 20244
rect 12068 20188 14476 20244
rect 14532 20188 14542 20244
rect 16818 20076 16828 20132
rect 16884 20076 17612 20132
rect 17668 20076 17678 20132
rect 20290 20076 20300 20132
rect 20356 20076 21532 20132
rect 21588 20076 21868 20132
rect 21924 20076 21934 20132
rect 22194 20076 22204 20132
rect 22260 20076 22270 20132
rect 22866 20076 22876 20132
rect 22932 20076 23996 20132
rect 24052 20076 24062 20132
rect 22204 20020 22260 20076
rect 16146 19964 16156 20020
rect 16212 19964 18060 20020
rect 18116 19964 18126 20020
rect 18610 19964 18620 20020
rect 18676 19964 19068 20020
rect 19124 19964 19852 20020
rect 19908 19964 19918 20020
rect 22204 19964 22764 20020
rect 22820 19964 23212 20020
rect 23268 19964 23278 20020
rect 12114 19852 12124 19908
rect 12180 19852 13356 19908
rect 13412 19852 13422 19908
rect 16034 19852 16044 19908
rect 16100 19852 18732 19908
rect 18788 19852 23772 19908
rect 23828 19852 23838 19908
rect 24098 19740 24108 19796
rect 24164 19740 25900 19796
rect 25956 19740 25966 19796
rect 13794 19628 13804 19684
rect 13860 19628 15932 19684
rect 15988 19628 18508 19684
rect 18564 19628 18574 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 4274 19180 4284 19236
rect 4340 19180 9996 19236
rect 10052 19180 13132 19236
rect 13188 19180 13804 19236
rect 13860 19180 13870 19236
rect 25666 19180 25676 19236
rect 25732 19180 27916 19236
rect 27972 19180 27982 19236
rect 31892 19180 37660 19236
rect 37716 19180 37726 19236
rect 31892 19124 31948 19180
rect 16482 19068 16492 19124
rect 16548 19068 29036 19124
rect 29092 19068 29102 19124
rect 29250 19068 29260 19124
rect 29316 19068 30156 19124
rect 30212 19068 31948 19124
rect 12898 18956 12908 19012
rect 12964 18956 14364 19012
rect 14420 18956 14430 19012
rect 15092 18956 15484 19012
rect 15540 18956 15550 19012
rect 15698 18956 15708 19012
rect 15764 18956 17164 19012
rect 17220 18956 18172 19012
rect 18228 18956 18238 19012
rect 25890 18956 25900 19012
rect 25956 18956 27356 19012
rect 27412 18956 27692 19012
rect 27748 18956 27758 19012
rect 28130 18956 28140 19012
rect 28196 18956 29484 19012
rect 29540 18956 29550 19012
rect 0 18900 800 18928
rect 0 18844 1932 18900
rect 1988 18844 1998 18900
rect 0 18816 800 18844
rect 15092 18788 15148 18956
rect 41200 18900 42000 18928
rect 40002 18844 40012 18900
rect 40068 18844 42000 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 41200 18816 42000 18844
rect 13906 18732 13916 18788
rect 13972 18732 14476 18788
rect 14532 18732 15148 18788
rect 15204 18732 15214 18788
rect 19842 18620 19852 18676
rect 19908 18620 22428 18676
rect 22484 18620 22494 18676
rect 19506 18508 19516 18564
rect 19572 18508 21644 18564
rect 21700 18508 21710 18564
rect 4274 18396 4284 18452
rect 4340 18396 12908 18452
rect 12964 18396 12974 18452
rect 17938 18396 17948 18452
rect 18004 18396 18620 18452
rect 18676 18396 18956 18452
rect 19012 18396 19628 18452
rect 19684 18396 19694 18452
rect 21746 18396 21756 18452
rect 21812 18396 22316 18452
rect 22372 18396 22988 18452
rect 23044 18396 23054 18452
rect 23538 18396 23548 18452
rect 23604 18396 25452 18452
rect 25508 18396 25518 18452
rect 16818 18284 16828 18340
rect 16884 18284 19180 18340
rect 19236 18284 20636 18340
rect 20692 18284 20702 18340
rect 22530 18284 22540 18340
rect 22596 18284 22876 18340
rect 22932 18284 22942 18340
rect 0 18228 800 18256
rect 41200 18228 42000 18256
rect 0 18172 1932 18228
rect 1988 18172 1998 18228
rect 18274 18172 18284 18228
rect 18340 18172 21420 18228
rect 21476 18172 21486 18228
rect 23202 18172 23212 18228
rect 23268 18172 25228 18228
rect 25284 18172 25294 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 0 18144 800 18172
rect 41200 18144 42000 18172
rect 18498 18060 18508 18116
rect 18564 18060 19964 18116
rect 20020 18060 20030 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 17490 17724 17500 17780
rect 17556 17724 18508 17780
rect 18564 17724 18574 17780
rect 23426 17612 23436 17668
rect 23492 17612 23996 17668
rect 24052 17612 37660 17668
rect 37716 17612 37726 17668
rect 41200 17556 42000 17584
rect 26338 17500 26348 17556
rect 26404 17500 26908 17556
rect 26964 17500 26974 17556
rect 29250 17500 29260 17556
rect 29316 17500 29932 17556
rect 29988 17500 37884 17556
rect 37940 17500 37950 17556
rect 40002 17500 40012 17556
rect 40068 17500 42000 17556
rect 41200 17472 42000 17500
rect 16706 17388 16716 17444
rect 16772 17388 17836 17444
rect 17892 17388 18620 17444
rect 18676 17388 19516 17444
rect 19572 17388 19852 17444
rect 19908 17388 19918 17444
rect 20514 17388 20524 17444
rect 20580 17388 22540 17444
rect 22596 17388 22606 17444
rect 28018 17388 28028 17444
rect 28084 17388 29484 17444
rect 29540 17388 29550 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 16594 16940 16604 16996
rect 16660 16940 17612 16996
rect 17668 16940 18172 16996
rect 18228 16940 23100 16996
rect 23156 16940 23166 16996
rect 17826 16828 17836 16884
rect 17892 16828 19180 16884
rect 19236 16828 20636 16884
rect 20692 16828 20702 16884
rect 15474 16716 15484 16772
rect 15540 16716 16492 16772
rect 16548 16716 16558 16772
rect 18946 16716 18956 16772
rect 19012 16716 20412 16772
rect 20468 16716 20478 16772
rect 21634 16716 21644 16772
rect 21700 16716 23548 16772
rect 23604 16716 23614 16772
rect 15250 16604 15260 16660
rect 15316 16604 16380 16660
rect 16436 16604 20300 16660
rect 20356 16604 20366 16660
rect 22754 16604 22764 16660
rect 22820 16604 23436 16660
rect 23492 16604 23502 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 20178 15820 20188 15876
rect 20244 15820 21644 15876
rect 21700 15820 21710 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 23538 15372 23548 15428
rect 23604 15372 25004 15428
rect 25060 15372 27580 15428
rect 27636 15372 27646 15428
rect 16482 15260 16492 15316
rect 16548 15260 16940 15316
rect 16996 15260 17006 15316
rect 17378 15260 17388 15316
rect 17444 15260 18284 15316
rect 18340 15260 23100 15316
rect 23156 15260 23166 15316
rect 17388 15204 17444 15260
rect 16828 15148 17444 15204
rect 21634 15148 21644 15204
rect 21700 15148 22932 15204
rect 23202 15148 23212 15204
rect 23268 15148 24108 15204
rect 24164 15148 24174 15204
rect 16828 15092 16884 15148
rect 22876 15092 22932 15148
rect 16818 15036 16828 15092
rect 16884 15036 16894 15092
rect 18834 15036 18844 15092
rect 18900 15036 19292 15092
rect 19348 15036 22316 15092
rect 22372 15036 22382 15092
rect 22866 15036 22876 15092
rect 22932 15036 22942 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 15586 14476 15596 14532
rect 15652 14476 16940 14532
rect 16996 14476 17006 14532
rect 20738 14476 20748 14532
rect 20804 14476 21420 14532
rect 21476 14476 21486 14532
rect 14690 14364 14700 14420
rect 14756 14364 15484 14420
rect 15540 14364 15550 14420
rect 17154 14364 17164 14420
rect 17220 14364 18396 14420
rect 18452 14364 18462 14420
rect 16594 14252 16604 14308
rect 16660 14252 17052 14308
rect 17108 14252 17118 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 24658 13580 24668 13636
rect 24724 13580 25788 13636
rect 25844 13580 25854 13636
rect 14018 13468 14028 13524
rect 14084 13468 15932 13524
rect 15988 13468 16716 13524
rect 16772 13468 17500 13524
rect 17556 13468 19292 13524
rect 19348 13468 19358 13524
rect 21746 13468 21756 13524
rect 21812 13468 25004 13524
rect 25060 13468 25070 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19282 13020 19292 13076
rect 19348 13020 21532 13076
rect 21588 13020 21598 13076
rect 22418 13020 22428 13076
rect 22484 13020 24444 13076
rect 24500 13020 24510 13076
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 18834 4060 18844 4116
rect 18900 4060 20076 4116
rect 20132 4060 20142 4116
rect 24210 4060 24220 4116
rect 24276 4060 26236 4116
rect 26292 4060 26302 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 23538 3612 23548 3668
rect 23604 3612 25564 3668
rect 25620 3612 25630 3668
rect 16818 3388 16828 3444
rect 16884 3388 18060 3444
rect 18116 3388 18126 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17696 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21056 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1698175906
transform -1 0 20832 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16240 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19376 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_
timestamp 1698175906
transform -1 0 20944 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18816 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18816 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _111_
timestamp 1698175906
transform -1 0 17696 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1698175906
transform -1 0 17920 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _113_
timestamp 1698175906
transform -1 0 17024 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16240 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _115_
timestamp 1698175906
transform -1 0 19376 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _116_
timestamp 1698175906
transform -1 0 18816 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform -1 0 16352 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698175906
transform -1 0 21840 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _119_
timestamp 1698175906
transform 1 0 17920 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19936 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17808 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _122_
timestamp 1698175906
transform -1 0 18144 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698175906
transform -1 0 17920 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14672 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _125_
timestamp 1698175906
transform 1 0 15904 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform -1 0 20944 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _127_
timestamp 1698175906
transform 1 0 18816 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _128_
timestamp 1698175906
transform 1 0 19152 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_
timestamp 1698175906
transform -1 0 20048 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19264 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _131_
timestamp 1698175906
transform -1 0 17920 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _132_
timestamp 1698175906
transform -1 0 16016 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _133_
timestamp 1698175906
transform -1 0 14112 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _134_
timestamp 1698175906
transform 1 0 21280 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _135_
timestamp 1698175906
transform 1 0 18928 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _136_
timestamp 1698175906
transform 1 0 19600 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _137_
timestamp 1698175906
transform -1 0 16016 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13104 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _139_
timestamp 1698175906
transform 1 0 21728 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _140_
timestamp 1698175906
transform -1 0 15680 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _141_
timestamp 1698175906
transform 1 0 14784 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _142_
timestamp 1698175906
transform 1 0 21168 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _143_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21056 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _144_
timestamp 1698175906
transform 1 0 22064 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _145_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19824 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _146_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18928 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _147_
timestamp 1698175906
transform 1 0 17808 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _148_
timestamp 1698175906
transform -1 0 15456 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _149_
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _150_
timestamp 1698175906
transform -1 0 17024 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _151_
timestamp 1698175906
transform 1 0 15456 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _152_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14000 0 -1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _153_
timestamp 1698175906
transform -1 0 20944 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _154_
timestamp 1698175906
transform 1 0 19488 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _155_
timestamp 1698175906
transform -1 0 22064 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _156_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18032 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _157_
timestamp 1698175906
transform 1 0 15344 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _158_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14224 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _159_
timestamp 1698175906
transform -1 0 21168 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _160_
timestamp 1698175906
transform 1 0 19712 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _161_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22064 0 -1 21952
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _162_
timestamp 1698175906
transform 1 0 20048 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _163_
timestamp 1698175906
transform 1 0 18928 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _164_
timestamp 1698175906
transform 1 0 19376 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _165_
timestamp 1698175906
transform 1 0 18704 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _166_
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _167_
timestamp 1698175906
transform 1 0 22400 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _168_
timestamp 1698175906
transform 1 0 23856 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _169_
timestamp 1698175906
transform -1 0 23744 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _170_
timestamp 1698175906
transform 1 0 22848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _171_
timestamp 1698175906
transform 1 0 22960 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _172_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _173_
timestamp 1698175906
transform 1 0 23856 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _174_
timestamp 1698175906
transform -1 0 23856 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _175_
timestamp 1698175906
transform 1 0 22624 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _176_
timestamp 1698175906
transform 1 0 24304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform -1 0 14224 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _178_
timestamp 1698175906
transform 1 0 14336 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _179_
timestamp 1698175906
transform 1 0 28224 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _180_
timestamp 1698175906
transform 1 0 23968 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _181_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 28224 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _182_
timestamp 1698175906
transform -1 0 14784 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _183_
timestamp 1698175906
transform 1 0 14000 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _184_
timestamp 1698175906
transform 1 0 25760 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _185_
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _186_
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _187_
timestamp 1698175906
transform 1 0 18144 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _188_
timestamp 1698175906
transform -1 0 17360 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _189_
timestamp 1698175906
transform -1 0 22848 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _190_
timestamp 1698175906
transform 1 0 22848 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _191_
timestamp 1698175906
transform 1 0 21280 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _192_
timestamp 1698175906
transform -1 0 27776 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _193_
timestamp 1698175906
transform 1 0 19936 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _194_
timestamp 1698175906
transform 1 0 25760 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _195_
timestamp 1698175906
transform 1 0 24192 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _196_
timestamp 1698175906
transform 1 0 22512 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _197_
timestamp 1698175906
transform -1 0 23856 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _198_
timestamp 1698175906
transform 1 0 22176 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _199_
timestamp 1698175906
transform 1 0 22736 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _200_
timestamp 1698175906
transform 1 0 19600 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _201_
timestamp 1698175906
transform 1 0 20160 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _202_
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _203_
timestamp 1698175906
transform 1 0 27552 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _204_
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _205_
timestamp 1698175906
transform 1 0 27216 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13776 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _207_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12992 0 -1 28224
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform 1 0 15680 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform -1 0 13104 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform -1 0 25984 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 13776 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform -1 0 20944 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform -1 0 12992 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform -1 0 14336 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 17248 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform -1 0 27104 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 21616 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 23856 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform -1 0 13104 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 26992 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform -1 0 14224 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 27328 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 15680 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 21168 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 25536 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform 1 0 22512 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 21392 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 17584 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 27104 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 26880 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _233_
timestamp 1698175906
transform -1 0 16912 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _234_
timestamp 1698175906
transform -1 0 13440 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _235_
timestamp 1698175906
transform 1 0 15232 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17472 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform -1 0 16912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 19152 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 14336 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 26208 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 17024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 16800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 21392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform -1 0 14224 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 15792 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 27328 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 26768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 13104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform -1 0 27216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 15008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 27104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform -1 0 19376 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 25760 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform -1 0 25088 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform -1 0 21280 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 26880 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 26656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 21168 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_165 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698175906
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_312 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 36288 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_328 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 38080 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_336
timestamp 1698175906
transform 1 0 38976 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698175906
transform 1 0 18144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_154
timestamp 1698175906
transform 1 0 18592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_156
timestamp 1698175906
transform 1 0 18816 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_183
timestamp 1698175906
transform 1 0 21840 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_199
timestamp 1698175906
transform 1 0 23632 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 28000 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 31584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_123
timestamp 1698175906
transform 1 0 15120 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_127
timestamp 1698175906
transform 1 0 15568 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_157
timestamp 1698175906
transform 1 0 18928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_161
timestamp 1698175906
transform 1 0 19376 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_169
timestamp 1698175906
transform 1 0 20272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698175906
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_208
timestamp 1698175906
transform 1 0 24640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_212
timestamp 1698175906
transform 1 0 25088 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698175906
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_104
timestamp 1698175906
transform 1 0 12992 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_108
timestamp 1698175906
transform 1 0 13440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_110
timestamp 1698175906
transform 1 0 13664 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_146
timestamp 1698175906
transform 1 0 17696 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_158
timestamp 1698175906
transform 1 0 19040 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_174
timestamp 1698175906
transform 1 0 20832 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_178
timestamp 1698175906
transform 1 0 21280 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_180
timestamp 1698175906
transform 1 0 21504 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_216
timestamp 1698175906
transform 1 0 25536 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_133
timestamp 1698175906
transform 1 0 16240 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_143
timestamp 1698175906
transform 1 0 17360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_145
timestamp 1698175906
transform 1 0 17584 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_181
timestamp 1698175906
transform 1 0 21616 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_185
timestamp 1698175906
transform 1 0 22064 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_220
timestamp 1698175906
transform 1 0 25984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_224
timestamp 1698175906
transform 1 0 26432 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_240
timestamp 1698175906
transform 1 0 28224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_104
timestamp 1698175906
transform 1 0 12992 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_120
timestamp 1698175906
transform 1 0 14784 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_128
timestamp 1698175906
transform 1 0 15680 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_132
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_148
timestamp 1698175906
transform 1 0 17920 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_180
timestamp 1698175906
transform 1 0 21504 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_188
timestamp 1698175906
transform 1 0 22400 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_190
timestamp 1698175906
transform 1 0 22624 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698175906
transform 1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_136
timestamp 1698175906
transform 1 0 16576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_140
timestamp 1698175906
transform 1 0 17024 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_156
timestamp 1698175906
transform 1 0 18816 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_164
timestamp 1698175906
transform 1 0 19712 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698175906
transform 1 0 20720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_185
timestamp 1698175906
transform 1 0 22064 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_189
timestamp 1698175906
transform 1 0 22512 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_199
timestamp 1698175906
transform 1 0 23632 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_230
timestamp 1698175906
transform 1 0 27104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_234
timestamp 1698175906
transform 1 0 27552 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698175906
transform 1 0 28448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_104
timestamp 1698175906
transform 1 0 12992 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_128
timestamp 1698175906
transform 1 0 15680 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_132
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_150
timestamp 1698175906
transform 1 0 18144 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_154
timestamp 1698175906
transform 1 0 18592 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_156
timestamp 1698175906
transform 1 0 18816 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_175
timestamp 1698175906
transform 1 0 20944 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_183
timestamp 1698175906
transform 1 0 21840 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_191
timestamp 1698175906
transform 1 0 22736 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_201
timestamp 1698175906
transform 1 0 23856 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_259
timestamp 1698175906
transform 1 0 30352 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_275
timestamp 1698175906
transform 1 0 32144 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_115
timestamp 1698175906
transform 1 0 14224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_119
timestamp 1698175906
transform 1 0 14672 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_121
timestamp 1698175906
transform 1 0 14896 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_128
timestamp 1698175906
transform 1 0 15680 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_136
timestamp 1698175906
transform 1 0 16576 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_227
timestamp 1698175906
transform 1 0 26768 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_239
timestamp 1698175906
transform 1 0 28112 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698175906
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_252
timestamp 1698175906
transform 1 0 29568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_284
timestamp 1698175906
transform 1 0 33152 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_300
timestamp 1698175906
transform 1 0 34944 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_308
timestamp 1698175906
transform 1 0 35840 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_312
timestamp 1698175906
transform 1 0 36288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698175906
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 4480 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 8064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_88
timestamp 1698175906
transform 1 0 11200 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_96
timestamp 1698175906
transform 1 0 12096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_100
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_108
timestamp 1698175906
transform 1 0 13440 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_110
timestamp 1698175906
transform 1 0 13664 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_183
timestamp 1698175906
transform 1 0 21840 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_191
timestamp 1698175906
transform 1 0 22736 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698175906
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_222
timestamp 1698175906
transform 1 0 26208 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_257
timestamp 1698175906
transform 1 0 30128 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_273
timestamp 1698175906
transform 1 0 31920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698175906
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698175906
transform 1 0 4928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 9072 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698175906
transform 1 0 9520 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_75
timestamp 1698175906
transform 1 0 9744 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_114
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_118
timestamp 1698175906
transform 1 0 14560 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_131
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_139
timestamp 1698175906
transform 1 0 16912 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_142
timestamp 1698175906
transform 1 0 17248 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698175906
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_183
timestamp 1698175906
transform 1 0 21840 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_191
timestamp 1698175906
transform 1 0 22736 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_200
timestamp 1698175906
transform 1 0 23744 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_232
timestamp 1698175906
transform 1 0 27328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_242
timestamp 1698175906
transform 1 0 28448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_252
timestamp 1698175906
transform 1 0 29568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_284
timestamp 1698175906
transform 1 0 33152 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_300
timestamp 1698175906
transform 1 0 34944 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_308
timestamp 1698175906
transform 1 0 35840 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698175906
transform 1 0 36288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698175906
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_74
timestamp 1698175906
transform 1 0 9632 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_104
timestamp 1698175906
transform 1 0 12992 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_124
timestamp 1698175906
transform 1 0 15232 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_146
timestamp 1698175906
transform 1 0 17696 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_157
timestamp 1698175906
transform 1 0 18928 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_161
timestamp 1698175906
transform 1 0 19376 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_163
timestamp 1698175906
transform 1 0 19600 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_170
timestamp 1698175906
transform 1 0 20384 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_174
timestamp 1698175906
transform 1 0 20832 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_177
timestamp 1698175906
transform 1 0 21168 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_206
timestamp 1698175906
transform 1 0 24416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698175906
transform 1 0 32256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 40320 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_111
timestamp 1698175906
transform 1 0 13776 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_115
timestamp 1698175906
transform 1 0 14224 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_123
timestamp 1698175906
transform 1 0 15120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_125
timestamp 1698175906
transform 1 0 15344 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_149
timestamp 1698175906
transform 1 0 18032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_227
timestamp 1698175906
transform 1 0 26768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_231
timestamp 1698175906
transform 1 0 27216 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_239
timestamp 1698175906
transform 1 0 28112 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698175906
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_252
timestamp 1698175906
transform 1 0 29568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_284
timestamp 1698175906
transform 1 0 33152 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_300
timestamp 1698175906
transform 1 0 34944 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_308
timestamp 1698175906
transform 1 0 35840 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_312
timestamp 1698175906
transform 1 0 36288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698175906
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 4480 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 8064 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_104
timestamp 1698175906
transform 1 0 12992 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_107
timestamp 1698175906
transform 1 0 13328 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_115
timestamp 1698175906
transform 1 0 14224 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_119
timestamp 1698175906
transform 1 0 14672 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_131
timestamp 1698175906
transform 1 0 16016 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698175906
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_146
timestamp 1698175906
transform 1 0 17696 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_185
timestamp 1698175906
transform 1 0 22064 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_189
timestamp 1698175906
transform 1 0 22512 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_201
timestamp 1698175906
transform 1 0 23856 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_223
timestamp 1698175906
transform 1 0 26320 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_258
timestamp 1698175906
transform 1 0 30240 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_274
timestamp 1698175906
transform 1 0 32032 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 4480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_69
timestamp 1698175906
transform 1 0 9072 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_73
timestamp 1698175906
transform 1 0 9520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_75
timestamp 1698175906
transform 1 0 9744 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_109
timestamp 1698175906
transform 1 0 13552 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_147
timestamp 1698175906
transform 1 0 17808 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_155
timestamp 1698175906
transform 1 0 18704 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_200
timestamp 1698175906
transform 1 0 23744 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_255
timestamp 1698175906
transform 1 0 29904 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_287
timestamp 1698175906
transform 1 0 33488 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_303
timestamp 1698175906
transform 1 0 35280 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 4480 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_80
timestamp 1698175906
transform 1 0 10304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_84
timestamp 1698175906
transform 1 0 10752 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_86
timestamp 1698175906
transform 1 0 10976 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_127
timestamp 1698175906
transform 1 0 15568 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_131
timestamp 1698175906
transform 1 0 16016 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_148
timestamp 1698175906
transform 1 0 17920 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_156
timestamp 1698175906
transform 1 0 18816 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_167
timestamp 1698175906
transform 1 0 20048 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_175
timestamp 1698175906
transform 1 0 20944 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_185
timestamp 1698175906
transform 1 0 22064 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_201
timestamp 1698175906
transform 1 0 23856 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_228
timestamp 1698175906
transform 1 0 26880 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_261
timestamp 1698175906
transform 1 0 30576 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_111
timestamp 1698175906
transform 1 0 13776 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_122
timestamp 1698175906
transform 1 0 15008 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_154
timestamp 1698175906
transform 1 0 18592 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_158
timestamp 1698175906
transform 1 0 19040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_160
timestamp 1698175906
transform 1 0 19264 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_169
timestamp 1698175906
transform 1 0 20272 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_173
timestamp 1698175906
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_227
timestamp 1698175906
transform 1 0 26768 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698175906
transform 1 0 10304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_84
timestamp 1698175906
transform 1 0 10752 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_115
timestamp 1698175906
transform 1 0 14224 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_120
timestamp 1698175906
transform 1 0 14784 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_124
timestamp 1698175906
transform 1 0 15232 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_148
timestamp 1698175906
transform 1 0 17920 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_150
timestamp 1698175906
transform 1 0 18144 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_160
timestamp 1698175906
transform 1 0 19264 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_176
timestamp 1698175906
transform 1 0 21056 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_184
timestamp 1698175906
transform 1 0 21952 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_188
timestamp 1698175906
transform 1 0 22400 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_199
timestamp 1698175906
transform 1 0 23632 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_203
timestamp 1698175906
transform 1 0 24080 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_245
timestamp 1698175906
transform 1 0 28784 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698175906
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_123
timestamp 1698175906
transform 1 0 15120 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_127
timestamp 1698175906
transform 1 0 15568 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_157
timestamp 1698175906
transform 1 0 18928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_161
timestamp 1698175906
transform 1 0 19376 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_165
timestamp 1698175906
transform 1 0 19824 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698175906
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_228
timestamp 1698175906
transform 1 0 26880 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_236
timestamp 1698175906
transform 1 0 27776 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_104
timestamp 1698175906
transform 1 0 12992 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_120
timestamp 1698175906
transform 1 0 14784 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_128
timestamp 1698175906
transform 1 0 15680 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_135
timestamp 1698175906
transform 1 0 16464 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_150
timestamp 1698175906
transform 1 0 18144 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_154
timestamp 1698175906
transform 1 0 18592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_206
timestamp 1698175906
transform 1 0 24416 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_216
timestamp 1698175906
transform 1 0 25536 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_220
timestamp 1698175906
transform 1 0 25984 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_252
timestamp 1698175906
transform 1 0 29568 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_268
timestamp 1698175906
transform 1 0 31360 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 36512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 37408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_115
timestamp 1698175906
transform 1 0 14224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_130
timestamp 1698175906
transform 1 0 15904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_132
timestamp 1698175906
transform 1 0 16128 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_139
timestamp 1698175906
transform 1 0 16912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_141
timestamp 1698175906
transform 1 0 17136 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_171
timestamp 1698175906
transform 1 0 20496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_185
timestamp 1698175906
transform 1 0 22064 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_189
timestamp 1698175906
transform 1 0 22512 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_191
timestamp 1698175906
transform 1 0 22736 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_198
timestamp 1698175906
transform 1 0 23520 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_230
timestamp 1698175906
transform 1 0 27104 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698175906
transform 1 0 28000 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_135
timestamp 1698175906
transform 1 0 16464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698175906
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_144
timestamp 1698175906
transform 1 0 17472 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_174
timestamp 1698175906
transform 1 0 20832 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_178
timestamp 1698175906
transform 1 0 21280 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_123
timestamp 1698175906
transform 1 0 15120 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_153
timestamp 1698175906
transform 1 0 18480 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_169
timestamp 1698175906
transform 1 0 20272 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_173
timestamp 1698175906
transform 1 0 20720 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_168
timestamp 1698175906
transform 1 0 20160 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_195
timestamp 1698175906
transform 1 0 23184 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698175906
transform 1 0 24080 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 25536 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_243
timestamp 1698175906
transform 1 0 28560 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698175906
transform 1 0 32144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_108
timestamp 1698175906
transform 1 0 13440 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698175906
transform 1 0 20832 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_201
timestamp 1698175906
transform 1 0 23856 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_203
timestamp 1698175906
transform 1 0 24080 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita33_26 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 36288 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 25648 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform -1 0 16576 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 4480 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform -1 0 4480 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 20272 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 37520 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 4480 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 18928 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 4480 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 16912 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 15568 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 4480 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 20944 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 37520 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 25536 41200 25648 42000 0 FreeSans 448 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 41200 17472 42000 17584 0 FreeSans 448 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 14784 41200 14896 42000 0 FreeSans 448 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 16128 41200 16240 42000 0 FreeSans 448 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 24192 41200 24304 42000 0 FreeSans 448 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 20160 41200 20272 42000 0 FreeSans 448 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 41200 25536 42000 25648 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 41200 21504 42000 21616 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 18816 41200 18928 42000 0 FreeSans 448 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 15456 41200 15568 42000 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 20832 41200 20944 42000 0 FreeSans 448 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 41200 18816 42000 18928 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal3 18592 26488 18592 26488 0 _000_
rlabel metal2 25984 16184 25984 16184 0 _001_
rlabel metal2 22680 13832 22680 13832 0 _002_
rlabel metal2 24808 22680 24808 22680 0 _003_
rlabel metal2 12152 22512 12152 22512 0 _004_
rlabel metal2 27944 21896 27944 21896 0 _005_
rlabel metal3 13888 24024 13888 24024 0 _006_
rlabel metal2 29288 22736 29288 22736 0 _007_
rlabel metal2 16632 13664 16632 13664 0 _008_
rlabel metal2 22176 26152 22176 26152 0 _009_
rlabel metal2 26488 25200 26488 25200 0 _010_
rlabel metal2 23464 25144 23464 25144 0 _011_
rlabel metal2 22680 12824 22680 12824 0 _012_
rlabel metal2 20440 26096 20440 26096 0 _013_
rlabel metal2 28000 16968 28000 16968 0 _014_
rlabel metal2 27496 18032 27496 18032 0 _015_
rlabel metal2 14728 14112 14728 14112 0 _016_
rlabel metal2 13944 27104 13944 27104 0 _017_
rlabel metal3 17136 24920 17136 24920 0 _018_
rlabel metal2 12152 19600 12152 19600 0 _019_
rlabel metal2 27608 16408 27608 16408 0 _020_
rlabel metal2 15176 18088 15176 18088 0 _021_
rlabel metal2 14280 16240 14280 16240 0 _022_
rlabel metal2 19992 14868 19992 14868 0 _023_
rlabel metal3 13272 20216 13272 20216 0 _024_
rlabel metal2 13384 22736 13384 22736 0 _025_
rlabel metal2 29176 19152 29176 19152 0 _026_
rlabel metal2 14616 20272 14616 20272 0 _027_
rlabel metal2 14728 22624 14728 22624 0 _028_
rlabel metal2 22512 19992 22512 19992 0 _029_
rlabel metal3 14952 23240 14952 23240 0 _030_
rlabel metal2 28056 22456 28056 22456 0 _031_
rlabel metal3 15512 22344 15512 22344 0 _032_
rlabel metal3 19992 26264 19992 26264 0 _033_
rlabel metal2 20216 21952 20216 21952 0 _034_
rlabel metal2 21560 25368 21560 25368 0 _035_
rlabel metal2 20328 22736 20328 22736 0 _036_
rlabel metal2 19208 23632 19208 23632 0 _037_
rlabel metal2 19656 25144 19656 25144 0 _038_
rlabel metal3 28616 22120 28616 22120 0 _039_
rlabel metal3 25312 21560 25312 21560 0 _040_
rlabel metal2 27384 18312 27384 18312 0 _041_
rlabel metal2 23352 23296 23352 23296 0 _042_
rlabel metal3 24528 18424 24528 18424 0 _043_
rlabel metal2 23240 17640 23240 17640 0 _044_
rlabel metal3 23688 15176 23688 15176 0 _045_
rlabel metal2 23800 21952 23800 21952 0 _046_
rlabel metal2 14056 22568 14056 22568 0 _047_
rlabel metal2 28504 22456 28504 22456 0 _048_
rlabel metal2 24360 22064 24360 22064 0 _049_
rlabel metal2 14280 24192 14280 24192 0 _050_
rlabel metal2 26320 21784 26320 21784 0 _051_
rlabel metal2 29568 20776 29568 20776 0 _052_
rlabel metal2 18424 14168 18424 14168 0 _053_
rlabel metal2 23128 27048 23128 27048 0 _054_
rlabel metal2 22568 26824 22568 26824 0 _055_
rlabel metal3 26824 25256 26824 25256 0 _056_
rlabel metal3 23352 25368 23352 25368 0 _057_
rlabel metal3 23968 24696 23968 24696 0 _058_
rlabel metal2 23296 16072 23296 16072 0 _059_
rlabel metal2 22792 15960 22792 15960 0 _060_
rlabel metal2 20216 26264 20216 26264 0 _061_
rlabel metal3 28840 18984 28840 18984 0 _062_
rlabel metal2 28056 17528 28056 17528 0 _063_
rlabel metal2 18200 17192 18200 17192 0 _064_
rlabel metal2 20552 17920 20552 17920 0 _065_
rlabel metal2 19992 16128 19992 16128 0 _066_
rlabel metal2 15568 14728 15568 14728 0 _067_
rlabel metal2 21336 22008 21336 22008 0 _068_
rlabel metal3 19264 19992 19264 19992 0 _069_
rlabel metal2 13832 19824 13832 19824 0 _070_
rlabel metal2 17528 18032 17528 18032 0 _071_
rlabel metal2 17192 17360 17192 17360 0 _072_
rlabel metal2 23128 15344 23128 15344 0 _073_
rlabel metal2 16072 14784 16072 14784 0 _074_
rlabel metal3 18312 18424 18312 18424 0 _075_
rlabel metal2 21448 17640 21448 17640 0 _076_
rlabel metal2 15736 21840 15736 21840 0 _077_
rlabel metal2 19824 21560 19824 21560 0 _078_
rlabel metal2 19768 22960 19768 22960 0 _079_
rlabel metal3 14728 23520 14728 23520 0 _080_
rlabel metal3 18200 25368 18200 25368 0 _081_
rlabel metal3 17248 20104 17248 20104 0 _082_
rlabel metal2 14840 25424 14840 25424 0 _083_
rlabel metal2 15176 26600 15176 26600 0 _084_
rlabel metal2 23240 22176 23240 22176 0 _085_
rlabel metal2 22344 14784 22344 14784 0 _086_
rlabel metal3 19488 23912 19488 23912 0 _087_
rlabel metal2 19488 23352 19488 23352 0 _088_
rlabel metal3 18256 24584 18256 24584 0 _089_
rlabel metal2 15064 17304 15064 17304 0 _090_
rlabel metal2 13608 19600 13608 19600 0 _091_
rlabel metal3 20944 20104 20944 20104 0 _092_
rlabel metal2 20664 22736 20664 22736 0 _093_
rlabel metal2 15848 21392 15848 21392 0 _094_
rlabel metal2 14840 22512 14840 22512 0 _095_
rlabel metal2 21672 16408 21672 16408 0 _096_
rlabel metal3 22680 18424 22680 18424 0 _097_
rlabel metal2 22568 17976 22568 17976 0 _098_
rlabel metal2 15064 20608 15064 20608 0 _099_
rlabel metal2 24136 21728 24136 21728 0 _100_
rlabel metal2 14392 21952 14392 21952 0 _101_
rlabel metal2 13608 20356 13608 20356 0 _102_
rlabel metal3 2478 27608 2478 27608 0 clk
rlabel metal2 23576 21000 23576 21000 0 clknet_0_clk
rlabel metal2 21560 12992 21560 12992 0 clknet_1_0__leaf_clk
rlabel metal2 20776 27440 20776 27440 0 clknet_1_1__leaf_clk
rlabel metal2 22904 14840 22904 14840 0 dut33.count\[0\]
rlabel metal2 19208 19544 19208 19544 0 dut33.count\[1\]
rlabel metal3 17304 17416 17304 17416 0 dut33.count\[2\]
rlabel metal3 18536 16856 18536 16856 0 dut33.count\[3\]
rlabel metal3 26936 21896 26936 21896 0 net1
rlabel metal3 23968 27048 23968 27048 0 net10
rlabel metal2 20440 27160 20440 27160 0 net11
rlabel metal2 4312 25032 4312 25032 0 net12
rlabel metal2 27608 25928 27608 25928 0 net13
rlabel metal3 11704 20664 11704 20664 0 net14
rlabel metal2 30408 21840 30408 21840 0 net15
rlabel metal2 19096 6356 19096 6356 0 net16
rlabel metal2 12936 18480 12936 18480 0 net17
rlabel metal3 18424 38024 18424 38024 0 net18
rlabel metal2 17080 5964 17080 5964 0 net19
rlabel metal2 25704 31920 25704 31920 0 net2
rlabel metal2 15736 31696 15736 31696 0 net20
rlabel metal3 6356 22344 6356 22344 0 net21
rlabel metal2 24528 13048 24528 13048 0 net22
rlabel metal2 20664 29820 20664 29820 0 net23
rlabel metal2 30184 17920 30184 17920 0 net24
rlabel metal2 29960 17920 29960 17920 0 net25
rlabel metal2 35672 2030 35672 2030 0 net26
rlabel metal2 23464 17304 23464 17304 0 net3
rlabel metal2 30072 21896 30072 21896 0 net4
rlabel metal2 16408 32480 16408 32480 0 net5
rlabel metal2 25592 6356 25592 6356 0 net6
rlabel metal2 10024 19264 10024 19264 0 net7
rlabel metal3 16800 28056 16800 28056 0 net8
rlabel metal2 10024 22344 10024 22344 0 net9
rlabel metal3 40642 22904 40642 22904 0 segm[10]
rlabel metal2 25592 39914 25592 39914 0 segm[11]
rlabel metal2 40040 17640 40040 17640 0 segm[12]
rlabel metal2 40040 22344 40040 22344 0 segm[13]
rlabel metal2 14840 39690 14840 39690 0 segm[1]
rlabel metal2 24248 2422 24248 2422 0 segm[2]
rlabel metal3 1358 18872 1358 18872 0 segm[3]
rlabel metal2 16184 39354 16184 39354 0 segm[4]
rlabel metal3 1358 22904 1358 22904 0 segm[5]
rlabel metal2 24248 39746 24248 39746 0 segm[6]
rlabel metal2 20216 39354 20216 39354 0 segm[7]
rlabel metal3 1358 24920 1358 24920 0 segm[8]
rlabel metal2 40040 25816 40040 25816 0 segm[9]
rlabel metal3 1358 20888 1358 20888 0 sel[0]
rlabel metal2 40040 21504 40040 21504 0 sel[10]
rlabel metal2 18872 2422 18872 2422 0 sel[11]
rlabel metal3 1358 18200 1358 18200 0 sel[1]
rlabel metal2 18872 39690 18872 39690 0 sel[2]
rlabel metal2 16856 2086 16856 2086 0 sel[3]
rlabel metal2 15512 38962 15512 38962 0 sel[4]
rlabel metal3 1358 22232 1358 22232 0 sel[5]
rlabel metal2 23576 2198 23576 2198 0 sel[6]
rlabel metal2 20888 39746 20888 39746 0 sel[7]
rlabel metal2 40040 19096 40040 19096 0 sel[8]
rlabel metal3 40642 18200 40642 18200 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
