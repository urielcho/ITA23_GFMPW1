magic
tech gf180mcuD
magscale 1 10
timestamp 1699642417
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 18622 38274 18674 38286
rect 18622 38210 18674 38222
rect 22430 38274 22482 38286
rect 22430 38210 22482 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 29374 38274 29426 38286
rect 29374 38210 29426 38222
rect 17714 37998 17726 38050
rect 17778 37998 17790 38050
rect 21410 37998 21422 38050
rect 21474 37998 21486 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 28578 37998 28590 38050
rect 28642 37998 28654 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 19854 37490 19906 37502
rect 19854 37426 19906 37438
rect 22766 37490 22818 37502
rect 22766 37426 22818 37438
rect 26238 37490 26290 37502
rect 26238 37426 26290 37438
rect 18834 37214 18846 37266
rect 18898 37214 18910 37266
rect 21858 37214 21870 37266
rect 21922 37214 21934 37266
rect 25218 37214 25230 37266
rect 25282 37214 25294 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 18062 36706 18114 36718
rect 18062 36642 18114 36654
rect 22318 36706 22370 36718
rect 22318 36642 22370 36654
rect 17266 36430 17278 36482
rect 17330 36430 17342 36482
rect 21298 36430 21310 36482
rect 21362 36430 21374 36482
rect 24334 36258 24386 36270
rect 24334 36194 24386 36206
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 21198 28642 21250 28654
rect 21198 28578 21250 28590
rect 21422 28530 21474 28542
rect 21422 28466 21474 28478
rect 21534 28530 21586 28542
rect 21534 28466 21586 28478
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 18498 27806 18510 27858
rect 18562 27806 18574 27858
rect 21858 27806 21870 27858
rect 21922 27806 21934 27858
rect 16158 27746 16210 27758
rect 16158 27682 16210 27694
rect 17502 27746 17554 27758
rect 17502 27682 17554 27694
rect 18286 27746 18338 27758
rect 19282 27694 19294 27746
rect 19346 27694 19358 27746
rect 21410 27694 21422 27746
rect 21474 27694 21486 27746
rect 22530 27694 22542 27746
rect 22594 27694 22606 27746
rect 24658 27694 24670 27746
rect 24722 27694 24734 27746
rect 18286 27682 18338 27694
rect 16046 27634 16098 27646
rect 16046 27570 16098 27582
rect 17390 27634 17442 27646
rect 17390 27570 17442 27582
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 23102 27298 23154 27310
rect 23102 27234 23154 27246
rect 16370 27134 16382 27186
rect 16434 27134 16446 27186
rect 18498 27134 18510 27186
rect 18562 27134 18574 27186
rect 19966 27074 20018 27086
rect 15698 27022 15710 27074
rect 15762 27022 15774 27074
rect 19966 27010 20018 27022
rect 21646 27074 21698 27086
rect 21646 27010 21698 27022
rect 22990 27074 23042 27086
rect 22990 27010 23042 27022
rect 24110 27074 24162 27086
rect 24110 27010 24162 27022
rect 18958 26962 19010 26974
rect 18958 26898 19010 26910
rect 19630 26962 19682 26974
rect 19630 26898 19682 26910
rect 19742 26962 19794 26974
rect 19742 26898 19794 26910
rect 21310 26962 21362 26974
rect 21310 26898 21362 26910
rect 21870 26962 21922 26974
rect 21870 26898 21922 26910
rect 21982 26962 22034 26974
rect 21982 26898 22034 26910
rect 23102 26962 23154 26974
rect 23102 26898 23154 26910
rect 23774 26962 23826 26974
rect 23774 26898 23826 26910
rect 23998 26962 24050 26974
rect 23998 26898 24050 26910
rect 21422 26850 21474 26862
rect 21422 26786 21474 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 17390 26514 17442 26526
rect 18398 26514 18450 26526
rect 17714 26462 17726 26514
rect 17778 26462 17790 26514
rect 17390 26450 17442 26462
rect 18398 26450 18450 26462
rect 18622 26514 18674 26526
rect 18622 26450 18674 26462
rect 25342 26514 25394 26526
rect 25342 26450 25394 26462
rect 25230 26402 25282 26414
rect 14690 26350 14702 26402
rect 14754 26350 14766 26402
rect 21746 26350 21758 26402
rect 21810 26350 21822 26402
rect 25230 26338 25282 26350
rect 18734 26290 18786 26302
rect 14018 26238 14030 26290
rect 14082 26238 14094 26290
rect 18162 26238 18174 26290
rect 18226 26238 18238 26290
rect 22530 26238 22542 26290
rect 22594 26238 22606 26290
rect 18734 26226 18786 26238
rect 16818 26126 16830 26178
rect 16882 26126 16894 26178
rect 18386 26126 18398 26178
rect 18450 26126 18462 26178
rect 19618 26126 19630 26178
rect 19682 26126 19694 26178
rect 25342 26066 25394 26078
rect 25342 26002 25394 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 1934 25618 1986 25630
rect 17378 25566 17390 25618
rect 17442 25566 17454 25618
rect 21746 25566 21758 25618
rect 21810 25566 21822 25618
rect 26450 25566 26462 25618
rect 26514 25566 26526 25618
rect 1934 25554 1986 25566
rect 17502 25506 17554 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 17502 25442 17554 25454
rect 18846 25506 18898 25518
rect 20178 25454 20190 25506
rect 20242 25454 20254 25506
rect 23650 25454 23662 25506
rect 23714 25454 23726 25506
rect 18846 25442 18898 25454
rect 17950 25394 18002 25406
rect 17950 25330 18002 25342
rect 18510 25394 18562 25406
rect 21310 25394 21362 25406
rect 20402 25342 20414 25394
rect 20466 25342 20478 25394
rect 18510 25330 18562 25342
rect 21310 25330 21362 25342
rect 21758 25394 21810 25406
rect 21758 25330 21810 25342
rect 21870 25394 21922 25406
rect 24322 25342 24334 25394
rect 24386 25342 24398 25394
rect 21870 25330 21922 25342
rect 16942 25282 16994 25294
rect 16942 25218 16994 25230
rect 17390 25282 17442 25294
rect 17390 25218 17442 25230
rect 17726 25282 17778 25294
rect 17726 25218 17778 25230
rect 18622 25282 18674 25294
rect 18622 25218 18674 25230
rect 21534 25282 21586 25294
rect 21534 25218 21586 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 24110 24946 24162 24958
rect 15474 24894 15486 24946
rect 15538 24894 15550 24946
rect 24110 24882 24162 24894
rect 24334 24834 24386 24846
rect 24334 24770 24386 24782
rect 24446 24834 24498 24846
rect 24446 24770 24498 24782
rect 4274 24670 4286 24722
rect 4338 24670 4350 24722
rect 15138 24670 15150 24722
rect 15202 24670 15214 24722
rect 15698 24670 15710 24722
rect 15762 24670 15774 24722
rect 16270 24610 16322 24622
rect 12226 24558 12238 24610
rect 12290 24558 12302 24610
rect 14354 24558 14366 24610
rect 14418 24558 14430 24610
rect 16270 24546 16322 24558
rect 17502 24610 17554 24622
rect 17502 24546 17554 24558
rect 1934 24498 1986 24510
rect 1934 24434 1986 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 1934 24050 1986 24062
rect 1934 23986 1986 23998
rect 17054 24050 17106 24062
rect 20402 23998 20414 24050
rect 20466 23998 20478 24050
rect 17054 23986 17106 23998
rect 15822 23938 15874 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 15026 23886 15038 23938
rect 15090 23886 15102 23938
rect 15822 23874 15874 23886
rect 16158 23938 16210 23950
rect 16158 23874 16210 23886
rect 16606 23938 16658 23950
rect 16606 23874 16658 23886
rect 16718 23938 16770 23950
rect 16718 23874 16770 23886
rect 16942 23938 16994 23950
rect 25454 23938 25506 23950
rect 17490 23886 17502 23938
rect 17554 23886 17566 23938
rect 16942 23874 16994 23886
rect 25454 23874 25506 23886
rect 26238 23938 26290 23950
rect 26238 23874 26290 23886
rect 15486 23826 15538 23838
rect 14802 23774 14814 23826
rect 14866 23774 14878 23826
rect 15486 23762 15538 23774
rect 15598 23826 15650 23838
rect 15598 23762 15650 23774
rect 17166 23826 17218 23838
rect 25118 23826 25170 23838
rect 18274 23774 18286 23826
rect 18338 23774 18350 23826
rect 17166 23762 17218 23774
rect 25118 23762 25170 23774
rect 25678 23826 25730 23838
rect 25678 23762 25730 23774
rect 26574 23826 26626 23838
rect 26574 23762 26626 23774
rect 21422 23714 21474 23726
rect 21422 23650 21474 23662
rect 25342 23714 25394 23726
rect 25342 23650 25394 23662
rect 26462 23714 26514 23726
rect 26462 23650 26514 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 17390 23378 17442 23390
rect 20190 23378 20242 23390
rect 18946 23326 18958 23378
rect 19010 23326 19022 23378
rect 17390 23314 17442 23326
rect 20190 23314 20242 23326
rect 20414 23378 20466 23390
rect 20414 23314 20466 23326
rect 14814 23266 14866 23278
rect 14814 23202 14866 23214
rect 17502 23266 17554 23278
rect 17502 23202 17554 23214
rect 18510 23266 18562 23278
rect 26002 23214 26014 23266
rect 26066 23214 26078 23266
rect 18510 23202 18562 23214
rect 14702 23154 14754 23166
rect 18062 23154 18114 23166
rect 4274 23102 4286 23154
rect 4338 23102 4350 23154
rect 14242 23102 14254 23154
rect 14306 23102 14318 23154
rect 17714 23102 17726 23154
rect 17778 23102 17790 23154
rect 14702 23090 14754 23102
rect 18062 23090 18114 23102
rect 18398 23154 18450 23166
rect 18398 23090 18450 23102
rect 18958 23154 19010 23166
rect 18958 23090 19010 23102
rect 19182 23154 19234 23166
rect 19182 23090 19234 23102
rect 19406 23154 19458 23166
rect 19406 23090 19458 23102
rect 19518 23154 19570 23166
rect 19954 23102 19966 23154
rect 20018 23102 20030 23154
rect 20626 23102 20638 23154
rect 20690 23102 20702 23154
rect 21074 23102 21086 23154
rect 21138 23102 21150 23154
rect 25330 23102 25342 23154
rect 25394 23102 25406 23154
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 19518 23090 19570 23102
rect 15374 23042 15426 23054
rect 11442 22990 11454 23042
rect 11506 22990 11518 23042
rect 13570 22990 13582 23042
rect 13634 22990 13646 23042
rect 20514 22990 20526 23042
rect 20578 22990 20590 23042
rect 21746 22990 21758 23042
rect 21810 22990 21822 23042
rect 23874 22990 23886 23042
rect 23938 22990 23950 23042
rect 28130 22990 28142 23042
rect 28194 22990 28206 23042
rect 15374 22978 15426 22990
rect 1934 22930 1986 22942
rect 1934 22866 1986 22878
rect 14814 22930 14866 22942
rect 14814 22866 14866 22878
rect 18510 22930 18562 22942
rect 18510 22866 18562 22878
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 19630 22594 19682 22606
rect 19630 22530 19682 22542
rect 21646 22594 21698 22606
rect 21646 22530 21698 22542
rect 1934 22482 1986 22494
rect 1934 22418 1986 22430
rect 21758 22482 21810 22494
rect 40014 22482 40066 22494
rect 28578 22430 28590 22482
rect 28642 22430 28654 22482
rect 21758 22418 21810 22430
rect 40014 22418 40066 22430
rect 14366 22370 14418 22382
rect 19854 22370 19906 22382
rect 4274 22318 4286 22370
rect 4338 22318 4350 22370
rect 18722 22318 18734 22370
rect 18786 22318 18798 22370
rect 14366 22306 14418 22318
rect 19854 22306 19906 22318
rect 20190 22370 20242 22382
rect 21970 22318 21982 22370
rect 22034 22318 22046 22370
rect 25778 22318 25790 22370
rect 25842 22318 25854 22370
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 20190 22306 20242 22318
rect 14030 22258 14082 22270
rect 14030 22194 14082 22206
rect 14142 22258 14194 22270
rect 14142 22194 14194 22206
rect 14702 22258 14754 22270
rect 19294 22258 19346 22270
rect 17826 22206 17838 22258
rect 17890 22206 17902 22258
rect 14702 22194 14754 22206
rect 19294 22194 19346 22206
rect 23550 22258 23602 22270
rect 26450 22206 26462 22258
rect 26514 22206 26526 22258
rect 23550 22194 23602 22206
rect 18174 22146 18226 22158
rect 19518 22146 19570 22158
rect 18498 22094 18510 22146
rect 18562 22094 18574 22146
rect 18174 22082 18226 22094
rect 19518 22082 19570 22094
rect 20078 22146 20130 22158
rect 20078 22082 20130 22094
rect 23662 22146 23714 22158
rect 23662 22082 23714 22094
rect 23886 22146 23938 22158
rect 23886 22082 23938 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 15038 21810 15090 21822
rect 18834 21758 18846 21810
rect 18898 21758 18910 21810
rect 25554 21758 25566 21810
rect 25618 21758 25630 21810
rect 26450 21758 26462 21810
rect 26514 21758 26526 21810
rect 15038 21746 15090 21758
rect 14814 21698 14866 21710
rect 14814 21634 14866 21646
rect 15486 21698 15538 21710
rect 15486 21634 15538 21646
rect 15598 21698 15650 21710
rect 26686 21698 26738 21710
rect 18386 21646 18398 21698
rect 18450 21646 18462 21698
rect 15598 21634 15650 21646
rect 26686 21634 26738 21646
rect 27806 21698 27858 21710
rect 27806 21634 27858 21646
rect 14478 21586 14530 21598
rect 14242 21534 14254 21586
rect 14306 21534 14318 21586
rect 14478 21522 14530 21534
rect 15262 21586 15314 21598
rect 15262 21522 15314 21534
rect 17614 21586 17666 21598
rect 25230 21586 25282 21598
rect 27694 21586 27746 21598
rect 18274 21534 18286 21586
rect 18338 21534 18350 21586
rect 19058 21534 19070 21586
rect 19122 21534 19134 21586
rect 19394 21534 19406 21586
rect 19458 21534 19470 21586
rect 25890 21534 25902 21586
rect 25954 21534 25966 21586
rect 26450 21534 26462 21586
rect 26514 21534 26526 21586
rect 37874 21534 37886 21586
rect 37938 21534 37950 21586
rect 17614 21522 17666 21534
rect 25230 21522 25282 21534
rect 27694 21522 27746 21534
rect 11330 21422 11342 21474
rect 11394 21422 11406 21474
rect 13458 21422 13470 21474
rect 13522 21422 13534 21474
rect 22866 21422 22878 21474
rect 22930 21422 22942 21474
rect 39890 21422 39902 21474
rect 39954 21422 39966 21474
rect 14702 21362 14754 21374
rect 26114 21310 26126 21362
rect 26178 21310 26190 21362
rect 14702 21298 14754 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 14926 21026 14978 21038
rect 14926 20962 14978 20974
rect 21198 21026 21250 21038
rect 21198 20962 21250 20974
rect 40014 20914 40066 20926
rect 40014 20850 40066 20862
rect 14030 20802 14082 20814
rect 14030 20738 14082 20750
rect 14366 20802 14418 20814
rect 14366 20738 14418 20750
rect 15150 20802 15202 20814
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 22194 20750 22206 20802
rect 22258 20750 22270 20802
rect 22866 20750 22878 20802
rect 22930 20750 22942 20802
rect 37986 20750 37998 20802
rect 38050 20750 38062 20802
rect 15150 20738 15202 20750
rect 14142 20690 14194 20702
rect 21534 20690 21586 20702
rect 15698 20638 15710 20690
rect 15762 20638 15774 20690
rect 14142 20626 14194 20638
rect 21534 20626 21586 20638
rect 21758 20690 21810 20702
rect 22418 20638 22430 20690
rect 22482 20638 22494 20690
rect 25778 20638 25790 20690
rect 25842 20638 25854 20690
rect 21758 20626 21810 20638
rect 21310 20578 21362 20590
rect 14578 20526 14590 20578
rect 14642 20526 14654 20578
rect 21310 20514 21362 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 22206 20242 22258 20254
rect 22206 20178 22258 20190
rect 13246 20130 13298 20142
rect 13246 20066 13298 20078
rect 13582 20130 13634 20142
rect 21646 20130 21698 20142
rect 17490 20078 17502 20130
rect 17554 20078 17566 20130
rect 18946 20078 18958 20130
rect 19010 20078 19022 20130
rect 13582 20066 13634 20078
rect 21646 20066 21698 20078
rect 22094 20130 22146 20142
rect 22094 20066 22146 20078
rect 23998 20130 24050 20142
rect 23998 20066 24050 20078
rect 24222 20130 24274 20142
rect 24222 20066 24274 20078
rect 25566 20130 25618 20142
rect 25566 20066 25618 20078
rect 25678 20130 25730 20142
rect 25678 20066 25730 20078
rect 26462 20130 26514 20142
rect 26462 20066 26514 20078
rect 27246 20130 27298 20142
rect 27246 20066 27298 20078
rect 27358 20130 27410 20142
rect 27358 20066 27410 20078
rect 29262 20130 29314 20142
rect 29262 20066 29314 20078
rect 17838 20018 17890 20030
rect 20526 20018 20578 20030
rect 21310 20018 21362 20030
rect 23774 20018 23826 20030
rect 18498 19966 18510 20018
rect 18562 19966 18574 20018
rect 18834 19966 18846 20018
rect 18898 19966 18910 20018
rect 19730 19966 19742 20018
rect 19794 19966 19806 20018
rect 20738 19966 20750 20018
rect 20802 19966 20814 20018
rect 21858 19966 21870 20018
rect 21922 19966 21934 20018
rect 17838 19954 17890 19966
rect 20526 19954 20578 19966
rect 21310 19954 21362 19966
rect 23774 19954 23826 19966
rect 24446 20018 24498 20030
rect 24446 19954 24498 19966
rect 25342 20018 25394 20030
rect 27022 20018 27074 20030
rect 26674 19966 26686 20018
rect 26738 19966 26750 20018
rect 25342 19954 25394 19966
rect 27022 19954 27074 19966
rect 29598 20018 29650 20030
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 29598 19954 29650 19966
rect 18386 19854 18398 19906
rect 18450 19854 18462 19906
rect 19506 19854 19518 19906
rect 19570 19854 19582 19906
rect 26450 19854 26462 19906
rect 26514 19854 26526 19906
rect 18174 19794 18226 19806
rect 18174 19730 18226 19742
rect 24334 19794 24386 19806
rect 24334 19730 24386 19742
rect 27358 19794 27410 19806
rect 27358 19730 27410 19742
rect 40014 19794 40066 19806
rect 40014 19730 40066 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 20638 19458 20690 19470
rect 17714 19406 17726 19458
rect 17778 19406 17790 19458
rect 19506 19406 19518 19458
rect 19570 19406 19582 19458
rect 20638 19394 20690 19406
rect 40014 19346 40066 19358
rect 20066 19294 20078 19346
rect 20130 19294 20142 19346
rect 24098 19294 24110 19346
rect 24162 19294 24174 19346
rect 26226 19294 26238 19346
rect 26290 19294 26302 19346
rect 40014 19282 40066 19294
rect 16606 19234 16658 19246
rect 15810 19182 15822 19234
rect 15874 19182 15886 19234
rect 16606 19170 16658 19182
rect 17054 19234 17106 19246
rect 17054 19170 17106 19182
rect 17502 19234 17554 19246
rect 27470 19234 27522 19246
rect 18498 19182 18510 19234
rect 18562 19182 18574 19234
rect 19954 19182 19966 19234
rect 20018 19182 20030 19234
rect 23314 19182 23326 19234
rect 23378 19182 23390 19234
rect 29250 19182 29262 19234
rect 29314 19182 29326 19234
rect 29922 19182 29934 19234
rect 29986 19182 29998 19234
rect 37650 19182 37662 19234
rect 37714 19182 37726 19234
rect 17502 19170 17554 19182
rect 27470 19170 27522 19182
rect 20526 19122 20578 19134
rect 14914 19070 14926 19122
rect 14978 19070 14990 19122
rect 20526 19058 20578 19070
rect 21310 19122 21362 19134
rect 21310 19058 21362 19070
rect 21422 19122 21474 19134
rect 29474 19070 29486 19122
rect 29538 19070 29550 19122
rect 21422 19058 21474 19070
rect 15262 19010 15314 19022
rect 20638 19010 20690 19022
rect 15586 18958 15598 19010
rect 15650 18958 15662 19010
rect 16258 18958 16270 19010
rect 16322 18958 16334 19010
rect 18722 18958 18734 19010
rect 18786 18958 18798 19010
rect 15262 18946 15314 18958
rect 20638 18946 20690 18958
rect 21646 19010 21698 19022
rect 21646 18946 21698 18958
rect 27582 19010 27634 19022
rect 27582 18946 27634 18958
rect 27806 19010 27858 19022
rect 30146 18958 30158 19010
rect 30210 18958 30222 19010
rect 27806 18946 27858 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 15710 18674 15762 18686
rect 15710 18610 15762 18622
rect 16270 18674 16322 18686
rect 16270 18610 16322 18622
rect 17614 18562 17666 18574
rect 12674 18510 12686 18562
rect 12738 18510 12750 18562
rect 17614 18498 17666 18510
rect 18398 18562 18450 18574
rect 26450 18510 26462 18562
rect 26514 18510 26526 18562
rect 29362 18510 29374 18562
rect 29426 18510 29438 18562
rect 18398 18498 18450 18510
rect 15486 18450 15538 18462
rect 4274 18398 4286 18450
rect 4338 18398 4350 18450
rect 12002 18398 12014 18450
rect 12066 18398 12078 18450
rect 15138 18398 15150 18450
rect 15202 18398 15214 18450
rect 15486 18386 15538 18398
rect 17838 18450 17890 18462
rect 17838 18386 17890 18398
rect 19518 18450 19570 18462
rect 19518 18386 19570 18398
rect 21086 18450 21138 18462
rect 21298 18398 21310 18450
rect 21362 18398 21374 18450
rect 22082 18398 22094 18450
rect 22146 18398 22158 18450
rect 25666 18398 25678 18450
rect 25730 18398 25742 18450
rect 29138 18398 29150 18450
rect 29202 18398 29214 18450
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 21086 18386 21138 18398
rect 15598 18338 15650 18350
rect 14802 18286 14814 18338
rect 14866 18286 14878 18338
rect 15598 18274 15650 18286
rect 16382 18338 16434 18350
rect 16382 18274 16434 18286
rect 16718 18338 16770 18350
rect 16718 18274 16770 18286
rect 17726 18338 17778 18350
rect 18498 18286 18510 18338
rect 18562 18286 18574 18338
rect 20738 18286 20750 18338
rect 20802 18286 20814 18338
rect 21970 18286 21982 18338
rect 22034 18286 22046 18338
rect 28578 18286 28590 18338
rect 28642 18286 28654 18338
rect 17726 18274 17778 18286
rect 1934 18226 1986 18238
rect 1934 18162 1986 18174
rect 16830 18226 16882 18238
rect 16830 18162 16882 18174
rect 18174 18226 18226 18238
rect 18174 18162 18226 18174
rect 19406 18226 19458 18238
rect 40014 18226 40066 18238
rect 20626 18174 20638 18226
rect 20690 18174 20702 18226
rect 22306 18174 22318 18226
rect 22370 18174 22382 18226
rect 19406 18162 19458 18174
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 14254 17890 14306 17902
rect 14254 17826 14306 17838
rect 16270 17890 16322 17902
rect 16270 17826 16322 17838
rect 20414 17890 20466 17902
rect 20414 17826 20466 17838
rect 23774 17890 23826 17902
rect 23774 17826 23826 17838
rect 24110 17890 24162 17902
rect 24110 17826 24162 17838
rect 40014 17778 40066 17790
rect 9986 17726 9998 17778
rect 10050 17726 10062 17778
rect 12114 17726 12126 17778
rect 12178 17726 12190 17778
rect 14018 17726 14030 17778
rect 14082 17726 14094 17778
rect 40014 17714 40066 17726
rect 13582 17666 13634 17678
rect 15038 17666 15090 17678
rect 12786 17614 12798 17666
rect 12850 17614 12862 17666
rect 13906 17614 13918 17666
rect 13970 17614 13982 17666
rect 13582 17602 13634 17614
rect 15038 17602 15090 17614
rect 16494 17666 16546 17678
rect 17278 17666 17330 17678
rect 16706 17614 16718 17666
rect 16770 17614 16782 17666
rect 16494 17602 16546 17614
rect 17278 17602 17330 17614
rect 17950 17666 18002 17678
rect 17950 17602 18002 17614
rect 18622 17666 18674 17678
rect 21310 17666 21362 17678
rect 19618 17614 19630 17666
rect 19682 17614 19694 17666
rect 20402 17614 20414 17666
rect 20466 17614 20478 17666
rect 18622 17602 18674 17614
rect 21310 17602 21362 17614
rect 21534 17666 21586 17678
rect 21534 17602 21586 17614
rect 21982 17666 22034 17678
rect 26462 17666 26514 17678
rect 23762 17614 23774 17666
rect 23826 17614 23838 17666
rect 21982 17602 22034 17614
rect 26462 17602 26514 17614
rect 26686 17666 26738 17678
rect 27122 17614 27134 17666
rect 27186 17614 27198 17666
rect 27682 17614 27694 17666
rect 27746 17614 27758 17666
rect 37874 17614 37886 17666
rect 37938 17614 37950 17666
rect 26686 17602 26738 17614
rect 16158 17554 16210 17566
rect 20078 17554 20130 17566
rect 21422 17554 21474 17566
rect 17602 17502 17614 17554
rect 17666 17502 17678 17554
rect 18274 17502 18286 17554
rect 18338 17502 18350 17554
rect 18946 17502 18958 17554
rect 19010 17502 19022 17554
rect 19394 17502 19406 17554
rect 19458 17502 19470 17554
rect 20514 17502 20526 17554
rect 20578 17551 20590 17554
rect 20850 17551 20862 17554
rect 20578 17505 20862 17551
rect 20578 17502 20590 17505
rect 20850 17502 20862 17505
rect 20914 17502 20926 17554
rect 16158 17490 16210 17502
rect 20078 17490 20130 17502
rect 21422 17490 21474 17502
rect 26574 17554 26626 17566
rect 26574 17490 26626 17502
rect 27470 17442 27522 17454
rect 27470 17378 27522 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 17502 17106 17554 17118
rect 20302 17106 20354 17118
rect 18050 17054 18062 17106
rect 18114 17054 18126 17106
rect 17502 17042 17554 17054
rect 20302 17042 20354 17054
rect 20526 17106 20578 17118
rect 20526 17042 20578 17054
rect 23774 17106 23826 17118
rect 23774 17042 23826 17054
rect 23438 16994 23490 17006
rect 14354 16942 14366 16994
rect 14418 16942 14430 16994
rect 23438 16930 23490 16942
rect 23886 16994 23938 17006
rect 23886 16930 23938 16942
rect 25230 16994 25282 17006
rect 25554 16942 25566 16994
rect 25618 16942 25630 16994
rect 27122 16942 27134 16994
rect 27186 16942 27198 16994
rect 25230 16930 25282 16942
rect 18398 16882 18450 16894
rect 13570 16830 13582 16882
rect 13634 16830 13646 16882
rect 18398 16818 18450 16830
rect 18622 16882 18674 16894
rect 18622 16818 18674 16830
rect 20190 16882 20242 16894
rect 22094 16882 22146 16894
rect 21634 16830 21646 16882
rect 21698 16830 21710 16882
rect 20190 16818 20242 16830
rect 22094 16818 22146 16830
rect 22430 16882 22482 16894
rect 23662 16882 23714 16894
rect 23090 16830 23102 16882
rect 23154 16830 23166 16882
rect 22430 16818 22482 16830
rect 23662 16818 23714 16830
rect 23998 16882 24050 16894
rect 26338 16830 26350 16882
rect 26402 16830 26414 16882
rect 37650 16830 37662 16882
rect 37714 16830 37726 16882
rect 23998 16818 24050 16830
rect 22878 16770 22930 16782
rect 16482 16718 16494 16770
rect 16546 16718 16558 16770
rect 21970 16718 21982 16770
rect 22034 16718 22046 16770
rect 29250 16718 29262 16770
rect 29314 16718 29326 16770
rect 22878 16706 22930 16718
rect 22766 16658 22818 16670
rect 22766 16594 22818 16606
rect 40014 16658 40066 16670
rect 40014 16594 40066 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 20526 16322 20578 16334
rect 20526 16258 20578 16270
rect 28254 16322 28306 16334
rect 28254 16258 28306 16270
rect 28366 16210 28418 16222
rect 23874 16158 23886 16210
rect 23938 16158 23950 16210
rect 26002 16158 26014 16210
rect 26066 16158 26078 16210
rect 28366 16146 28418 16158
rect 19630 16098 19682 16110
rect 19394 16046 19406 16098
rect 19458 16046 19470 16098
rect 19630 16034 19682 16046
rect 22094 16098 22146 16110
rect 22094 16034 22146 16046
rect 22654 16098 22706 16110
rect 23090 16046 23102 16098
rect 23154 16046 23166 16098
rect 22654 16034 22706 16046
rect 20414 15986 20466 15998
rect 20414 15922 20466 15934
rect 22542 15986 22594 15998
rect 22542 15922 22594 15934
rect 19966 15874 20018 15886
rect 19966 15810 20018 15822
rect 22430 15874 22482 15886
rect 22430 15810 22482 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 18834 15486 18846 15538
rect 18898 15486 18910 15538
rect 20750 15426 20802 15438
rect 20066 15374 20078 15426
rect 20130 15374 20142 15426
rect 20750 15362 20802 15374
rect 20862 15426 20914 15438
rect 22530 15374 22542 15426
rect 22594 15374 22606 15426
rect 20862 15362 20914 15374
rect 18510 15314 18562 15326
rect 18510 15250 18562 15262
rect 19182 15314 19234 15326
rect 19182 15250 19234 15262
rect 19406 15314 19458 15326
rect 20290 15262 20302 15314
rect 20354 15262 20366 15314
rect 21858 15262 21870 15314
rect 21922 15262 21934 15314
rect 19406 15250 19458 15262
rect 18050 15150 18062 15202
rect 18114 15150 18126 15202
rect 24658 15150 24670 15202
rect 24722 15150 24734 15202
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 16818 14590 16830 14642
rect 16882 14590 16894 14642
rect 18946 14590 18958 14642
rect 19010 14590 19022 14642
rect 19618 14590 19630 14642
rect 19682 14590 19694 14642
rect 21310 14530 21362 14542
rect 16146 14478 16158 14530
rect 16210 14478 16222 14530
rect 19954 14478 19966 14530
rect 20018 14478 20030 14530
rect 21310 14466 21362 14478
rect 19294 14418 19346 14430
rect 21634 14366 21646 14418
rect 21698 14366 21710 14418
rect 19294 14354 19346 14366
rect 20750 14306 20802 14318
rect 20750 14242 20802 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 16830 13970 16882 13982
rect 16830 13906 16882 13918
rect 17826 13694 17838 13746
rect 17890 13694 17902 13746
rect 18498 13582 18510 13634
rect 18562 13582 18574 13634
rect 20626 13582 20638 13634
rect 20690 13582 20702 13634
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 18846 12962 18898 12974
rect 18846 12898 18898 12910
rect 18510 12850 18562 12862
rect 18510 12786 18562 12798
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 25218 4286 25230 4338
rect 25282 4286 25294 4338
rect 26238 4114 26290 4126
rect 26238 4050 26290 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 18622 38222 18674 38274
rect 22430 38222 22482 38274
rect 25566 38222 25618 38274
rect 29374 38222 29426 38274
rect 17726 37998 17778 38050
rect 21422 37998 21474 38050
rect 24558 37998 24610 38050
rect 28590 37998 28642 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 19854 37438 19906 37490
rect 22766 37438 22818 37490
rect 26238 37438 26290 37490
rect 18846 37214 18898 37266
rect 21870 37214 21922 37266
rect 25230 37214 25282 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 18062 36654 18114 36706
rect 22318 36654 22370 36706
rect 17278 36430 17330 36482
rect 21310 36430 21362 36482
rect 24334 36206 24386 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 21198 28590 21250 28642
rect 21422 28478 21474 28530
rect 21534 28478 21586 28530
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 18510 27806 18562 27858
rect 21870 27806 21922 27858
rect 16158 27694 16210 27746
rect 17502 27694 17554 27746
rect 18286 27694 18338 27746
rect 19294 27694 19346 27746
rect 21422 27694 21474 27746
rect 22542 27694 22594 27746
rect 24670 27694 24722 27746
rect 16046 27582 16098 27634
rect 17390 27582 17442 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 23102 27246 23154 27298
rect 16382 27134 16434 27186
rect 18510 27134 18562 27186
rect 15710 27022 15762 27074
rect 19966 27022 20018 27074
rect 21646 27022 21698 27074
rect 22990 27022 23042 27074
rect 24110 27022 24162 27074
rect 18958 26910 19010 26962
rect 19630 26910 19682 26962
rect 19742 26910 19794 26962
rect 21310 26910 21362 26962
rect 21870 26910 21922 26962
rect 21982 26910 22034 26962
rect 23102 26910 23154 26962
rect 23774 26910 23826 26962
rect 23998 26910 24050 26962
rect 21422 26798 21474 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 17390 26462 17442 26514
rect 17726 26462 17778 26514
rect 18398 26462 18450 26514
rect 18622 26462 18674 26514
rect 25342 26462 25394 26514
rect 14702 26350 14754 26402
rect 21758 26350 21810 26402
rect 25230 26350 25282 26402
rect 14030 26238 14082 26290
rect 18174 26238 18226 26290
rect 18734 26238 18786 26290
rect 22542 26238 22594 26290
rect 16830 26126 16882 26178
rect 18398 26126 18450 26178
rect 19630 26126 19682 26178
rect 25342 26014 25394 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 1934 25566 1986 25618
rect 17390 25566 17442 25618
rect 21758 25566 21810 25618
rect 26462 25566 26514 25618
rect 4286 25454 4338 25506
rect 17502 25454 17554 25506
rect 18846 25454 18898 25506
rect 20190 25454 20242 25506
rect 23662 25454 23714 25506
rect 17950 25342 18002 25394
rect 18510 25342 18562 25394
rect 20414 25342 20466 25394
rect 21310 25342 21362 25394
rect 21758 25342 21810 25394
rect 21870 25342 21922 25394
rect 24334 25342 24386 25394
rect 16942 25230 16994 25282
rect 17390 25230 17442 25282
rect 17726 25230 17778 25282
rect 18622 25230 18674 25282
rect 21534 25230 21586 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 15486 24894 15538 24946
rect 24110 24894 24162 24946
rect 24334 24782 24386 24834
rect 24446 24782 24498 24834
rect 4286 24670 4338 24722
rect 15150 24670 15202 24722
rect 15710 24670 15762 24722
rect 12238 24558 12290 24610
rect 14366 24558 14418 24610
rect 16270 24558 16322 24610
rect 17502 24558 17554 24610
rect 1934 24446 1986 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 1934 23998 1986 24050
rect 17054 23998 17106 24050
rect 20414 23998 20466 24050
rect 4286 23886 4338 23938
rect 15038 23886 15090 23938
rect 15822 23886 15874 23938
rect 16158 23886 16210 23938
rect 16606 23886 16658 23938
rect 16718 23886 16770 23938
rect 16942 23886 16994 23938
rect 17502 23886 17554 23938
rect 25454 23886 25506 23938
rect 26238 23886 26290 23938
rect 14814 23774 14866 23826
rect 15486 23774 15538 23826
rect 15598 23774 15650 23826
rect 17166 23774 17218 23826
rect 18286 23774 18338 23826
rect 25118 23774 25170 23826
rect 25678 23774 25730 23826
rect 26574 23774 26626 23826
rect 21422 23662 21474 23714
rect 25342 23662 25394 23714
rect 26462 23662 26514 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 17390 23326 17442 23378
rect 18958 23326 19010 23378
rect 20190 23326 20242 23378
rect 20414 23326 20466 23378
rect 14814 23214 14866 23266
rect 17502 23214 17554 23266
rect 18510 23214 18562 23266
rect 26014 23214 26066 23266
rect 4286 23102 4338 23154
rect 14254 23102 14306 23154
rect 14702 23102 14754 23154
rect 17726 23102 17778 23154
rect 18062 23102 18114 23154
rect 18398 23102 18450 23154
rect 18958 23102 19010 23154
rect 19182 23102 19234 23154
rect 19406 23102 19458 23154
rect 19518 23102 19570 23154
rect 19966 23102 20018 23154
rect 20638 23102 20690 23154
rect 21086 23102 21138 23154
rect 25342 23102 25394 23154
rect 37662 23102 37714 23154
rect 11454 22990 11506 23042
rect 13582 22990 13634 23042
rect 15374 22990 15426 23042
rect 20526 22990 20578 23042
rect 21758 22990 21810 23042
rect 23886 22990 23938 23042
rect 28142 22990 28194 23042
rect 1934 22878 1986 22930
rect 14814 22878 14866 22930
rect 18510 22878 18562 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 19630 22542 19682 22594
rect 21646 22542 21698 22594
rect 1934 22430 1986 22482
rect 21758 22430 21810 22482
rect 28590 22430 28642 22482
rect 40014 22430 40066 22482
rect 4286 22318 4338 22370
rect 14366 22318 14418 22370
rect 18734 22318 18786 22370
rect 19854 22318 19906 22370
rect 20190 22318 20242 22370
rect 21982 22318 22034 22370
rect 25790 22318 25842 22370
rect 37662 22318 37714 22370
rect 14030 22206 14082 22258
rect 14142 22206 14194 22258
rect 14702 22206 14754 22258
rect 17838 22206 17890 22258
rect 19294 22206 19346 22258
rect 23550 22206 23602 22258
rect 26462 22206 26514 22258
rect 18174 22094 18226 22146
rect 18510 22094 18562 22146
rect 19518 22094 19570 22146
rect 20078 22094 20130 22146
rect 23662 22094 23714 22146
rect 23886 22094 23938 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 15038 21758 15090 21810
rect 18846 21758 18898 21810
rect 25566 21758 25618 21810
rect 26462 21758 26514 21810
rect 14814 21646 14866 21698
rect 15486 21646 15538 21698
rect 15598 21646 15650 21698
rect 18398 21646 18450 21698
rect 26686 21646 26738 21698
rect 27806 21646 27858 21698
rect 14254 21534 14306 21586
rect 14478 21534 14530 21586
rect 15262 21534 15314 21586
rect 17614 21534 17666 21586
rect 18286 21534 18338 21586
rect 19070 21534 19122 21586
rect 19406 21534 19458 21586
rect 25230 21534 25282 21586
rect 25902 21534 25954 21586
rect 26462 21534 26514 21586
rect 27694 21534 27746 21586
rect 37886 21534 37938 21586
rect 11342 21422 11394 21474
rect 13470 21422 13522 21474
rect 22878 21422 22930 21474
rect 39902 21422 39954 21474
rect 14702 21310 14754 21362
rect 26126 21310 26178 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 14926 20974 14978 21026
rect 21198 20974 21250 21026
rect 40014 20862 40066 20914
rect 14030 20750 14082 20802
rect 14366 20750 14418 20802
rect 15150 20750 15202 20802
rect 20078 20750 20130 20802
rect 22206 20750 22258 20802
rect 22878 20750 22930 20802
rect 37998 20750 38050 20802
rect 14142 20638 14194 20690
rect 15710 20638 15762 20690
rect 21534 20638 21586 20690
rect 21758 20638 21810 20690
rect 22430 20638 22482 20690
rect 25790 20638 25842 20690
rect 14590 20526 14642 20578
rect 21310 20526 21362 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 22206 20190 22258 20242
rect 13246 20078 13298 20130
rect 13582 20078 13634 20130
rect 17502 20078 17554 20130
rect 18958 20078 19010 20130
rect 21646 20078 21698 20130
rect 22094 20078 22146 20130
rect 23998 20078 24050 20130
rect 24222 20078 24274 20130
rect 25566 20078 25618 20130
rect 25678 20078 25730 20130
rect 26462 20078 26514 20130
rect 27246 20078 27298 20130
rect 27358 20078 27410 20130
rect 29262 20078 29314 20130
rect 17838 19966 17890 20018
rect 18510 19966 18562 20018
rect 18846 19966 18898 20018
rect 19742 19966 19794 20018
rect 20526 19966 20578 20018
rect 20750 19966 20802 20018
rect 21310 19966 21362 20018
rect 21870 19966 21922 20018
rect 23774 19966 23826 20018
rect 24446 19966 24498 20018
rect 25342 19966 25394 20018
rect 26686 19966 26738 20018
rect 27022 19966 27074 20018
rect 29598 19966 29650 20018
rect 37662 19966 37714 20018
rect 18398 19854 18450 19906
rect 19518 19854 19570 19906
rect 26462 19854 26514 19906
rect 18174 19742 18226 19794
rect 24334 19742 24386 19794
rect 27358 19742 27410 19794
rect 40014 19742 40066 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 17726 19406 17778 19458
rect 19518 19406 19570 19458
rect 20638 19406 20690 19458
rect 20078 19294 20130 19346
rect 24110 19294 24162 19346
rect 26238 19294 26290 19346
rect 40014 19294 40066 19346
rect 15822 19182 15874 19234
rect 16606 19182 16658 19234
rect 17054 19182 17106 19234
rect 17502 19182 17554 19234
rect 18510 19182 18562 19234
rect 19966 19182 20018 19234
rect 23326 19182 23378 19234
rect 27470 19182 27522 19234
rect 29262 19182 29314 19234
rect 29934 19182 29986 19234
rect 37662 19182 37714 19234
rect 14926 19070 14978 19122
rect 20526 19070 20578 19122
rect 21310 19070 21362 19122
rect 21422 19070 21474 19122
rect 29486 19070 29538 19122
rect 15262 18958 15314 19010
rect 15598 18958 15650 19010
rect 16270 18958 16322 19010
rect 18734 18958 18786 19010
rect 20638 18958 20690 19010
rect 21646 18958 21698 19010
rect 27582 18958 27634 19010
rect 27806 18958 27858 19010
rect 30158 18958 30210 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 15710 18622 15762 18674
rect 16270 18622 16322 18674
rect 12686 18510 12738 18562
rect 17614 18510 17666 18562
rect 18398 18510 18450 18562
rect 26462 18510 26514 18562
rect 29374 18510 29426 18562
rect 4286 18398 4338 18450
rect 12014 18398 12066 18450
rect 15150 18398 15202 18450
rect 15486 18398 15538 18450
rect 17838 18398 17890 18450
rect 19518 18398 19570 18450
rect 21086 18398 21138 18450
rect 21310 18398 21362 18450
rect 22094 18398 22146 18450
rect 25678 18398 25730 18450
rect 29150 18398 29202 18450
rect 37662 18398 37714 18450
rect 14814 18286 14866 18338
rect 15598 18286 15650 18338
rect 16382 18286 16434 18338
rect 16718 18286 16770 18338
rect 17726 18286 17778 18338
rect 18510 18286 18562 18338
rect 20750 18286 20802 18338
rect 21982 18286 22034 18338
rect 28590 18286 28642 18338
rect 1934 18174 1986 18226
rect 16830 18174 16882 18226
rect 18174 18174 18226 18226
rect 19406 18174 19458 18226
rect 20638 18174 20690 18226
rect 22318 18174 22370 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 14254 17838 14306 17890
rect 16270 17838 16322 17890
rect 20414 17838 20466 17890
rect 23774 17838 23826 17890
rect 24110 17838 24162 17890
rect 9998 17726 10050 17778
rect 12126 17726 12178 17778
rect 14030 17726 14082 17778
rect 40014 17726 40066 17778
rect 12798 17614 12850 17666
rect 13582 17614 13634 17666
rect 13918 17614 13970 17666
rect 15038 17614 15090 17666
rect 16494 17614 16546 17666
rect 16718 17614 16770 17666
rect 17278 17614 17330 17666
rect 17950 17614 18002 17666
rect 18622 17614 18674 17666
rect 19630 17614 19682 17666
rect 20414 17614 20466 17666
rect 21310 17614 21362 17666
rect 21534 17614 21586 17666
rect 21982 17614 22034 17666
rect 23774 17614 23826 17666
rect 26462 17614 26514 17666
rect 26686 17614 26738 17666
rect 27134 17614 27186 17666
rect 27694 17614 27746 17666
rect 37886 17614 37938 17666
rect 16158 17502 16210 17554
rect 17614 17502 17666 17554
rect 18286 17502 18338 17554
rect 18958 17502 19010 17554
rect 19406 17502 19458 17554
rect 20078 17502 20130 17554
rect 20526 17502 20578 17554
rect 20862 17502 20914 17554
rect 21422 17502 21474 17554
rect 26574 17502 26626 17554
rect 27470 17390 27522 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 17502 17054 17554 17106
rect 18062 17054 18114 17106
rect 20302 17054 20354 17106
rect 20526 17054 20578 17106
rect 23774 17054 23826 17106
rect 14366 16942 14418 16994
rect 23438 16942 23490 16994
rect 23886 16942 23938 16994
rect 25230 16942 25282 16994
rect 25566 16942 25618 16994
rect 27134 16942 27186 16994
rect 13582 16830 13634 16882
rect 18398 16830 18450 16882
rect 18622 16830 18674 16882
rect 20190 16830 20242 16882
rect 21646 16830 21698 16882
rect 22094 16830 22146 16882
rect 22430 16830 22482 16882
rect 23102 16830 23154 16882
rect 23662 16830 23714 16882
rect 23998 16830 24050 16882
rect 26350 16830 26402 16882
rect 37662 16830 37714 16882
rect 16494 16718 16546 16770
rect 21982 16718 22034 16770
rect 22878 16718 22930 16770
rect 29262 16718 29314 16770
rect 22766 16606 22818 16658
rect 40014 16606 40066 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 20526 16270 20578 16322
rect 28254 16270 28306 16322
rect 23886 16158 23938 16210
rect 26014 16158 26066 16210
rect 28366 16158 28418 16210
rect 19406 16046 19458 16098
rect 19630 16046 19682 16098
rect 22094 16046 22146 16098
rect 22654 16046 22706 16098
rect 23102 16046 23154 16098
rect 20414 15934 20466 15986
rect 22542 15934 22594 15986
rect 19966 15822 20018 15874
rect 22430 15822 22482 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 18846 15486 18898 15538
rect 20078 15374 20130 15426
rect 20750 15374 20802 15426
rect 20862 15374 20914 15426
rect 22542 15374 22594 15426
rect 18510 15262 18562 15314
rect 19182 15262 19234 15314
rect 19406 15262 19458 15314
rect 20302 15262 20354 15314
rect 21870 15262 21922 15314
rect 18062 15150 18114 15202
rect 24670 15150 24722 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 16830 14590 16882 14642
rect 18958 14590 19010 14642
rect 19630 14590 19682 14642
rect 16158 14478 16210 14530
rect 19966 14478 20018 14530
rect 21310 14478 21362 14530
rect 19294 14366 19346 14418
rect 21646 14366 21698 14418
rect 20750 14254 20802 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 16830 13918 16882 13970
rect 17838 13694 17890 13746
rect 18510 13582 18562 13634
rect 20638 13582 20690 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 18846 12910 18898 12962
rect 18510 12798 18562 12850
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 25230 4286 25282 4338
rect 26238 4062 26290 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 25566 3614 25618 3666
rect 24558 3502 24610 3554
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 16800 41200 16912 42000
rect 17472 41200 17584 42000
rect 18816 41200 18928 42000
rect 20160 41200 20272 42000
rect 21504 41200 21616 42000
rect 22176 41200 22288 42000
rect 23520 41200 23632 42000
rect 24864 41200 24976 42000
rect 26208 41200 26320 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 16828 36708 16884 41200
rect 17500 38276 17556 41200
rect 17500 38210 17556 38220
rect 18620 38276 18676 38286
rect 18620 38182 18676 38220
rect 16828 36642 16884 36652
rect 17724 38050 17780 38062
rect 17724 37998 17726 38050
rect 17778 37998 17780 38050
rect 17276 36482 17332 36494
rect 17276 36430 17278 36482
rect 17330 36430 17332 36482
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 16156 27746 16212 27758
rect 16156 27694 16158 27746
rect 16210 27694 16212 27746
rect 4172 27636 4228 27646
rect 1932 25618 1988 25630
rect 1932 25566 1934 25618
rect 1986 25566 1988 25618
rect 1932 24948 1988 25566
rect 1932 24882 1988 24892
rect 1932 24500 1988 24510
rect 1932 24406 1988 24444
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 1932 23538 1988 23548
rect 1932 22932 1988 22942
rect 1932 22838 1988 22876
rect 1932 22482 1988 22494
rect 1932 22430 1934 22482
rect 1986 22430 1988 22482
rect 1932 21588 1988 22430
rect 1932 21522 1988 21532
rect 4172 21476 4228 27580
rect 14700 27636 14756 27646
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 14700 26402 14756 27580
rect 16044 27636 16100 27646
rect 16044 27542 16100 27580
rect 15708 27074 15764 27086
rect 15708 27022 15710 27074
rect 15762 27022 15764 27074
rect 15708 26964 15764 27022
rect 15708 26898 15764 26908
rect 14700 26350 14702 26402
rect 14754 26350 14756 26402
rect 14700 26338 14756 26350
rect 14028 26292 14084 26302
rect 14028 26290 14308 26292
rect 14028 26238 14030 26290
rect 14082 26238 14308 26290
rect 14028 26236 14308 26238
rect 14028 26226 14084 26236
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4284 25508 4340 25518
rect 4284 25414 4340 25452
rect 4284 24724 4340 24734
rect 4284 24630 4340 24668
rect 12236 24610 12292 24622
rect 12236 24558 12238 24610
rect 12290 24558 12292 24610
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4284 23940 4340 23950
rect 4284 23846 4340 23884
rect 12236 23940 12292 24558
rect 12236 23874 12292 23884
rect 4284 23156 4340 23166
rect 4284 23062 4340 23100
rect 11452 23156 11508 23166
rect 11452 23042 11508 23100
rect 14140 23156 14196 23166
rect 11452 22990 11454 23042
rect 11506 22990 11508 23042
rect 11452 22978 11508 22990
rect 13580 23042 13636 23054
rect 13580 22990 13582 23042
rect 13634 22990 13636 23042
rect 13580 22932 13636 22990
rect 13692 22932 13748 22942
rect 13580 22876 13692 22932
rect 13692 22866 13748 22876
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4284 22370 4340 22382
rect 4284 22318 4286 22370
rect 4338 22318 4340 22370
rect 4284 21588 4340 22318
rect 14028 22258 14084 22270
rect 14028 22206 14030 22258
rect 14082 22206 14084 22258
rect 4284 21522 4340 21532
rect 11340 21588 11396 21598
rect 4172 21410 4228 21420
rect 11340 21474 11396 21532
rect 11340 21422 11342 21474
rect 11394 21422 11396 21474
rect 11340 21410 11396 21422
rect 13468 21474 13524 21486
rect 13468 21422 13470 21474
rect 13522 21422 13524 21474
rect 13468 21364 13524 21422
rect 13692 21364 13748 21374
rect 13468 21308 13692 21364
rect 13692 21298 13748 21308
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 14028 20804 14084 22206
rect 14140 22258 14196 23100
rect 14140 22206 14142 22258
rect 14194 22206 14196 22258
rect 14140 22194 14196 22206
rect 14252 23154 14308 26236
rect 16156 25620 16212 27694
rect 16380 27636 16436 27646
rect 16380 27186 16436 27580
rect 17276 27188 17332 36430
rect 17500 27748 17556 27758
rect 17500 27746 17668 27748
rect 17500 27694 17502 27746
rect 17554 27694 17668 27746
rect 17500 27692 17668 27694
rect 17500 27682 17556 27692
rect 17388 27636 17444 27646
rect 17388 27542 17444 27580
rect 16380 27134 16382 27186
rect 16434 27134 16436 27186
rect 16380 27122 16436 27134
rect 16828 27132 17332 27188
rect 16828 26178 16884 27132
rect 16828 26126 16830 26178
rect 16882 26126 16884 26178
rect 16828 26114 16884 26126
rect 16940 26964 16996 26974
rect 16156 25554 16212 25564
rect 15484 25508 15540 25518
rect 15484 24946 15540 25452
rect 15484 24894 15486 24946
rect 15538 24894 15540 24946
rect 15484 24882 15540 24894
rect 16940 25282 16996 26908
rect 17276 26908 17332 27132
rect 17276 26852 17444 26908
rect 17388 26516 17444 26852
rect 17388 26514 17556 26516
rect 17388 26462 17390 26514
rect 17442 26462 17556 26514
rect 17388 26460 17556 26462
rect 17388 26450 17444 26460
rect 17276 26292 17332 26302
rect 16940 25230 16942 25282
rect 16994 25230 16996 25282
rect 14812 24724 14868 24734
rect 14364 24610 14420 24622
rect 14364 24558 14366 24610
rect 14418 24558 14420 24610
rect 14364 24052 14420 24558
rect 14364 23986 14420 23996
rect 14812 23826 14868 24668
rect 15148 24722 15204 24734
rect 15148 24670 15150 24722
rect 15202 24670 15204 24722
rect 15148 24612 15204 24670
rect 15036 23940 15092 23950
rect 15036 23846 15092 23884
rect 14812 23774 14814 23826
rect 14866 23774 14868 23826
rect 14812 23762 14868 23774
rect 14812 23268 14868 23278
rect 14812 23266 14980 23268
rect 14812 23214 14814 23266
rect 14866 23214 14980 23266
rect 14812 23212 14980 23214
rect 14812 23202 14868 23212
rect 14252 23102 14254 23154
rect 14306 23102 14308 23154
rect 14252 22148 14308 23102
rect 14700 23154 14756 23166
rect 14700 23102 14702 23154
rect 14754 23102 14756 23154
rect 14700 22708 14756 23102
rect 14812 22932 14868 22942
rect 14812 22838 14868 22876
rect 14364 22652 14756 22708
rect 14364 22370 14420 22652
rect 14924 22596 14980 23212
rect 14924 22530 14980 22540
rect 15148 22484 15204 24556
rect 15708 24722 15764 24734
rect 15708 24670 15710 24722
rect 15762 24670 15764 24722
rect 15708 23940 15764 24670
rect 16268 24612 16324 24622
rect 16268 24518 16324 24556
rect 16940 24612 16996 25230
rect 16940 24546 16996 24556
rect 17164 25284 17220 25294
rect 17276 25284 17332 26236
rect 17388 25620 17444 25630
rect 17388 25526 17444 25564
rect 17500 25506 17556 26460
rect 17612 26068 17668 27692
rect 17724 26514 17780 37998
rect 18844 37492 18900 41200
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 18844 37426 18900 37436
rect 19852 37492 19908 37502
rect 19852 37398 19908 37436
rect 18844 37266 18900 37278
rect 18844 37214 18846 37266
rect 18898 37214 18900 37266
rect 18060 36708 18116 36718
rect 18060 36614 18116 36652
rect 18844 31948 18900 37214
rect 20188 36708 20244 41200
rect 20188 36642 20244 36652
rect 21420 38050 21476 38062
rect 21420 37998 21422 38050
rect 21474 37998 21476 38050
rect 21308 36484 21364 36494
rect 20300 36482 21364 36484
rect 20300 36430 21310 36482
rect 21362 36430 21364 36482
rect 20300 36428 21364 36430
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 18620 31892 18900 31948
rect 18508 27858 18564 27870
rect 18508 27806 18510 27858
rect 18562 27806 18564 27858
rect 18284 27748 18340 27758
rect 18508 27748 18564 27806
rect 18284 27746 18564 27748
rect 18284 27694 18286 27746
rect 18338 27694 18564 27746
rect 18284 27692 18564 27694
rect 18284 26964 18340 27692
rect 18508 27188 18564 27198
rect 18620 27188 18676 31892
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20188 28644 20244 28654
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20188 28084 20244 28588
rect 20076 28028 20244 28084
rect 19292 27748 19348 27758
rect 19292 27746 20020 27748
rect 19292 27694 19294 27746
rect 19346 27694 20020 27746
rect 19292 27692 20020 27694
rect 19292 27682 19348 27692
rect 18284 26898 18340 26908
rect 18396 27186 18676 27188
rect 18396 27134 18510 27186
rect 18562 27134 18676 27186
rect 18396 27132 18676 27134
rect 17724 26462 17726 26514
rect 17778 26462 17780 26514
rect 17724 26450 17780 26462
rect 18396 26514 18452 27132
rect 18508 27122 18564 27132
rect 19964 27074 20020 27692
rect 19964 27022 19966 27074
rect 20018 27022 20020 27074
rect 19964 27010 20020 27022
rect 18956 26964 19012 26974
rect 19628 26964 19684 26974
rect 18956 26870 19012 26908
rect 19068 26962 19684 26964
rect 19068 26910 19630 26962
rect 19682 26910 19684 26962
rect 19068 26908 19684 26910
rect 18396 26462 18398 26514
rect 18450 26462 18452 26514
rect 18396 26450 18452 26462
rect 18620 26852 18676 26862
rect 18620 26514 18676 26796
rect 18620 26462 18622 26514
rect 18674 26462 18676 26514
rect 18620 26450 18676 26462
rect 18172 26292 18228 26302
rect 18172 26198 18228 26236
rect 18732 26290 18788 26302
rect 18732 26238 18734 26290
rect 18786 26238 18788 26290
rect 18396 26178 18452 26190
rect 18396 26126 18398 26178
rect 18450 26126 18452 26178
rect 18396 26068 18452 26126
rect 17612 26012 18452 26068
rect 17500 25454 17502 25506
rect 17554 25454 17556 25506
rect 17500 25442 17556 25454
rect 17948 25396 18004 25406
rect 17948 25302 18004 25340
rect 18508 25394 18564 25406
rect 18508 25342 18510 25394
rect 18562 25342 18564 25394
rect 17388 25284 17444 25294
rect 17276 25282 17444 25284
rect 17276 25230 17390 25282
rect 17442 25230 17444 25282
rect 17276 25228 17444 25230
rect 17052 24052 17108 24062
rect 17052 23958 17108 23996
rect 15484 23826 15540 23838
rect 15484 23774 15486 23826
rect 15538 23774 15540 23826
rect 15372 23042 15428 23054
rect 15372 22990 15374 23042
rect 15426 22990 15428 23042
rect 15372 22484 15428 22990
rect 14364 22318 14366 22370
rect 14418 22318 14420 22370
rect 14364 22306 14420 22318
rect 15036 22428 15428 22484
rect 14700 22260 14756 22270
rect 15036 22260 15092 22428
rect 14588 22258 15092 22260
rect 14588 22206 14702 22258
rect 14754 22206 15092 22258
rect 14588 22204 15092 22206
rect 14588 22148 14644 22204
rect 14700 22194 14756 22204
rect 14252 22092 14644 22148
rect 14028 20710 14084 20748
rect 14140 21588 14196 21598
rect 14140 20690 14196 21532
rect 14140 20638 14142 20690
rect 14194 20638 14196 20690
rect 14140 20626 14196 20638
rect 14252 21586 14308 22092
rect 14924 22036 14980 22046
rect 15484 22036 15540 23774
rect 15596 23828 15652 23838
rect 15708 23828 15764 23884
rect 15820 23940 15876 23950
rect 16156 23940 16212 23950
rect 15820 23938 16212 23940
rect 15820 23886 15822 23938
rect 15874 23886 16158 23938
rect 16210 23886 16212 23938
rect 15820 23884 16212 23886
rect 15820 23874 15876 23884
rect 16156 23874 16212 23884
rect 16604 23938 16660 23950
rect 16604 23886 16606 23938
rect 16658 23886 16660 23938
rect 15596 23826 15764 23828
rect 15596 23774 15598 23826
rect 15650 23774 15764 23826
rect 15596 23772 15764 23774
rect 15596 23762 15652 23772
rect 16604 23380 16660 23886
rect 16716 23940 16772 23950
rect 16828 23940 16884 23950
rect 16716 23938 16828 23940
rect 16716 23886 16718 23938
rect 16770 23886 16828 23938
rect 16716 23884 16828 23886
rect 16716 23874 16772 23884
rect 16604 23314 16660 23324
rect 14980 21980 15092 22036
rect 14924 21970 14980 21980
rect 15036 21812 15092 21980
rect 15036 21718 15092 21756
rect 15372 21980 15484 22036
rect 14812 21700 14868 21710
rect 14812 21606 14868 21644
rect 14252 21534 14254 21586
rect 14306 21534 14308 21586
rect 14252 20692 14308 21534
rect 14476 21586 14532 21598
rect 14476 21534 14478 21586
rect 14530 21534 14532 21586
rect 14364 20804 14420 20814
rect 14476 20804 14532 21534
rect 15260 21586 15316 21598
rect 15260 21534 15262 21586
rect 15314 21534 15316 21586
rect 14700 21364 14756 21374
rect 14700 21270 14756 21308
rect 14924 21028 14980 21038
rect 15260 21028 15316 21534
rect 14924 21026 15316 21028
rect 14924 20974 14926 21026
rect 14978 20974 15316 21026
rect 14924 20972 15316 20974
rect 14924 20962 14980 20972
rect 15372 20916 15428 21980
rect 15484 21970 15540 21980
rect 15596 22148 15652 22158
rect 15148 20860 15428 20916
rect 15484 21698 15540 21710
rect 15484 21646 15486 21698
rect 15538 21646 15540 21698
rect 14364 20802 14532 20804
rect 14364 20750 14366 20802
rect 14418 20750 14532 20802
rect 14364 20748 14532 20750
rect 14924 20804 14980 20814
rect 14364 20738 14420 20748
rect 14252 20626 14308 20636
rect 14588 20580 14644 20590
rect 14364 20578 14644 20580
rect 14364 20526 14590 20578
rect 14642 20526 14644 20578
rect 14364 20524 14644 20526
rect 14364 20244 14420 20524
rect 14588 20514 14644 20524
rect 13580 20188 14420 20244
rect 13244 20132 13300 20142
rect 12684 20130 13300 20132
rect 12684 20078 13246 20130
rect 13298 20078 13300 20130
rect 12684 20076 13300 20078
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 12684 18562 12740 20076
rect 13244 20066 13300 20076
rect 13580 20130 13636 20188
rect 13580 20078 13582 20130
rect 13634 20078 13636 20130
rect 13580 20066 13636 20078
rect 12684 18510 12686 18562
rect 12738 18510 12740 18562
rect 12684 18498 12740 18510
rect 14924 19122 14980 20748
rect 15148 20802 15204 20860
rect 15148 20750 15150 20802
rect 15202 20750 15204 20802
rect 15148 20738 15204 20750
rect 15484 20804 15540 21646
rect 15596 21698 15652 22092
rect 15596 21646 15598 21698
rect 15650 21646 15652 21698
rect 15596 21634 15652 21646
rect 15484 20738 15540 20748
rect 15708 20692 15764 20702
rect 15708 20598 15764 20636
rect 16156 20132 16212 20142
rect 14924 19070 14926 19122
rect 14978 19070 14980 19122
rect 4284 18452 4340 18462
rect 4284 18358 4340 18396
rect 9996 18452 10052 18462
rect 1932 18228 1988 18238
rect 1932 18134 1988 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 9996 17778 10052 18396
rect 12012 18452 12068 18462
rect 12012 18358 12068 18396
rect 12796 18452 12852 18462
rect 14924 18452 14980 19070
rect 15820 19234 15876 19246
rect 15820 19182 15822 19234
rect 15874 19182 15876 19234
rect 15260 19012 15316 19022
rect 15596 19012 15652 19022
rect 15260 19010 15652 19012
rect 15260 18958 15262 19010
rect 15314 18958 15598 19010
rect 15650 18958 15652 19010
rect 15260 18956 15652 18958
rect 15260 18946 15316 18956
rect 15596 18564 15652 18956
rect 15708 19012 15764 19022
rect 15708 18674 15764 18956
rect 15708 18622 15710 18674
rect 15762 18622 15764 18674
rect 15708 18610 15764 18622
rect 15596 18498 15652 18508
rect 15148 18452 15204 18462
rect 14924 18450 15204 18452
rect 14924 18398 15150 18450
rect 15202 18398 15204 18450
rect 14924 18396 15204 18398
rect 9996 17726 9998 17778
rect 10050 17726 10052 17778
rect 9996 17714 10052 17726
rect 12124 17780 12180 17790
rect 12124 17686 12180 17724
rect 12796 17668 12852 18396
rect 15148 18386 15204 18396
rect 15484 18452 15540 18462
rect 15484 18358 15540 18396
rect 14252 18340 14308 18350
rect 13916 17892 13972 17902
rect 12796 17574 12852 17612
rect 13580 17668 13636 17678
rect 13580 16882 13636 17612
rect 13916 17666 13972 17836
rect 14252 17890 14308 18284
rect 14812 18338 14868 18350
rect 14812 18286 14814 18338
rect 14866 18286 14868 18338
rect 14812 18228 14868 18286
rect 15596 18340 15652 18350
rect 15596 18246 15652 18284
rect 14812 18162 14868 18172
rect 15820 18228 15876 19182
rect 15820 18162 15876 18172
rect 14252 17838 14254 17890
rect 14306 17838 14308 17890
rect 14252 17826 14308 17838
rect 16156 17892 16212 20076
rect 16716 20132 16772 20142
rect 16828 20132 16884 23884
rect 16940 23938 16996 23950
rect 16940 23886 16942 23938
rect 16994 23886 16996 23938
rect 16940 23156 16996 23886
rect 16940 23090 16996 23100
rect 17164 23826 17220 25228
rect 17388 24948 17444 25228
rect 17724 25284 17780 25294
rect 18508 25284 18564 25342
rect 18732 25396 18788 26238
rect 19068 26068 19124 26908
rect 19628 26898 19684 26908
rect 19740 26964 19796 26974
rect 19740 26962 19908 26964
rect 19740 26910 19742 26962
rect 19794 26910 19908 26962
rect 19740 26908 19908 26910
rect 20076 26908 20132 28028
rect 19740 26898 19796 26908
rect 19852 26852 20132 26908
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20188 26292 20244 26302
rect 19628 26180 19684 26190
rect 19628 26086 19684 26124
rect 18844 26012 19124 26068
rect 18844 25506 18900 26012
rect 18844 25454 18846 25506
rect 18898 25454 18900 25506
rect 18844 25442 18900 25454
rect 20188 25506 20244 26236
rect 20188 25454 20190 25506
rect 20242 25454 20244 25506
rect 20188 25442 20244 25454
rect 18732 25330 18788 25340
rect 19292 25396 19348 25406
rect 17724 25190 17780 25228
rect 18172 25228 18564 25284
rect 18620 25284 18676 25294
rect 17388 24892 17668 24948
rect 17500 24612 17556 24622
rect 17500 23938 17556 24556
rect 17500 23886 17502 23938
rect 17554 23886 17556 23938
rect 17500 23874 17556 23886
rect 17164 23774 17166 23826
rect 17218 23774 17220 23826
rect 17164 22148 17220 23774
rect 17388 23380 17444 23390
rect 17388 23286 17444 23324
rect 17500 23266 17556 23278
rect 17500 23214 17502 23266
rect 17554 23214 17556 23266
rect 17500 22372 17556 23214
rect 17500 22306 17556 22316
rect 17164 22082 17220 22092
rect 17612 22036 17668 24892
rect 17724 23154 17780 23166
rect 18060 23156 18116 23166
rect 18172 23156 18228 25228
rect 18620 25190 18676 25228
rect 18284 23826 18340 23838
rect 18284 23774 18286 23826
rect 18338 23774 18340 23826
rect 18284 23492 18340 23774
rect 18284 23426 18340 23436
rect 18956 23492 19012 23502
rect 18844 23380 18900 23390
rect 18732 23324 18844 23380
rect 18508 23268 18564 23278
rect 18508 23174 18564 23212
rect 17724 23102 17726 23154
rect 17778 23102 17780 23154
rect 17724 22260 17780 23102
rect 17724 22194 17780 22204
rect 17836 23100 18060 23156
rect 18116 23100 18228 23156
rect 18396 23154 18452 23166
rect 18396 23102 18398 23154
rect 18450 23102 18452 23154
rect 17836 22258 17892 23100
rect 18060 23062 18116 23100
rect 18396 22596 18452 23102
rect 18732 23044 18788 23324
rect 18844 23314 18900 23324
rect 18956 23378 19012 23436
rect 18956 23326 18958 23378
rect 19010 23326 19012 23378
rect 18956 23314 19012 23326
rect 18508 22988 18788 23044
rect 18956 23154 19012 23166
rect 18956 23102 18958 23154
rect 19010 23102 19012 23154
rect 18508 22930 18564 22988
rect 18508 22878 18510 22930
rect 18562 22878 18564 22930
rect 18508 22866 18564 22878
rect 18396 22540 18900 22596
rect 18732 22372 18788 22382
rect 17836 22206 17838 22258
rect 17890 22206 17892 22258
rect 17836 22194 17892 22206
rect 17948 22370 18788 22372
rect 17948 22318 18734 22370
rect 18786 22318 18788 22370
rect 17948 22316 18788 22318
rect 17612 21980 17780 22036
rect 17612 21588 17668 21598
rect 17612 21494 17668 21532
rect 17724 21476 17780 21980
rect 17836 21476 17892 21486
rect 17724 21420 17836 21476
rect 17836 21410 17892 21420
rect 17276 20692 17332 20702
rect 17332 20636 17444 20692
rect 17276 20626 17332 20636
rect 16772 20076 16884 20132
rect 16716 20066 16772 20076
rect 16604 19236 16660 19246
rect 17052 19236 17108 19246
rect 16380 19234 17108 19236
rect 16380 19182 16606 19234
rect 16658 19182 17054 19234
rect 17106 19182 17108 19234
rect 16380 19180 17108 19182
rect 16268 19012 16324 19022
rect 16268 18918 16324 18956
rect 16268 18676 16324 18686
rect 16380 18676 16436 19180
rect 16604 19170 16660 19180
rect 17052 19170 17108 19180
rect 16268 18674 16436 18676
rect 16268 18622 16270 18674
rect 16322 18622 16436 18674
rect 16268 18620 16436 18622
rect 16268 18610 16324 18620
rect 16716 18452 16772 18462
rect 16380 18338 16436 18350
rect 16380 18286 16382 18338
rect 16434 18286 16436 18338
rect 16268 17892 16324 17902
rect 16156 17890 16324 17892
rect 16156 17838 16270 17890
rect 16322 17838 16324 17890
rect 16156 17836 16324 17838
rect 16268 17826 16324 17836
rect 14028 17780 14084 17790
rect 14028 17686 14084 17724
rect 16380 17780 16436 18286
rect 16716 18338 16772 18396
rect 16716 18286 16718 18338
rect 16770 18286 16772 18338
rect 16492 18228 16548 18238
rect 16716 18228 16772 18286
rect 16548 18172 16772 18228
rect 16828 18228 16884 18238
rect 16492 18162 16548 18172
rect 16828 18134 16884 18172
rect 13916 17614 13918 17666
rect 13970 17614 13972 17666
rect 13916 17602 13972 17614
rect 15036 17668 15092 17678
rect 14364 17556 14420 17566
rect 14364 16994 14420 17500
rect 14364 16942 14366 16994
rect 14418 16942 14420 16994
rect 14364 16930 14420 16942
rect 13580 16830 13582 16882
rect 13634 16830 13636 16882
rect 13580 16818 13636 16830
rect 15036 16660 15092 17612
rect 16156 17556 16212 17566
rect 16156 17462 16212 17500
rect 16380 16772 16436 17724
rect 16716 17892 16772 17902
rect 16492 17668 16548 17678
rect 16492 17574 16548 17612
rect 16716 17666 16772 17836
rect 16716 17614 16718 17666
rect 16770 17614 16772 17666
rect 16716 17602 16772 17614
rect 17276 17780 17332 17790
rect 17276 17666 17332 17724
rect 17276 17614 17278 17666
rect 17330 17614 17332 17666
rect 17276 17602 17332 17614
rect 17388 17108 17444 20636
rect 17500 20132 17556 20142
rect 17500 20038 17556 20076
rect 17836 20020 17892 20030
rect 17836 19926 17892 19964
rect 17724 19460 17780 19470
rect 17724 19366 17780 19404
rect 17500 19234 17556 19246
rect 17500 19182 17502 19234
rect 17554 19182 17556 19234
rect 17500 18564 17556 19182
rect 17500 18498 17556 18508
rect 17612 18562 17668 18574
rect 17612 18510 17614 18562
rect 17666 18510 17668 18562
rect 17612 18340 17668 18510
rect 17836 18452 17892 18462
rect 17948 18452 18004 22316
rect 18172 22146 18228 22158
rect 18172 22094 18174 22146
rect 18226 22094 18228 22146
rect 18172 21588 18228 22094
rect 18396 21698 18452 22316
rect 18732 22306 18788 22316
rect 18508 22148 18564 22158
rect 18844 22148 18900 22540
rect 18508 22054 18564 22092
rect 18732 22092 18900 22148
rect 18396 21646 18398 21698
rect 18450 21646 18452 21698
rect 18396 21634 18452 21646
rect 18732 22036 18788 22092
rect 18284 21588 18340 21598
rect 18172 21586 18340 21588
rect 18172 21534 18286 21586
rect 18338 21534 18340 21586
rect 18172 21532 18340 21534
rect 18172 19794 18228 19806
rect 18172 19742 18174 19794
rect 18226 19742 18228 19794
rect 18172 19012 18228 19742
rect 18284 19460 18340 21532
rect 18396 21476 18452 21486
rect 18396 19906 18452 21420
rect 18508 20020 18564 20030
rect 18508 20018 18676 20020
rect 18508 19966 18510 20018
rect 18562 19966 18676 20018
rect 18508 19964 18676 19966
rect 18508 19954 18564 19964
rect 18396 19854 18398 19906
rect 18450 19854 18452 19906
rect 18396 19842 18452 19854
rect 18284 19394 18340 19404
rect 18172 18676 18228 18956
rect 18172 18610 18228 18620
rect 18508 19236 18564 19246
rect 18396 18562 18452 18574
rect 18396 18510 18398 18562
rect 18450 18510 18452 18562
rect 18396 18452 18452 18510
rect 17836 18450 18340 18452
rect 17836 18398 17838 18450
rect 17890 18398 18340 18450
rect 17836 18396 18340 18398
rect 17836 18386 17892 18396
rect 17612 17554 17668 18284
rect 17724 18338 17780 18350
rect 17724 18286 17726 18338
rect 17778 18286 17780 18338
rect 17724 17892 17780 18286
rect 17724 17826 17780 17836
rect 17948 18228 18004 18238
rect 17948 17666 18004 18172
rect 18172 18226 18228 18238
rect 18172 18174 18174 18226
rect 18226 18174 18228 18226
rect 18172 17780 18228 18174
rect 18284 18228 18340 18396
rect 18396 18386 18452 18396
rect 18508 18338 18564 19180
rect 18620 19124 18676 19964
rect 18732 19236 18788 21980
rect 18844 21812 18900 21822
rect 18956 21812 19012 23102
rect 18900 21756 19012 21812
rect 19180 23154 19236 23166
rect 19180 23102 19182 23154
rect 19234 23102 19236 23154
rect 18844 21718 18900 21756
rect 19068 21586 19124 21598
rect 19068 21534 19070 21586
rect 19122 21534 19124 21586
rect 18956 20130 19012 20142
rect 18956 20078 18958 20130
rect 19010 20078 19012 20130
rect 18844 20018 18900 20030
rect 18844 19966 18846 20018
rect 18898 19966 18900 20018
rect 18844 19460 18900 19966
rect 18844 19394 18900 19404
rect 18956 19796 19012 20078
rect 19068 20020 19124 21534
rect 19180 20692 19236 23102
rect 19292 22820 19348 25340
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20300 24052 20356 36428
rect 21308 36418 21364 36428
rect 21420 31948 21476 37998
rect 21532 37492 21588 41200
rect 22204 38276 22260 41200
rect 22428 38276 22484 38286
rect 22204 38274 22484 38276
rect 22204 38222 22430 38274
rect 22482 38222 22484 38274
rect 22204 38220 22484 38222
rect 22428 38210 22484 38220
rect 23548 38276 23604 41200
rect 23548 38210 23604 38220
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 21532 37426 21588 37436
rect 22764 37492 22820 37502
rect 22764 37398 22820 37436
rect 21084 31892 21476 31948
rect 21868 37266 21924 37278
rect 21868 37214 21870 37266
rect 21922 37214 21924 37266
rect 21084 26180 21140 31892
rect 21196 28644 21252 28654
rect 21196 28550 21252 28588
rect 21420 28532 21476 28542
rect 21420 27746 21476 28476
rect 21420 27694 21422 27746
rect 21474 27694 21476 27746
rect 21420 27682 21476 27694
rect 21532 28530 21588 28542
rect 21532 28478 21534 28530
rect 21586 28478 21588 28530
rect 21532 27188 21588 28478
rect 21868 28532 21924 37214
rect 22316 36708 22372 36718
rect 22316 36614 22372 36652
rect 24332 36260 24388 36270
rect 24556 36260 24612 37998
rect 24892 37492 24948 41200
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 26236 38276 26292 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 26236 38210 26292 38220
rect 29372 38276 29428 38286
rect 29372 38182 29428 38220
rect 28588 38050 28644 38062
rect 28588 37998 28590 38050
rect 28642 37998 28644 38050
rect 24892 37426 24948 37436
rect 26236 37492 26292 37502
rect 26236 37398 26292 37436
rect 24332 36258 24612 36260
rect 24332 36206 24334 36258
rect 24386 36206 24612 36258
rect 24332 36204 24612 36206
rect 25228 37266 25284 37278
rect 25228 37214 25230 37266
rect 25282 37214 25284 37266
rect 24332 31948 24388 36204
rect 21868 28466 21924 28476
rect 23884 31892 24388 31948
rect 21868 27860 21924 27870
rect 21868 27858 22484 27860
rect 21868 27806 21870 27858
rect 21922 27806 22484 27858
rect 21868 27804 22484 27806
rect 21868 27794 21924 27804
rect 20412 25396 20468 25406
rect 20412 25302 20468 25340
rect 21084 25284 21140 26124
rect 21196 27132 21532 27188
rect 21196 25396 21252 27132
rect 21532 27094 21588 27132
rect 21644 27076 21700 27086
rect 21644 26982 21700 27020
rect 21308 26962 21364 26974
rect 21868 26964 21924 26974
rect 21308 26910 21310 26962
rect 21362 26910 21364 26962
rect 21308 25732 21364 26910
rect 21756 26962 21924 26964
rect 21756 26910 21870 26962
rect 21922 26910 21924 26962
rect 21756 26908 21924 26910
rect 21420 26852 21476 26862
rect 21476 26796 21700 26852
rect 21420 26758 21476 26796
rect 21308 25676 21588 25732
rect 21196 25330 21252 25340
rect 21308 25394 21364 25406
rect 21308 25342 21310 25394
rect 21362 25342 21364 25394
rect 21084 25218 21140 25228
rect 20412 24052 20468 24062
rect 20300 24050 20468 24052
rect 20300 23998 20414 24050
rect 20466 23998 20468 24050
rect 20300 23996 20468 23998
rect 19628 23828 19684 23838
rect 19516 23380 19572 23390
rect 19404 23154 19460 23166
rect 19404 23102 19406 23154
rect 19458 23102 19460 23154
rect 19404 22932 19460 23102
rect 19516 23154 19572 23324
rect 19516 23102 19518 23154
rect 19570 23102 19572 23154
rect 19516 23090 19572 23102
rect 19628 22932 19684 23772
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20188 23380 20244 23390
rect 19964 23156 20020 23166
rect 19964 23062 20020 23100
rect 19404 22876 19684 22932
rect 19292 22764 19460 22820
rect 19180 20626 19236 20636
rect 19292 22260 19348 22270
rect 19068 19954 19124 19964
rect 19292 19796 19348 22204
rect 19404 21924 19460 22764
rect 19516 22372 19572 22876
rect 19628 22596 19684 22606
rect 20188 22596 20244 23324
rect 20300 23268 20356 23996
rect 20412 23986 20468 23996
rect 20412 23492 20468 23502
rect 20412 23378 20468 23436
rect 20412 23326 20414 23378
rect 20466 23326 20468 23378
rect 20412 23314 20468 23326
rect 21308 23380 21364 25342
rect 21532 25282 21588 25676
rect 21532 25230 21534 25282
rect 21586 25230 21588 25282
rect 21532 23940 21588 25230
rect 21532 23874 21588 23884
rect 21420 23714 21476 23726
rect 21420 23662 21422 23714
rect 21474 23662 21476 23714
rect 21420 23492 21476 23662
rect 21420 23426 21476 23436
rect 21308 23314 21364 23324
rect 21644 23268 21700 26796
rect 21756 26402 21812 26908
rect 21868 26898 21924 26908
rect 21980 26962 22036 26974
rect 21980 26910 21982 26962
rect 22034 26910 22036 26962
rect 21980 26516 22036 26910
rect 22428 26908 22484 27804
rect 22540 27748 22596 27758
rect 22540 27746 23156 27748
rect 22540 27694 22542 27746
rect 22594 27694 23156 27746
rect 22540 27692 23156 27694
rect 22540 27682 22596 27692
rect 23100 27298 23156 27692
rect 23100 27246 23102 27298
rect 23154 27246 23156 27298
rect 23100 27234 23156 27246
rect 22988 27076 23044 27086
rect 22988 26982 23044 27020
rect 23100 26964 23156 26974
rect 22428 26852 22596 26908
rect 23100 26870 23156 26908
rect 23772 26964 23828 26974
rect 23772 26870 23828 26908
rect 21756 26350 21758 26402
rect 21810 26350 21812 26402
rect 21756 26338 21812 26350
rect 21868 26460 22036 26516
rect 21868 26180 21924 26460
rect 21756 26124 21924 26180
rect 22540 26290 22596 26852
rect 22540 26238 22542 26290
rect 22594 26238 22596 26290
rect 21756 25618 21812 26124
rect 21756 25566 21758 25618
rect 21810 25566 21812 25618
rect 21756 25554 21812 25566
rect 22540 25508 22596 26238
rect 22540 25442 22596 25452
rect 23660 25508 23716 25518
rect 21756 25394 21812 25406
rect 21756 25342 21758 25394
rect 21810 25342 21812 25394
rect 21756 25284 21812 25342
rect 21868 25396 21924 25406
rect 21868 25302 21924 25340
rect 21756 25218 21812 25228
rect 20300 23202 20356 23212
rect 21532 23212 21700 23268
rect 20636 23156 20692 23166
rect 21084 23156 21140 23166
rect 20636 23154 21028 23156
rect 20636 23102 20638 23154
rect 20690 23102 21028 23154
rect 20636 23100 21028 23102
rect 20636 23090 20692 23100
rect 20524 23044 20580 23054
rect 20524 22950 20580 22988
rect 19628 22594 20244 22596
rect 19628 22542 19630 22594
rect 19682 22542 20244 22594
rect 19628 22540 20244 22542
rect 19628 22530 19684 22540
rect 19852 22372 19908 22382
rect 19516 22370 19908 22372
rect 19516 22318 19854 22370
rect 19906 22318 19908 22370
rect 19516 22316 19908 22318
rect 19852 22306 19908 22316
rect 20188 22370 20244 22540
rect 20188 22318 20190 22370
rect 20242 22318 20244 22370
rect 20188 22306 20244 22318
rect 19516 22148 19572 22158
rect 20076 22148 20132 22158
rect 19516 22054 19572 22092
rect 19628 22146 20132 22148
rect 19628 22094 20078 22146
rect 20130 22094 20132 22146
rect 19628 22092 20132 22094
rect 19628 21924 19684 22092
rect 20076 22082 20132 22092
rect 20300 22148 20356 22158
rect 19404 21868 19684 21924
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19404 21588 19460 21598
rect 19404 21494 19460 21532
rect 19628 21364 19684 21868
rect 18956 19740 19348 19796
rect 19404 21308 19684 21364
rect 18956 19348 19012 19740
rect 18956 19292 19124 19348
rect 18732 19180 18900 19236
rect 18620 19058 18676 19068
rect 18732 19012 18788 19022
rect 18732 18918 18788 18956
rect 18508 18286 18510 18338
rect 18562 18286 18564 18338
rect 18508 18274 18564 18286
rect 18620 18228 18676 18238
rect 18284 18172 18452 18228
rect 18172 17714 18228 17724
rect 17948 17614 17950 17666
rect 18002 17614 18004 17666
rect 17948 17602 18004 17614
rect 18060 17668 18116 17678
rect 17612 17502 17614 17554
rect 17666 17502 17668 17554
rect 17612 17490 17668 17502
rect 17500 17108 17556 17118
rect 17388 17106 17556 17108
rect 17388 17054 17502 17106
rect 17554 17054 17556 17106
rect 17388 17052 17556 17054
rect 16492 16772 16548 16782
rect 16380 16770 16548 16772
rect 16380 16718 16494 16770
rect 16546 16718 16548 16770
rect 16380 16716 16548 16718
rect 16492 16706 16548 16716
rect 15036 16604 15204 16660
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 15148 14308 15204 16604
rect 16828 15428 16884 15438
rect 16828 14642 16884 15372
rect 16828 14590 16830 14642
rect 16882 14590 16884 14642
rect 16828 14578 16884 14590
rect 15148 14242 15204 14252
rect 16156 14530 16212 14542
rect 16156 14478 16158 14530
rect 16210 14478 16212 14530
rect 16156 14308 16212 14478
rect 16156 14242 16212 14252
rect 16940 14308 16996 14318
rect 16828 13972 16884 13982
rect 16940 13972 16996 14252
rect 17500 14308 17556 17052
rect 18060 17106 18116 17612
rect 18284 17668 18340 17678
rect 18284 17554 18340 17612
rect 18284 17502 18286 17554
rect 18338 17502 18340 17554
rect 18284 17490 18340 17502
rect 18060 17054 18062 17106
rect 18114 17054 18116 17106
rect 18060 17042 18116 17054
rect 18396 16882 18452 18172
rect 18620 17666 18676 18172
rect 18844 18228 18900 19180
rect 18844 18162 18900 18172
rect 18956 19124 19012 19134
rect 18844 17780 18900 17790
rect 18620 17614 18622 17666
rect 18674 17614 18676 17666
rect 18620 17602 18676 17614
rect 18732 17724 18844 17780
rect 18396 16830 18398 16882
rect 18450 16830 18452 16882
rect 18396 16548 18452 16830
rect 18620 16884 18676 16894
rect 18732 16884 18788 17724
rect 18844 17714 18900 17724
rect 18956 17554 19012 19068
rect 18956 17502 18958 17554
rect 19010 17502 19012 17554
rect 18956 17490 19012 17502
rect 18620 16882 18788 16884
rect 18620 16830 18622 16882
rect 18674 16830 18788 16882
rect 18620 16828 18788 16830
rect 18620 16818 18676 16828
rect 18396 16492 18900 16548
rect 18844 15538 18900 16492
rect 18844 15486 18846 15538
rect 18898 15486 18900 15538
rect 18844 15474 18900 15486
rect 18508 15316 18564 15326
rect 18060 15204 18116 15242
rect 18508 15222 18564 15260
rect 18060 15138 18116 15148
rect 19068 15204 19124 19292
rect 19404 19012 19460 21308
rect 20076 20804 20132 20814
rect 20076 20710 20132 20748
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19740 20020 19796 20030
rect 19516 19908 19572 19918
rect 19516 19814 19572 19852
rect 19516 19460 19572 19470
rect 19740 19460 19796 19964
rect 20076 20020 20132 20030
rect 20076 19460 20132 19964
rect 19516 19458 19796 19460
rect 19516 19406 19518 19458
rect 19570 19406 19796 19458
rect 19516 19404 19796 19406
rect 19852 19404 20132 19460
rect 19516 19394 19572 19404
rect 19516 19012 19572 19022
rect 19852 19012 19908 19404
rect 20076 19346 20132 19404
rect 20076 19294 20078 19346
rect 20130 19294 20132 19346
rect 20076 19282 20132 19294
rect 19964 19234 20020 19246
rect 19964 19182 19966 19234
rect 20018 19182 20020 19234
rect 19964 19124 20020 19182
rect 19964 19058 20020 19068
rect 19404 18956 19516 19012
rect 19516 18946 19572 18956
rect 19628 18956 19908 19012
rect 19516 18450 19572 18462
rect 19516 18398 19518 18450
rect 19570 18398 19572 18450
rect 19404 18228 19460 18238
rect 19404 18134 19460 18172
rect 19404 17780 19460 17790
rect 19404 17554 19460 17724
rect 19516 17668 19572 18398
rect 19516 17602 19572 17612
rect 19628 18340 19684 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 17666 19684 18284
rect 19628 17614 19630 17666
rect 19682 17614 19684 17666
rect 19628 17602 19684 17614
rect 20076 18564 20132 18574
rect 19404 17502 19406 17554
rect 19458 17502 19460 17554
rect 19404 17490 19460 17502
rect 20076 17556 20132 18508
rect 20300 18116 20356 22092
rect 20972 20804 21028 23100
rect 21084 23062 21140 23100
rect 21196 21588 21252 21598
rect 21196 21026 21252 21532
rect 21532 21252 21588 23212
rect 23660 23156 23716 25452
rect 23660 23090 23716 23100
rect 23884 23492 23940 31892
rect 25228 28532 25284 37214
rect 24668 28476 25284 28532
rect 24668 27746 24724 28476
rect 24668 27694 24670 27746
rect 24722 27694 24724 27746
rect 24108 27188 24164 27198
rect 24108 27074 24164 27132
rect 24108 27022 24110 27074
rect 24162 27022 24164 27074
rect 24108 27010 24164 27022
rect 23996 26964 24052 26974
rect 23996 26870 24052 26908
rect 24668 26964 24724 27694
rect 25004 27188 25060 27198
rect 25060 27132 25172 27188
rect 25004 27122 25060 27132
rect 24668 26898 24724 26908
rect 25116 26908 25172 27132
rect 25116 26852 25284 26908
rect 25228 26402 25284 26852
rect 25340 26852 25396 26862
rect 25340 26514 25396 26796
rect 25340 26462 25342 26514
rect 25394 26462 25396 26514
rect 25340 26450 25396 26462
rect 26460 26852 26516 26862
rect 25228 26350 25230 26402
rect 25282 26350 25284 26402
rect 25228 26338 25284 26350
rect 24444 26068 24500 26078
rect 24332 25396 24388 25406
rect 24108 25394 24388 25396
rect 24108 25342 24334 25394
rect 24386 25342 24388 25394
rect 24108 25340 24388 25342
rect 24108 24946 24164 25340
rect 24332 25330 24388 25340
rect 24108 24894 24110 24946
rect 24162 24894 24164 24946
rect 24108 24882 24164 24894
rect 24332 24836 24388 24846
rect 21644 23044 21700 23054
rect 21644 22594 21700 22988
rect 21644 22542 21646 22594
rect 21698 22542 21700 22594
rect 21644 22530 21700 22542
rect 21756 23042 21812 23054
rect 21756 22990 21758 23042
rect 21810 22990 21812 23042
rect 21756 22482 21812 22990
rect 23884 23042 23940 23436
rect 23884 22990 23886 23042
rect 23938 22990 23940 23042
rect 23884 22978 23940 22990
rect 24220 24834 24388 24836
rect 24220 24782 24334 24834
rect 24386 24782 24388 24834
rect 24220 24780 24388 24782
rect 21756 22430 21758 22482
rect 21810 22430 21812 22482
rect 21756 22418 21812 22430
rect 21980 22370 22036 22382
rect 21980 22318 21982 22370
rect 22034 22318 22036 22370
rect 21980 22260 22036 22318
rect 22092 22260 22148 22270
rect 21980 22204 22092 22260
rect 22092 22194 22148 22204
rect 22316 22260 22372 22270
rect 22204 22148 22260 22158
rect 21532 21196 21700 21252
rect 21196 20974 21198 21026
rect 21250 20974 21252 21026
rect 21196 20962 21252 20974
rect 20972 20748 21476 20804
rect 21308 20578 21364 20590
rect 21308 20526 21310 20578
rect 21362 20526 21364 20578
rect 21308 20188 21364 20526
rect 20636 20132 21364 20188
rect 20524 20020 20580 20030
rect 20636 20020 20692 20132
rect 20300 18050 20356 18060
rect 20412 20018 20692 20020
rect 20412 19966 20526 20018
rect 20578 19966 20692 20018
rect 20412 19964 20692 19966
rect 20748 20018 20804 20030
rect 20748 19966 20750 20018
rect 20802 19966 20804 20018
rect 20412 17890 20468 19964
rect 20524 19954 20580 19964
rect 20636 19460 20692 19470
rect 20636 19366 20692 19404
rect 20748 19236 20804 19966
rect 21308 20020 21364 20030
rect 21420 20020 21476 20748
rect 21532 20692 21588 20702
rect 21532 20598 21588 20636
rect 21644 20132 21700 21196
rect 22204 20802 22260 22092
rect 22204 20750 22206 20802
rect 22258 20750 22260 20802
rect 21308 20018 21476 20020
rect 21308 19966 21310 20018
rect 21362 19966 21476 20018
rect 21308 19964 21476 19966
rect 21308 19954 21364 19964
rect 21420 19796 21476 19964
rect 21420 19730 21476 19740
rect 21532 20130 21700 20132
rect 21532 20078 21646 20130
rect 21698 20078 21700 20130
rect 21532 20076 21700 20078
rect 20748 19170 20804 19180
rect 20524 19122 20580 19134
rect 20524 19070 20526 19122
rect 20578 19070 20580 19122
rect 20524 19012 20580 19070
rect 21308 19122 21364 19134
rect 21308 19070 21310 19122
rect 21362 19070 21364 19122
rect 20524 18946 20580 18956
rect 20636 19012 20692 19022
rect 20636 19010 20804 19012
rect 20636 18958 20638 19010
rect 20690 18958 20804 19010
rect 20636 18956 20804 18958
rect 20636 18946 20692 18956
rect 20412 17838 20414 17890
rect 20466 17838 20468 17890
rect 20412 17826 20468 17838
rect 20636 18676 20692 18686
rect 20636 18226 20692 18620
rect 20748 18564 20804 18956
rect 21308 18788 21364 19070
rect 21420 19124 21476 19134
rect 21420 19030 21476 19068
rect 21308 18732 21476 18788
rect 20748 18498 20804 18508
rect 21084 18450 21140 18462
rect 21308 18452 21364 18462
rect 21084 18398 21086 18450
rect 21138 18398 21140 18450
rect 20748 18340 20804 18350
rect 20748 18246 20804 18284
rect 20636 18174 20638 18226
rect 20690 18174 20692 18226
rect 20412 17666 20468 17678
rect 20412 17614 20414 17666
rect 20466 17614 20468 17666
rect 20076 17554 20244 17556
rect 20076 17502 20078 17554
rect 20130 17502 20244 17554
rect 20076 17500 20244 17502
rect 20076 17490 20132 17500
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19964 17108 20020 17118
rect 20188 17108 20244 17500
rect 20300 17108 20356 17118
rect 20188 17106 20356 17108
rect 20188 17054 20302 17106
rect 20354 17054 20356 17106
rect 20188 17052 20356 17054
rect 19404 16100 19460 16110
rect 19292 16098 19460 16100
rect 19292 16046 19406 16098
rect 19458 16046 19460 16098
rect 19292 16044 19460 16046
rect 19180 15316 19236 15326
rect 19292 15316 19348 16044
rect 19404 16034 19460 16044
rect 19628 16098 19684 16110
rect 19628 16046 19630 16098
rect 19682 16046 19684 16098
rect 19236 15260 19348 15316
rect 19404 15316 19460 15326
rect 19628 15316 19684 16046
rect 19964 15874 20020 17052
rect 20300 17042 20356 17052
rect 20188 16884 20244 16894
rect 20188 16790 20244 16828
rect 20412 16212 20468 17614
rect 20524 17554 20580 17566
rect 20524 17502 20526 17554
rect 20578 17502 20580 17554
rect 20524 17106 20580 17502
rect 20524 17054 20526 17106
rect 20578 17054 20580 17106
rect 20524 17042 20580 17054
rect 20636 16996 20692 18174
rect 20636 16930 20692 16940
rect 20748 18116 20804 18126
rect 21084 18116 21140 18398
rect 20804 18060 21140 18116
rect 21196 18450 21364 18452
rect 21196 18398 21310 18450
rect 21362 18398 21364 18450
rect 21196 18396 21364 18398
rect 20524 16884 20580 16894
rect 20524 16322 20580 16828
rect 20524 16270 20526 16322
rect 20578 16270 20580 16322
rect 20524 16258 20580 16270
rect 19964 15822 19966 15874
rect 20018 15822 20020 15874
rect 19964 15810 20020 15822
rect 20300 16156 20468 16212
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19404 15314 19684 15316
rect 19404 15262 19406 15314
rect 19458 15262 19684 15314
rect 19404 15260 19684 15262
rect 20076 15426 20132 15438
rect 20076 15374 20078 15426
rect 20130 15374 20132 15426
rect 20076 15316 20132 15374
rect 19180 15222 19236 15260
rect 19404 15250 19460 15260
rect 19068 15138 19124 15148
rect 18956 14644 19012 14654
rect 18956 14550 19012 14588
rect 19516 14644 19572 15260
rect 20076 15250 20132 15260
rect 20300 15314 20356 16156
rect 20300 15262 20302 15314
rect 20354 15262 20356 15314
rect 19740 15204 19796 15214
rect 19516 14578 19572 14588
rect 19628 15092 19796 15148
rect 20300 15148 20356 15262
rect 20412 15986 20468 15998
rect 20412 15934 20414 15986
rect 20466 15934 20468 15986
rect 20412 15316 20468 15934
rect 20748 15428 20804 18060
rect 20860 17556 20916 17566
rect 21196 17556 21252 18396
rect 21308 18386 21364 18396
rect 21308 17892 21364 17902
rect 21308 17666 21364 17836
rect 21420 17780 21476 18732
rect 21420 17714 21476 17724
rect 21308 17614 21310 17666
rect 21362 17614 21364 17666
rect 21308 17602 21364 17614
rect 21532 17666 21588 20076
rect 21644 20066 21700 20076
rect 21756 20690 21812 20702
rect 21756 20638 21758 20690
rect 21810 20638 21812 20690
rect 21756 20132 21812 20638
rect 22204 20242 22260 20750
rect 22204 20190 22206 20242
rect 22258 20190 22260 20242
rect 22204 20178 22260 20190
rect 21756 19460 21812 20076
rect 22092 20130 22148 20142
rect 22092 20078 22094 20130
rect 22146 20078 22148 20130
rect 21868 20020 21924 20030
rect 21868 19926 21924 19964
rect 21756 19394 21812 19404
rect 22092 19124 22148 20078
rect 22092 19058 22148 19068
rect 21644 19012 21700 19022
rect 21644 19010 21812 19012
rect 21644 18958 21646 19010
rect 21698 18958 21812 19010
rect 21644 18956 21812 18958
rect 21644 18946 21700 18956
rect 21532 17614 21534 17666
rect 21586 17614 21588 17666
rect 20860 17554 21252 17556
rect 20860 17502 20862 17554
rect 20914 17502 21252 17554
rect 20860 17500 21252 17502
rect 21420 17556 21476 17566
rect 20860 17490 20916 17500
rect 21420 17462 21476 17500
rect 21532 17108 21588 17614
rect 21532 17042 21588 17052
rect 21644 18564 21700 18574
rect 21644 16882 21700 18508
rect 21756 18452 21812 18956
rect 21756 18396 22036 18452
rect 21980 18338 22036 18396
rect 21980 18286 21982 18338
rect 22034 18286 22036 18338
rect 21980 18274 22036 18286
rect 22092 18450 22148 18462
rect 22092 18398 22094 18450
rect 22146 18398 22148 18450
rect 22092 18340 22148 18398
rect 21644 16830 21646 16882
rect 21698 16830 21700 16882
rect 20748 15334 20804 15372
rect 20860 15428 20916 15438
rect 21644 15428 21700 16830
rect 21868 17780 21924 17790
rect 21868 16772 21924 17724
rect 21980 17668 22036 17678
rect 21980 16996 22036 17612
rect 21980 16930 22036 16940
rect 22092 16884 22148 18284
rect 22316 18228 22372 22204
rect 23548 22258 23604 22270
rect 23548 22206 23550 22258
rect 23602 22206 23604 22258
rect 22876 21474 22932 21486
rect 22876 21422 22878 21474
rect 22930 21422 22932 21474
rect 22876 20804 22932 21422
rect 22876 20710 22932 20748
rect 22428 20692 22484 20702
rect 22428 20598 22484 20636
rect 23548 20132 23604 22206
rect 23660 22148 23716 22158
rect 23660 22054 23716 22092
rect 23884 22146 23940 22158
rect 23884 22094 23886 22146
rect 23938 22094 23940 22146
rect 23884 21588 23940 22094
rect 24220 21812 24276 24780
rect 24332 24770 24388 24780
rect 24444 24834 24500 26012
rect 25340 26068 25396 26078
rect 25340 25974 25396 26012
rect 26460 25618 26516 26796
rect 28588 26852 28644 37998
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 28588 26786 28644 26796
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 26460 25566 26462 25618
rect 26514 25566 26516 25618
rect 26460 25554 26516 25566
rect 24444 24782 24446 24834
rect 24498 24782 24500 24834
rect 24444 24770 24500 24782
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 25452 23996 25844 24052
rect 25452 23938 25508 23996
rect 25452 23886 25454 23938
rect 25506 23886 25508 23938
rect 25452 23874 25508 23886
rect 25788 23940 25844 23996
rect 26236 23940 26292 23950
rect 25788 23938 26292 23940
rect 25788 23886 26238 23938
rect 26290 23886 26292 23938
rect 25788 23884 26292 23886
rect 26236 23874 26292 23884
rect 25116 23828 25172 23838
rect 25116 23734 25172 23772
rect 25676 23828 25732 23838
rect 25676 23826 26180 23828
rect 25676 23774 25678 23826
rect 25730 23774 26180 23826
rect 25676 23772 26180 23774
rect 25676 23762 25732 23772
rect 25340 23716 25396 23726
rect 25340 23714 25620 23716
rect 25340 23662 25342 23714
rect 25394 23662 25620 23714
rect 25340 23660 25620 23662
rect 25340 23650 25396 23660
rect 25564 23380 25620 23660
rect 25564 23324 26068 23380
rect 26012 23266 26068 23324
rect 26012 23214 26014 23266
rect 26066 23214 26068 23266
rect 26012 23202 26068 23214
rect 25340 23156 25396 23166
rect 25340 22372 25396 23100
rect 25788 22372 25844 22382
rect 25340 22370 25844 22372
rect 25340 22318 25790 22370
rect 25842 22318 25844 22370
rect 25340 22316 25844 22318
rect 23884 21522 23940 21532
rect 23996 21756 24276 21812
rect 25564 21810 25620 21822
rect 25564 21758 25566 21810
rect 25618 21758 25620 21810
rect 23548 20066 23604 20076
rect 23996 20692 24052 21756
rect 25564 21700 25620 21758
rect 25676 21700 25732 21710
rect 25564 21644 25676 21700
rect 23996 20130 24052 20636
rect 25228 21586 25284 21598
rect 25228 21534 25230 21586
rect 25282 21534 25284 21586
rect 23996 20078 23998 20130
rect 24050 20078 24052 20130
rect 23996 20066 24052 20078
rect 24220 20132 24276 20142
rect 24220 20038 24276 20076
rect 23772 20018 23828 20030
rect 23772 19966 23774 20018
rect 23826 19966 23828 20018
rect 23772 19908 23828 19966
rect 24444 20020 24500 20030
rect 24444 19926 24500 19964
rect 23772 19842 23828 19852
rect 24332 19796 24388 19806
rect 24108 19794 24388 19796
rect 24108 19742 24334 19794
rect 24386 19742 24388 19794
rect 24108 19740 24388 19742
rect 24108 19346 24164 19740
rect 24332 19730 24388 19740
rect 24444 19796 24500 19806
rect 24108 19294 24110 19346
rect 24162 19294 24164 19346
rect 24108 19282 24164 19294
rect 22316 18134 22372 18172
rect 23324 19234 23380 19246
rect 23324 19182 23326 19234
rect 23378 19182 23380 19234
rect 23324 18564 23380 19182
rect 23100 16996 23156 17006
rect 22092 16790 22148 16828
rect 22428 16884 22484 16894
rect 22652 16884 22708 16894
rect 22428 16882 22652 16884
rect 22428 16830 22430 16882
rect 22482 16830 22652 16882
rect 22428 16828 22652 16830
rect 22428 16818 22484 16828
rect 21980 16772 22036 16782
rect 21868 16770 22036 16772
rect 21868 16718 21982 16770
rect 22034 16718 22036 16770
rect 21868 16716 22036 16718
rect 21980 16100 22036 16716
rect 22092 16100 22148 16110
rect 21980 16098 22148 16100
rect 21980 16046 22094 16098
rect 22146 16046 22148 16098
rect 21980 16044 22148 16046
rect 22092 16034 22148 16044
rect 22652 16098 22708 16828
rect 23100 16882 23156 16940
rect 23100 16830 23102 16882
rect 23154 16830 23156 16882
rect 23100 16818 23156 16830
rect 22876 16770 22932 16782
rect 22876 16718 22878 16770
rect 22930 16718 22932 16770
rect 22652 16046 22654 16098
rect 22706 16046 22708 16098
rect 22652 16034 22708 16046
rect 22764 16658 22820 16670
rect 22764 16606 22766 16658
rect 22818 16606 22820 16658
rect 22540 15988 22596 15998
rect 22540 15894 22596 15932
rect 22428 15874 22484 15886
rect 22428 15822 22430 15874
rect 22482 15822 22484 15874
rect 22428 15764 22484 15822
rect 22764 15764 22820 16606
rect 22428 15708 22820 15764
rect 22876 15652 22932 16718
rect 20860 15426 21700 15428
rect 20860 15374 20862 15426
rect 20914 15374 21700 15426
rect 20860 15372 21700 15374
rect 20860 15362 20916 15372
rect 20412 15250 20468 15260
rect 20300 15092 20692 15148
rect 19628 14642 19684 15092
rect 19628 14590 19630 14642
rect 19682 14590 19684 14642
rect 19628 14578 19684 14590
rect 19964 14532 20020 14542
rect 19964 14438 20020 14476
rect 19292 14420 19348 14430
rect 18844 14418 19348 14420
rect 18844 14366 19294 14418
rect 19346 14366 19348 14418
rect 18844 14364 19348 14366
rect 17500 14242 17556 14252
rect 17836 14308 17892 14318
rect 16828 13970 16996 13972
rect 16828 13918 16830 13970
rect 16882 13918 16996 13970
rect 16828 13916 16996 13918
rect 16828 13906 16884 13916
rect 17836 13746 17892 14252
rect 17836 13694 17838 13746
rect 17890 13694 17892 13746
rect 17836 13682 17892 13694
rect 18508 13634 18564 13646
rect 18508 13582 18510 13634
rect 18562 13582 18564 13634
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 18508 12850 18564 13582
rect 18844 12962 18900 14364
rect 19292 14354 19348 14364
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20636 13634 20692 15092
rect 21308 14644 21364 14654
rect 21308 14530 21364 14588
rect 21308 14478 21310 14530
rect 21362 14478 21364 14530
rect 21308 14466 21364 14478
rect 21644 14532 21700 15372
rect 22540 15596 22932 15652
rect 23100 16100 23156 16110
rect 23324 16100 23380 18508
rect 24108 18228 24164 18238
rect 23772 17892 23828 17902
rect 23548 17890 23828 17892
rect 23548 17838 23774 17890
rect 23826 17838 23828 17890
rect 23548 17836 23828 17838
rect 23436 16996 23492 17006
rect 23436 16902 23492 16940
rect 23548 16660 23604 17836
rect 23772 17826 23828 17836
rect 24108 17890 24164 18172
rect 24108 17838 24110 17890
rect 24162 17838 24164 17890
rect 24108 17826 24164 17838
rect 23772 17666 23828 17678
rect 23772 17614 23774 17666
rect 23826 17614 23828 17666
rect 23772 17106 23828 17614
rect 24444 17220 24500 19740
rect 25228 19796 25284 21534
rect 25564 20132 25620 20142
rect 25564 20038 25620 20076
rect 25676 20130 25732 21644
rect 25676 20078 25678 20130
rect 25730 20078 25732 20130
rect 25340 20020 25396 20030
rect 25340 19926 25396 19964
rect 25676 20020 25732 20078
rect 25676 19954 25732 19964
rect 25788 20690 25844 22316
rect 26124 22260 26180 23772
rect 26572 23826 26628 23838
rect 26572 23774 26574 23826
rect 26626 23774 26628 23826
rect 26460 23716 26516 23726
rect 26460 23622 26516 23660
rect 25900 21588 25956 21598
rect 25900 21494 25956 21532
rect 26124 21362 26180 22204
rect 26460 22258 26516 22270
rect 26460 22206 26462 22258
rect 26514 22206 26516 22258
rect 26460 21810 26516 22206
rect 26460 21758 26462 21810
rect 26514 21758 26516 21810
rect 26460 21746 26516 21758
rect 26572 21700 26628 23774
rect 28140 23716 28196 23726
rect 28140 23044 28196 23660
rect 37660 23156 37716 23166
rect 37660 23062 37716 23100
rect 28140 22950 28196 22988
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 27804 22484 27860 22494
rect 26684 21700 26740 21710
rect 26628 21698 26740 21700
rect 26628 21646 26686 21698
rect 26738 21646 26740 21698
rect 26628 21644 26740 21646
rect 26572 21606 26628 21644
rect 26684 21634 26740 21644
rect 27804 21698 27860 22428
rect 28588 22484 28644 22494
rect 28588 22390 28644 22428
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 37660 22372 37716 22382
rect 37660 22278 37716 22316
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 27804 21646 27806 21698
rect 27858 21646 27860 21698
rect 27804 21634 27860 21646
rect 26460 21588 26516 21598
rect 26460 21494 26516 21532
rect 27692 21588 27748 21598
rect 27692 21494 27748 21532
rect 37884 21586 37940 21598
rect 37884 21534 37886 21586
rect 37938 21534 37940 21586
rect 26124 21310 26126 21362
rect 26178 21310 26180 21362
rect 26124 21298 26180 21310
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 25788 20638 25790 20690
rect 25842 20638 25844 20690
rect 25228 19236 25284 19740
rect 25228 19170 25284 19180
rect 25676 18564 25732 18574
rect 25676 18452 25732 18508
rect 25788 18452 25844 20638
rect 26236 20132 26292 20142
rect 26460 20132 26516 20142
rect 26236 19796 26292 20076
rect 26236 19346 26292 19740
rect 26236 19294 26238 19346
rect 26290 19294 26292 19346
rect 26236 19282 26292 19294
rect 26348 20130 26516 20132
rect 26348 20078 26462 20130
rect 26514 20078 26516 20130
rect 26348 20076 26516 20078
rect 26348 19908 26404 20076
rect 26460 20066 26516 20076
rect 27244 20132 27300 20142
rect 27244 20038 27300 20076
rect 27356 20130 27412 20142
rect 27356 20078 27358 20130
rect 27410 20078 27412 20130
rect 26684 20020 26740 20030
rect 26572 20018 26740 20020
rect 26572 19966 26686 20018
rect 26738 19966 26740 20018
rect 26572 19964 26740 19966
rect 26348 18788 26404 19852
rect 26236 18732 26404 18788
rect 26460 19906 26516 19918
rect 26460 19854 26462 19906
rect 26514 19854 26516 19906
rect 25676 18450 26180 18452
rect 25676 18398 25678 18450
rect 25730 18398 26180 18450
rect 25676 18396 26180 18398
rect 25676 18386 25732 18396
rect 23772 17054 23774 17106
rect 23826 17054 23828 17106
rect 23772 17042 23828 17054
rect 24220 17164 24500 17220
rect 23884 16996 23940 17006
rect 23884 16902 23940 16940
rect 23660 16884 23716 16894
rect 23660 16790 23716 16828
rect 23996 16884 24052 16894
rect 24220 16884 24276 17164
rect 23996 16882 24276 16884
rect 23996 16830 23998 16882
rect 24050 16830 24276 16882
rect 23996 16828 24276 16830
rect 25228 16996 25284 17006
rect 23996 16818 24052 16828
rect 23548 16604 23940 16660
rect 23884 16210 23940 16604
rect 23884 16158 23886 16210
rect 23938 16158 23940 16210
rect 23884 16146 23940 16158
rect 23100 16098 23380 16100
rect 23100 16046 23102 16098
rect 23154 16046 23380 16098
rect 23100 16044 23380 16046
rect 22540 15426 22596 15596
rect 22540 15374 22542 15426
rect 22594 15374 22596 15426
rect 22540 15362 22596 15374
rect 21868 15316 21924 15326
rect 21868 15314 22484 15316
rect 21868 15262 21870 15314
rect 21922 15262 22484 15314
rect 21868 15260 22484 15262
rect 21868 15250 21924 15260
rect 22428 15204 22484 15260
rect 23100 15204 23156 16044
rect 22428 15148 23156 15204
rect 24668 15988 24724 15998
rect 24668 15202 24724 15932
rect 24668 15150 24670 15202
rect 24722 15150 24724 15202
rect 21644 14418 21700 14476
rect 21644 14366 21646 14418
rect 21698 14366 21700 14418
rect 21644 14354 21700 14366
rect 20748 14308 20804 14318
rect 20748 14214 20804 14252
rect 20636 13582 20638 13634
rect 20690 13582 20692 13634
rect 20636 13570 20692 13582
rect 18844 12910 18846 12962
rect 18898 12910 18900 12962
rect 18844 12898 18900 12910
rect 18508 12798 18510 12850
rect 18562 12798 18564 12850
rect 18508 12786 18564 12798
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 24668 8428 24724 15150
rect 24556 8372 24724 8428
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 24220 4116 24276 4126
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 23548 3668 23604 3678
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 23548 800 23604 3612
rect 24220 800 24276 4060
rect 24556 3554 24612 8372
rect 25228 4338 25284 16940
rect 25564 16994 25620 17006
rect 25564 16942 25566 16994
rect 25618 16942 25620 16994
rect 25564 16660 25620 16942
rect 25564 16594 25620 16604
rect 26012 16996 26068 17006
rect 26012 16210 26068 16940
rect 26124 16884 26180 18396
rect 26236 17668 26292 18732
rect 26460 18562 26516 19854
rect 26460 18510 26462 18562
rect 26514 18510 26516 18562
rect 26460 18498 26516 18510
rect 26460 17668 26516 17678
rect 26236 17666 26516 17668
rect 26236 17614 26462 17666
rect 26514 17614 26516 17666
rect 26236 17612 26516 17614
rect 26460 17602 26516 17612
rect 26572 17556 26628 19964
rect 26684 19954 26740 19964
rect 27020 20018 27076 20030
rect 27020 19966 27022 20018
rect 27074 19966 27076 20018
rect 27020 19796 27076 19966
rect 27356 20020 27412 20078
rect 27356 19954 27412 19964
rect 29260 20130 29316 20142
rect 29260 20078 29262 20130
rect 29314 20078 29316 20130
rect 29260 20020 29316 20078
rect 27356 19796 27412 19806
rect 27020 19794 27412 19796
rect 27020 19742 27358 19794
rect 27410 19742 27412 19794
rect 27020 19740 27412 19742
rect 27356 19730 27412 19740
rect 27468 19236 27524 19246
rect 29260 19236 29316 19964
rect 27468 19142 27524 19180
rect 29148 19180 29260 19236
rect 26684 19012 26740 19022
rect 26684 17666 26740 18956
rect 27580 19010 27636 19022
rect 27580 18958 27582 19010
rect 27634 18958 27636 19010
rect 27580 17892 27636 18958
rect 27804 19012 27860 19022
rect 27804 18918 27860 18956
rect 28588 18564 28644 18574
rect 28588 18338 28644 18508
rect 29148 18450 29204 19180
rect 29260 19142 29316 19180
rect 29596 20018 29652 20030
rect 37660 20020 37716 20030
rect 29596 19966 29598 20018
rect 29650 19966 29652 20018
rect 29484 19124 29540 19134
rect 29484 19030 29540 19068
rect 29148 18398 29150 18450
rect 29202 18398 29204 18450
rect 29148 18386 29204 18398
rect 29372 18562 29428 18574
rect 29372 18510 29374 18562
rect 29426 18510 29428 18562
rect 29372 18452 29428 18510
rect 29596 18564 29652 19966
rect 37548 20018 37716 20020
rect 37548 19966 37662 20018
rect 37714 19966 37716 20018
rect 37548 19964 37716 19966
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 29932 19236 29988 19246
rect 29932 19142 29988 19180
rect 30156 19012 30212 19022
rect 30156 18918 30212 18956
rect 37548 19012 37604 19964
rect 37660 19954 37716 19964
rect 37884 19796 37940 21534
rect 39900 21474 39956 21486
rect 39900 21422 39902 21474
rect 39954 21422 39956 21474
rect 39900 20916 39956 21422
rect 39900 20850 39956 20860
rect 40012 20914 40068 20926
rect 40012 20862 40014 20914
rect 40066 20862 40068 20914
rect 37884 19730 37940 19740
rect 37996 20802 38052 20814
rect 37996 20750 37998 20802
rect 38050 20750 38052 20802
rect 37548 18946 37604 18956
rect 37660 19234 37716 19246
rect 37660 19182 37662 19234
rect 37714 19182 37716 19234
rect 37660 18676 37716 19182
rect 37996 19124 38052 20750
rect 40012 20244 40068 20862
rect 40012 20178 40068 20188
rect 40012 19794 40068 19806
rect 40012 19742 40014 19794
rect 40066 19742 40068 19794
rect 40012 19572 40068 19742
rect 40012 19506 40068 19516
rect 37996 19058 38052 19068
rect 40012 19346 40068 19358
rect 40012 19294 40014 19346
rect 40066 19294 40068 19346
rect 40012 18900 40068 19294
rect 40012 18834 40068 18844
rect 37660 18610 37716 18620
rect 29596 18498 29652 18508
rect 29372 18386 29428 18396
rect 37660 18452 37716 18462
rect 37660 18358 37716 18396
rect 28588 18286 28590 18338
rect 28642 18286 28644 18338
rect 28588 18274 28644 18286
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 27580 17836 28308 17892
rect 26684 17614 26686 17666
rect 26738 17614 26740 17666
rect 26684 17602 26740 17614
rect 27132 17668 27188 17678
rect 27692 17668 27748 17678
rect 27132 17666 27748 17668
rect 27132 17614 27134 17666
rect 27186 17614 27694 17666
rect 27746 17614 27748 17666
rect 27132 17612 27748 17614
rect 27132 17602 27188 17612
rect 27692 17602 27748 17612
rect 26572 17462 26628 17500
rect 27468 17444 27524 17454
rect 27132 17442 27524 17444
rect 27132 17390 27470 17442
rect 27522 17390 27524 17442
rect 27132 17388 27524 17390
rect 27132 16994 27188 17388
rect 27468 17378 27524 17388
rect 27132 16942 27134 16994
rect 27186 16942 27188 16994
rect 27132 16930 27188 16942
rect 26348 16884 26404 16894
rect 26124 16882 26404 16884
rect 26124 16830 26350 16882
rect 26402 16830 26404 16882
rect 26124 16828 26404 16830
rect 26348 16818 26404 16828
rect 28252 16322 28308 17836
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 37884 17666 37940 17678
rect 37884 17614 37886 17666
rect 37938 17614 37940 17666
rect 37660 16882 37716 16894
rect 37660 16830 37662 16882
rect 37714 16830 37716 16882
rect 28252 16270 28254 16322
rect 28306 16270 28308 16322
rect 28252 16258 28308 16270
rect 28364 16772 28420 16782
rect 26012 16158 26014 16210
rect 26066 16158 26068 16210
rect 26012 16146 26068 16158
rect 28364 16210 28420 16716
rect 29260 16772 29316 16782
rect 29260 16678 29316 16716
rect 37660 16660 37716 16830
rect 37884 16772 37940 17614
rect 40012 16884 40068 17726
rect 40012 16818 40068 16828
rect 37884 16706 37940 16716
rect 37660 16594 37716 16604
rect 40012 16658 40068 16670
rect 40012 16606 40014 16658
rect 40066 16606 40068 16658
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 28364 16158 28366 16210
rect 28418 16158 28420 16210
rect 28364 16146 28420 16158
rect 40012 16212 40068 16606
rect 40012 16146 40068 16156
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 25228 4286 25230 4338
rect 25282 4286 25284 4338
rect 25228 4274 25284 4286
rect 26236 4116 26292 4126
rect 26236 4022 26292 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 23520 0 23632 800
rect 24192 0 24304 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 17500 38220 17556 38276
rect 18620 38274 18676 38276
rect 18620 38222 18622 38274
rect 18622 38222 18674 38274
rect 18674 38222 18676 38274
rect 18620 38220 18676 38222
rect 16828 36652 16884 36708
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4172 27580 4228 27636
rect 1932 24892 1988 24948
rect 1932 24498 1988 24500
rect 1932 24446 1934 24498
rect 1934 24446 1986 24498
rect 1986 24446 1988 24498
rect 1932 24444 1988 24446
rect 1932 23548 1988 23604
rect 1932 22930 1988 22932
rect 1932 22878 1934 22930
rect 1934 22878 1986 22930
rect 1986 22878 1988 22930
rect 1932 22876 1988 22878
rect 1932 21532 1988 21588
rect 14700 27580 14756 27636
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 16044 27634 16100 27636
rect 16044 27582 16046 27634
rect 16046 27582 16098 27634
rect 16098 27582 16100 27634
rect 16044 27580 16100 27582
rect 15708 26908 15764 26964
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4284 25506 4340 25508
rect 4284 25454 4286 25506
rect 4286 25454 4338 25506
rect 4338 25454 4340 25506
rect 4284 25452 4340 25454
rect 4284 24722 4340 24724
rect 4284 24670 4286 24722
rect 4286 24670 4338 24722
rect 4338 24670 4340 24722
rect 4284 24668 4340 24670
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4284 23938 4340 23940
rect 4284 23886 4286 23938
rect 4286 23886 4338 23938
rect 4338 23886 4340 23938
rect 4284 23884 4340 23886
rect 12236 23884 12292 23940
rect 4284 23154 4340 23156
rect 4284 23102 4286 23154
rect 4286 23102 4338 23154
rect 4338 23102 4340 23154
rect 4284 23100 4340 23102
rect 11452 23100 11508 23156
rect 14140 23100 14196 23156
rect 13692 22876 13748 22932
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4284 21532 4340 21588
rect 11340 21532 11396 21588
rect 4172 21420 4228 21476
rect 13692 21308 13748 21364
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 16380 27580 16436 27636
rect 17388 27634 17444 27636
rect 17388 27582 17390 27634
rect 17390 27582 17442 27634
rect 17442 27582 17444 27634
rect 17388 27580 17444 27582
rect 16940 26908 16996 26964
rect 16156 25564 16212 25620
rect 15484 25452 15540 25508
rect 17276 26236 17332 26292
rect 14812 24668 14868 24724
rect 14364 23996 14420 24052
rect 15148 24556 15204 24612
rect 15036 23938 15092 23940
rect 15036 23886 15038 23938
rect 15038 23886 15090 23938
rect 15090 23886 15092 23938
rect 15036 23884 15092 23886
rect 14812 22930 14868 22932
rect 14812 22878 14814 22930
rect 14814 22878 14866 22930
rect 14866 22878 14868 22930
rect 14812 22876 14868 22878
rect 14924 22540 14980 22596
rect 16268 24610 16324 24612
rect 16268 24558 16270 24610
rect 16270 24558 16322 24610
rect 16322 24558 16324 24610
rect 16268 24556 16324 24558
rect 16940 24556 16996 24612
rect 17164 25228 17220 25284
rect 17388 25618 17444 25620
rect 17388 25566 17390 25618
rect 17390 25566 17442 25618
rect 17442 25566 17444 25618
rect 17388 25564 17444 25566
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 18844 37436 18900 37492
rect 19852 37490 19908 37492
rect 19852 37438 19854 37490
rect 19854 37438 19906 37490
rect 19906 37438 19908 37490
rect 19852 37436 19908 37438
rect 18060 36706 18116 36708
rect 18060 36654 18062 36706
rect 18062 36654 18114 36706
rect 18114 36654 18116 36706
rect 18060 36652 18116 36654
rect 20188 36652 20244 36708
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 20188 28588 20244 28644
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 18284 26908 18340 26964
rect 18956 26962 19012 26964
rect 18956 26910 18958 26962
rect 18958 26910 19010 26962
rect 19010 26910 19012 26962
rect 18956 26908 19012 26910
rect 18620 26796 18676 26852
rect 18172 26290 18228 26292
rect 18172 26238 18174 26290
rect 18174 26238 18226 26290
rect 18226 26238 18228 26290
rect 18172 26236 18228 26238
rect 17948 25394 18004 25396
rect 17948 25342 17950 25394
rect 17950 25342 18002 25394
rect 18002 25342 18004 25394
rect 17948 25340 18004 25342
rect 17052 24050 17108 24052
rect 17052 23998 17054 24050
rect 17054 23998 17106 24050
rect 17106 23998 17108 24050
rect 17052 23996 17108 23998
rect 15708 23884 15764 23940
rect 14028 20802 14084 20804
rect 14028 20750 14030 20802
rect 14030 20750 14082 20802
rect 14082 20750 14084 20802
rect 14028 20748 14084 20750
rect 14140 21532 14196 21588
rect 16828 23884 16884 23940
rect 16604 23324 16660 23380
rect 14924 21980 14980 22036
rect 15036 21810 15092 21812
rect 15036 21758 15038 21810
rect 15038 21758 15090 21810
rect 15090 21758 15092 21810
rect 15036 21756 15092 21758
rect 15484 21980 15540 22036
rect 14812 21698 14868 21700
rect 14812 21646 14814 21698
rect 14814 21646 14866 21698
rect 14866 21646 14868 21698
rect 14812 21644 14868 21646
rect 14700 21362 14756 21364
rect 14700 21310 14702 21362
rect 14702 21310 14754 21362
rect 14754 21310 14756 21362
rect 14700 21308 14756 21310
rect 15596 22092 15652 22148
rect 14924 20748 14980 20804
rect 14252 20636 14308 20692
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 15484 20748 15540 20804
rect 15708 20690 15764 20692
rect 15708 20638 15710 20690
rect 15710 20638 15762 20690
rect 15762 20638 15764 20690
rect 15708 20636 15764 20638
rect 16156 20076 16212 20132
rect 4284 18450 4340 18452
rect 4284 18398 4286 18450
rect 4286 18398 4338 18450
rect 4338 18398 4340 18450
rect 4284 18396 4340 18398
rect 9996 18396 10052 18452
rect 1932 18226 1988 18228
rect 1932 18174 1934 18226
rect 1934 18174 1986 18226
rect 1986 18174 1988 18226
rect 1932 18172 1988 18174
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 12012 18450 12068 18452
rect 12012 18398 12014 18450
rect 12014 18398 12066 18450
rect 12066 18398 12068 18450
rect 12012 18396 12068 18398
rect 12796 18396 12852 18452
rect 15708 18956 15764 19012
rect 15596 18508 15652 18564
rect 12124 17778 12180 17780
rect 12124 17726 12126 17778
rect 12126 17726 12178 17778
rect 12178 17726 12180 17778
rect 12124 17724 12180 17726
rect 15484 18450 15540 18452
rect 15484 18398 15486 18450
rect 15486 18398 15538 18450
rect 15538 18398 15540 18450
rect 15484 18396 15540 18398
rect 14252 18284 14308 18340
rect 13916 17836 13972 17892
rect 12796 17666 12852 17668
rect 12796 17614 12798 17666
rect 12798 17614 12850 17666
rect 12850 17614 12852 17666
rect 12796 17612 12852 17614
rect 13580 17666 13636 17668
rect 13580 17614 13582 17666
rect 13582 17614 13634 17666
rect 13634 17614 13636 17666
rect 13580 17612 13636 17614
rect 15596 18338 15652 18340
rect 15596 18286 15598 18338
rect 15598 18286 15650 18338
rect 15650 18286 15652 18338
rect 15596 18284 15652 18286
rect 14812 18172 14868 18228
rect 15820 18172 15876 18228
rect 16940 23100 16996 23156
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20188 26236 20244 26292
rect 19628 26178 19684 26180
rect 19628 26126 19630 26178
rect 19630 26126 19682 26178
rect 19682 26126 19684 26178
rect 19628 26124 19684 26126
rect 18732 25340 18788 25396
rect 19292 25340 19348 25396
rect 17724 25282 17780 25284
rect 17724 25230 17726 25282
rect 17726 25230 17778 25282
rect 17778 25230 17780 25282
rect 17724 25228 17780 25230
rect 18620 25282 18676 25284
rect 18620 25230 18622 25282
rect 18622 25230 18674 25282
rect 18674 25230 18676 25282
rect 18620 25228 18676 25230
rect 17500 24610 17556 24612
rect 17500 24558 17502 24610
rect 17502 24558 17554 24610
rect 17554 24558 17556 24610
rect 17500 24556 17556 24558
rect 17388 23378 17444 23380
rect 17388 23326 17390 23378
rect 17390 23326 17442 23378
rect 17442 23326 17444 23378
rect 17388 23324 17444 23326
rect 17500 22316 17556 22372
rect 17164 22092 17220 22148
rect 18284 23436 18340 23492
rect 18956 23436 19012 23492
rect 18844 23324 18900 23380
rect 18508 23266 18564 23268
rect 18508 23214 18510 23266
rect 18510 23214 18562 23266
rect 18562 23214 18564 23266
rect 18508 23212 18564 23214
rect 17724 22204 17780 22260
rect 18060 23154 18116 23156
rect 18060 23102 18062 23154
rect 18062 23102 18114 23154
rect 18114 23102 18116 23154
rect 18060 23100 18116 23102
rect 17612 21586 17668 21588
rect 17612 21534 17614 21586
rect 17614 21534 17666 21586
rect 17666 21534 17668 21586
rect 17612 21532 17668 21534
rect 17836 21420 17892 21476
rect 17276 20636 17332 20692
rect 16716 20076 16772 20132
rect 16268 19010 16324 19012
rect 16268 18958 16270 19010
rect 16270 18958 16322 19010
rect 16322 18958 16324 19010
rect 16268 18956 16324 18958
rect 16716 18396 16772 18452
rect 14028 17778 14084 17780
rect 14028 17726 14030 17778
rect 14030 17726 14082 17778
rect 14082 17726 14084 17778
rect 14028 17724 14084 17726
rect 16492 18172 16548 18228
rect 16828 18226 16884 18228
rect 16828 18174 16830 18226
rect 16830 18174 16882 18226
rect 16882 18174 16884 18226
rect 16828 18172 16884 18174
rect 16380 17724 16436 17780
rect 15036 17666 15092 17668
rect 15036 17614 15038 17666
rect 15038 17614 15090 17666
rect 15090 17614 15092 17666
rect 15036 17612 15092 17614
rect 14364 17500 14420 17556
rect 16156 17554 16212 17556
rect 16156 17502 16158 17554
rect 16158 17502 16210 17554
rect 16210 17502 16212 17554
rect 16156 17500 16212 17502
rect 16716 17836 16772 17892
rect 16492 17666 16548 17668
rect 16492 17614 16494 17666
rect 16494 17614 16546 17666
rect 16546 17614 16548 17666
rect 16492 17612 16548 17614
rect 17276 17724 17332 17780
rect 17500 20130 17556 20132
rect 17500 20078 17502 20130
rect 17502 20078 17554 20130
rect 17554 20078 17556 20130
rect 17500 20076 17556 20078
rect 17836 20018 17892 20020
rect 17836 19966 17838 20018
rect 17838 19966 17890 20018
rect 17890 19966 17892 20018
rect 17836 19964 17892 19966
rect 17724 19458 17780 19460
rect 17724 19406 17726 19458
rect 17726 19406 17778 19458
rect 17778 19406 17780 19458
rect 17724 19404 17780 19406
rect 17500 18508 17556 18564
rect 18508 22146 18564 22148
rect 18508 22094 18510 22146
rect 18510 22094 18562 22146
rect 18562 22094 18564 22146
rect 18508 22092 18564 22094
rect 18732 21980 18788 22036
rect 18396 21420 18452 21476
rect 18284 19404 18340 19460
rect 18172 18956 18228 19012
rect 18172 18620 18228 18676
rect 18508 19234 18564 19236
rect 18508 19182 18510 19234
rect 18510 19182 18562 19234
rect 18562 19182 18564 19234
rect 18508 19180 18564 19182
rect 17612 18284 17668 18340
rect 17724 17836 17780 17892
rect 17948 18172 18004 18228
rect 18396 18396 18452 18452
rect 18844 21810 18900 21812
rect 18844 21758 18846 21810
rect 18846 21758 18898 21810
rect 18898 21758 18900 21810
rect 18844 21756 18900 21758
rect 18844 19404 18900 19460
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 23548 38220 23604 38276
rect 21532 37436 21588 37492
rect 22764 37490 22820 37492
rect 22764 37438 22766 37490
rect 22766 37438 22818 37490
rect 22818 37438 22820 37490
rect 22764 37436 22820 37438
rect 21196 28642 21252 28644
rect 21196 28590 21198 28642
rect 21198 28590 21250 28642
rect 21250 28590 21252 28642
rect 21196 28588 21252 28590
rect 21420 28530 21476 28532
rect 21420 28478 21422 28530
rect 21422 28478 21474 28530
rect 21474 28478 21476 28530
rect 21420 28476 21476 28478
rect 22316 36706 22372 36708
rect 22316 36654 22318 36706
rect 22318 36654 22370 36706
rect 22370 36654 22372 36706
rect 22316 36652 22372 36654
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 26236 38220 26292 38276
rect 29372 38274 29428 38276
rect 29372 38222 29374 38274
rect 29374 38222 29426 38274
rect 29426 38222 29428 38274
rect 29372 38220 29428 38222
rect 24892 37436 24948 37492
rect 26236 37490 26292 37492
rect 26236 37438 26238 37490
rect 26238 37438 26290 37490
rect 26290 37438 26292 37490
rect 26236 37436 26292 37438
rect 21868 28476 21924 28532
rect 21084 26124 21140 26180
rect 20412 25394 20468 25396
rect 20412 25342 20414 25394
rect 20414 25342 20466 25394
rect 20466 25342 20468 25394
rect 20412 25340 20468 25342
rect 21532 27132 21588 27188
rect 21644 27074 21700 27076
rect 21644 27022 21646 27074
rect 21646 27022 21698 27074
rect 21698 27022 21700 27074
rect 21644 27020 21700 27022
rect 21420 26850 21476 26852
rect 21420 26798 21422 26850
rect 21422 26798 21474 26850
rect 21474 26798 21476 26850
rect 21420 26796 21476 26798
rect 21196 25340 21252 25396
rect 21084 25228 21140 25284
rect 19628 23772 19684 23828
rect 19516 23324 19572 23380
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20188 23378 20244 23380
rect 20188 23326 20190 23378
rect 20190 23326 20242 23378
rect 20242 23326 20244 23378
rect 20188 23324 20244 23326
rect 19964 23154 20020 23156
rect 19964 23102 19966 23154
rect 19966 23102 20018 23154
rect 20018 23102 20020 23154
rect 19964 23100 20020 23102
rect 19180 20636 19236 20692
rect 19292 22258 19348 22260
rect 19292 22206 19294 22258
rect 19294 22206 19346 22258
rect 19346 22206 19348 22258
rect 19292 22204 19348 22206
rect 19068 19964 19124 20020
rect 20412 23436 20468 23492
rect 21532 23884 21588 23940
rect 21420 23436 21476 23492
rect 21308 23324 21364 23380
rect 22988 27074 23044 27076
rect 22988 27022 22990 27074
rect 22990 27022 23042 27074
rect 23042 27022 23044 27074
rect 22988 27020 23044 27022
rect 23100 26962 23156 26964
rect 23100 26910 23102 26962
rect 23102 26910 23154 26962
rect 23154 26910 23156 26962
rect 23100 26908 23156 26910
rect 23772 26962 23828 26964
rect 23772 26910 23774 26962
rect 23774 26910 23826 26962
rect 23826 26910 23828 26962
rect 23772 26908 23828 26910
rect 22540 25452 22596 25508
rect 23660 25506 23716 25508
rect 23660 25454 23662 25506
rect 23662 25454 23714 25506
rect 23714 25454 23716 25506
rect 23660 25452 23716 25454
rect 21868 25394 21924 25396
rect 21868 25342 21870 25394
rect 21870 25342 21922 25394
rect 21922 25342 21924 25394
rect 21868 25340 21924 25342
rect 21756 25228 21812 25284
rect 20300 23212 20356 23268
rect 20524 23042 20580 23044
rect 20524 22990 20526 23042
rect 20526 22990 20578 23042
rect 20578 22990 20580 23042
rect 20524 22988 20580 22990
rect 19516 22146 19572 22148
rect 19516 22094 19518 22146
rect 19518 22094 19570 22146
rect 19570 22094 19572 22146
rect 19516 22092 19572 22094
rect 20300 22092 20356 22148
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19404 21586 19460 21588
rect 19404 21534 19406 21586
rect 19406 21534 19458 21586
rect 19458 21534 19460 21586
rect 19404 21532 19460 21534
rect 18620 19068 18676 19124
rect 18732 19010 18788 19012
rect 18732 18958 18734 19010
rect 18734 18958 18786 19010
rect 18786 18958 18788 19010
rect 18732 18956 18788 18958
rect 18172 17724 18228 17780
rect 18060 17612 18116 17668
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 16828 15372 16884 15428
rect 15148 14252 15204 14308
rect 16156 14252 16212 14308
rect 16940 14252 16996 14308
rect 18284 17612 18340 17668
rect 18620 18172 18676 18228
rect 18844 18172 18900 18228
rect 18956 19068 19012 19124
rect 18844 17724 18900 17780
rect 18508 15314 18564 15316
rect 18508 15262 18510 15314
rect 18510 15262 18562 15314
rect 18562 15262 18564 15314
rect 18508 15260 18564 15262
rect 18060 15202 18116 15204
rect 18060 15150 18062 15202
rect 18062 15150 18114 15202
rect 18114 15150 18116 15202
rect 18060 15148 18116 15150
rect 20076 20802 20132 20804
rect 20076 20750 20078 20802
rect 20078 20750 20130 20802
rect 20130 20750 20132 20802
rect 20076 20748 20132 20750
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19740 20018 19796 20020
rect 19740 19966 19742 20018
rect 19742 19966 19794 20018
rect 19794 19966 19796 20018
rect 19740 19964 19796 19966
rect 19516 19906 19572 19908
rect 19516 19854 19518 19906
rect 19518 19854 19570 19906
rect 19570 19854 19572 19906
rect 19516 19852 19572 19854
rect 20076 19964 20132 20020
rect 19964 19068 20020 19124
rect 19516 18956 19572 19012
rect 19404 18226 19460 18228
rect 19404 18174 19406 18226
rect 19406 18174 19458 18226
rect 19458 18174 19460 18226
rect 19404 18172 19460 18174
rect 19404 17724 19460 17780
rect 19516 17612 19572 17668
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19628 18284 19684 18340
rect 20076 18508 20132 18564
rect 21084 23154 21140 23156
rect 21084 23102 21086 23154
rect 21086 23102 21138 23154
rect 21138 23102 21140 23154
rect 21084 23100 21140 23102
rect 21196 21532 21252 21588
rect 23660 23100 23716 23156
rect 24108 27132 24164 27188
rect 23996 26962 24052 26964
rect 23996 26910 23998 26962
rect 23998 26910 24050 26962
rect 24050 26910 24052 26962
rect 23996 26908 24052 26910
rect 25004 27132 25060 27188
rect 24668 26908 24724 26964
rect 25340 26796 25396 26852
rect 26460 26796 26516 26852
rect 24444 26012 24500 26068
rect 23884 23436 23940 23492
rect 21644 22988 21700 23044
rect 22092 22204 22148 22260
rect 22316 22204 22372 22260
rect 22204 22092 22260 22148
rect 20300 18060 20356 18116
rect 20636 19458 20692 19460
rect 20636 19406 20638 19458
rect 20638 19406 20690 19458
rect 20690 19406 20692 19458
rect 20636 19404 20692 19406
rect 21532 20690 21588 20692
rect 21532 20638 21534 20690
rect 21534 20638 21586 20690
rect 21586 20638 21588 20690
rect 21532 20636 21588 20638
rect 21420 19740 21476 19796
rect 20748 19180 20804 19236
rect 20524 18956 20580 19012
rect 20636 18620 20692 18676
rect 21420 19122 21476 19124
rect 21420 19070 21422 19122
rect 21422 19070 21474 19122
rect 21474 19070 21476 19122
rect 21420 19068 21476 19070
rect 20748 18508 20804 18564
rect 20748 18338 20804 18340
rect 20748 18286 20750 18338
rect 20750 18286 20802 18338
rect 20802 18286 20804 18338
rect 20748 18284 20804 18286
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19964 17052 20020 17108
rect 19180 15314 19236 15316
rect 19180 15262 19182 15314
rect 19182 15262 19234 15314
rect 19234 15262 19236 15314
rect 19180 15260 19236 15262
rect 20188 16882 20244 16884
rect 20188 16830 20190 16882
rect 20190 16830 20242 16882
rect 20242 16830 20244 16882
rect 20188 16828 20244 16830
rect 20636 16940 20692 16996
rect 20748 18060 20804 18116
rect 20524 16828 20580 16884
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20076 15260 20132 15316
rect 19068 15148 19124 15204
rect 18956 14642 19012 14644
rect 18956 14590 18958 14642
rect 18958 14590 19010 14642
rect 19010 14590 19012 14642
rect 18956 14588 19012 14590
rect 19740 15148 19796 15204
rect 19516 14588 19572 14644
rect 21308 17836 21364 17892
rect 21420 17724 21476 17780
rect 21756 20076 21812 20132
rect 21868 20018 21924 20020
rect 21868 19966 21870 20018
rect 21870 19966 21922 20018
rect 21922 19966 21924 20018
rect 21868 19964 21924 19966
rect 21756 19404 21812 19460
rect 22092 19068 22148 19124
rect 21420 17554 21476 17556
rect 21420 17502 21422 17554
rect 21422 17502 21474 17554
rect 21474 17502 21476 17554
rect 21420 17500 21476 17502
rect 21532 17052 21588 17108
rect 21644 18508 21700 18564
rect 22092 18284 22148 18340
rect 20748 15426 20804 15428
rect 20748 15374 20750 15426
rect 20750 15374 20802 15426
rect 20802 15374 20804 15426
rect 20748 15372 20804 15374
rect 21868 17724 21924 17780
rect 21980 17666 22036 17668
rect 21980 17614 21982 17666
rect 21982 17614 22034 17666
rect 22034 17614 22036 17666
rect 21980 17612 22036 17614
rect 21980 16940 22036 16996
rect 22876 20802 22932 20804
rect 22876 20750 22878 20802
rect 22878 20750 22930 20802
rect 22930 20750 22932 20802
rect 22876 20748 22932 20750
rect 22428 20690 22484 20692
rect 22428 20638 22430 20690
rect 22430 20638 22482 20690
rect 22482 20638 22484 20690
rect 22428 20636 22484 20638
rect 23660 22146 23716 22148
rect 23660 22094 23662 22146
rect 23662 22094 23714 22146
rect 23714 22094 23716 22146
rect 23660 22092 23716 22094
rect 25340 26066 25396 26068
rect 25340 26014 25342 26066
rect 25342 26014 25394 26066
rect 25394 26014 25396 26066
rect 25340 26012 25396 26014
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 28588 26796 28644 26852
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 25116 23826 25172 23828
rect 25116 23774 25118 23826
rect 25118 23774 25170 23826
rect 25170 23774 25172 23826
rect 25116 23772 25172 23774
rect 25340 23154 25396 23156
rect 25340 23102 25342 23154
rect 25342 23102 25394 23154
rect 25394 23102 25396 23154
rect 25340 23100 25396 23102
rect 23884 21532 23940 21588
rect 23548 20076 23604 20132
rect 25676 21644 25732 21700
rect 23996 20636 24052 20692
rect 24220 20130 24276 20132
rect 24220 20078 24222 20130
rect 24222 20078 24274 20130
rect 24274 20078 24276 20130
rect 24220 20076 24276 20078
rect 24444 20018 24500 20020
rect 24444 19966 24446 20018
rect 24446 19966 24498 20018
rect 24498 19966 24500 20018
rect 24444 19964 24500 19966
rect 23772 19852 23828 19908
rect 24444 19740 24500 19796
rect 22316 18226 22372 18228
rect 22316 18174 22318 18226
rect 22318 18174 22370 18226
rect 22370 18174 22372 18226
rect 22316 18172 22372 18174
rect 23324 18508 23380 18564
rect 23100 16940 23156 16996
rect 22092 16882 22148 16884
rect 22092 16830 22094 16882
rect 22094 16830 22146 16882
rect 22146 16830 22148 16882
rect 22092 16828 22148 16830
rect 22652 16828 22708 16884
rect 22540 15986 22596 15988
rect 22540 15934 22542 15986
rect 22542 15934 22594 15986
rect 22594 15934 22596 15986
rect 22540 15932 22596 15934
rect 20412 15260 20468 15316
rect 19964 14530 20020 14532
rect 19964 14478 19966 14530
rect 19966 14478 20018 14530
rect 20018 14478 20020 14530
rect 19964 14476 20020 14478
rect 17500 14252 17556 14308
rect 17836 14252 17892 14308
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 21308 14588 21364 14644
rect 24108 18172 24164 18228
rect 23436 16994 23492 16996
rect 23436 16942 23438 16994
rect 23438 16942 23490 16994
rect 23490 16942 23492 16994
rect 23436 16940 23492 16942
rect 25564 20130 25620 20132
rect 25564 20078 25566 20130
rect 25566 20078 25618 20130
rect 25618 20078 25620 20130
rect 25564 20076 25620 20078
rect 25340 20018 25396 20020
rect 25340 19966 25342 20018
rect 25342 19966 25394 20018
rect 25394 19966 25396 20018
rect 25340 19964 25396 19966
rect 25676 19964 25732 20020
rect 26460 23714 26516 23716
rect 26460 23662 26462 23714
rect 26462 23662 26514 23714
rect 26514 23662 26516 23714
rect 26460 23660 26516 23662
rect 26124 22204 26180 22260
rect 25900 21586 25956 21588
rect 25900 21534 25902 21586
rect 25902 21534 25954 21586
rect 25954 21534 25956 21586
rect 25900 21532 25956 21534
rect 28140 23660 28196 23716
rect 37660 23154 37716 23156
rect 37660 23102 37662 23154
rect 37662 23102 37714 23154
rect 37714 23102 37716 23154
rect 37660 23100 37716 23102
rect 28140 23042 28196 23044
rect 28140 22990 28142 23042
rect 28142 22990 28194 23042
rect 28194 22990 28196 23042
rect 28140 22988 28196 22990
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 27804 22428 27860 22484
rect 26572 21644 26628 21700
rect 28588 22482 28644 22484
rect 28588 22430 28590 22482
rect 28590 22430 28642 22482
rect 28642 22430 28644 22482
rect 28588 22428 28644 22430
rect 37660 22370 37716 22372
rect 37660 22318 37662 22370
rect 37662 22318 37714 22370
rect 37714 22318 37716 22370
rect 37660 22316 37716 22318
rect 40012 22204 40068 22260
rect 26460 21586 26516 21588
rect 26460 21534 26462 21586
rect 26462 21534 26514 21586
rect 26514 21534 26516 21586
rect 26460 21532 26516 21534
rect 27692 21586 27748 21588
rect 27692 21534 27694 21586
rect 27694 21534 27746 21586
rect 27746 21534 27748 21586
rect 27692 21532 27748 21534
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 25228 19740 25284 19796
rect 25228 19180 25284 19236
rect 25676 18508 25732 18564
rect 26236 20076 26292 20132
rect 26236 19740 26292 19796
rect 27244 20130 27300 20132
rect 27244 20078 27246 20130
rect 27246 20078 27298 20130
rect 27298 20078 27300 20130
rect 27244 20076 27300 20078
rect 26348 19852 26404 19908
rect 23884 16994 23940 16996
rect 23884 16942 23886 16994
rect 23886 16942 23938 16994
rect 23938 16942 23940 16994
rect 23884 16940 23940 16942
rect 23660 16882 23716 16884
rect 23660 16830 23662 16882
rect 23662 16830 23714 16882
rect 23714 16830 23716 16882
rect 23660 16828 23716 16830
rect 25228 16994 25284 16996
rect 25228 16942 25230 16994
rect 25230 16942 25282 16994
rect 25282 16942 25284 16994
rect 25228 16940 25284 16942
rect 24668 15932 24724 15988
rect 21644 14476 21700 14532
rect 20748 14306 20804 14308
rect 20748 14254 20750 14306
rect 20750 14254 20802 14306
rect 20802 14254 20804 14306
rect 20748 14252 20804 14254
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 24220 4060 24276 4116
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 23548 3612 23604 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 25564 16604 25620 16660
rect 26012 16940 26068 16996
rect 27356 19964 27412 20020
rect 29260 19964 29316 20020
rect 27468 19234 27524 19236
rect 27468 19182 27470 19234
rect 27470 19182 27522 19234
rect 27522 19182 27524 19234
rect 27468 19180 27524 19182
rect 29260 19234 29316 19236
rect 29260 19182 29262 19234
rect 29262 19182 29314 19234
rect 29314 19182 29316 19234
rect 29260 19180 29316 19182
rect 26684 18956 26740 19012
rect 27804 19010 27860 19012
rect 27804 18958 27806 19010
rect 27806 18958 27858 19010
rect 27858 18958 27860 19010
rect 27804 18956 27860 18958
rect 28588 18508 28644 18564
rect 29484 19122 29540 19124
rect 29484 19070 29486 19122
rect 29486 19070 29538 19122
rect 29538 19070 29540 19122
rect 29484 19068 29540 19070
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 29932 19234 29988 19236
rect 29932 19182 29934 19234
rect 29934 19182 29986 19234
rect 29986 19182 29988 19234
rect 29932 19180 29988 19182
rect 30156 19010 30212 19012
rect 30156 18958 30158 19010
rect 30158 18958 30210 19010
rect 30210 18958 30212 19010
rect 30156 18956 30212 18958
rect 39900 20860 39956 20916
rect 37884 19740 37940 19796
rect 37548 18956 37604 19012
rect 40012 20188 40068 20244
rect 40012 19516 40068 19572
rect 37996 19068 38052 19124
rect 40012 18844 40068 18900
rect 37660 18620 37716 18676
rect 29596 18508 29652 18564
rect 29372 18396 29428 18452
rect 37660 18450 37716 18452
rect 37660 18398 37662 18450
rect 37662 18398 37714 18450
rect 37714 18398 37716 18450
rect 37660 18396 37716 18398
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 26572 17554 26628 17556
rect 26572 17502 26574 17554
rect 26574 17502 26626 17554
rect 26626 17502 26628 17554
rect 26572 17500 26628 17502
rect 28364 16716 28420 16772
rect 29260 16770 29316 16772
rect 29260 16718 29262 16770
rect 29262 16718 29314 16770
rect 29314 16718 29316 16770
rect 29260 16716 29316 16718
rect 40012 16828 40068 16884
rect 37884 16716 37940 16772
rect 37660 16604 37716 16660
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 40012 16156 40068 16212
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 26236 4114 26292 4116
rect 26236 4062 26238 4114
rect 26238 4062 26290 4114
rect 26290 4062 26292 4114
rect 26236 4060 26292 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 17490 38220 17500 38276
rect 17556 38220 18620 38276
rect 18676 38220 18686 38276
rect 23538 38220 23548 38276
rect 23604 38220 25564 38276
rect 25620 38220 25630 38276
rect 26226 38220 26236 38276
rect 26292 38220 29372 38276
rect 29428 38220 29438 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 18834 37436 18844 37492
rect 18900 37436 19852 37492
rect 19908 37436 19918 37492
rect 21522 37436 21532 37492
rect 21588 37436 22764 37492
rect 22820 37436 22830 37492
rect 24882 37436 24892 37492
rect 24948 37436 26236 37492
rect 26292 37436 26302 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 16818 36652 16828 36708
rect 16884 36652 18060 36708
rect 18116 36652 18126 36708
rect 20178 36652 20188 36708
rect 20244 36652 22316 36708
rect 22372 36652 22382 36708
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 20178 28588 20188 28644
rect 20244 28588 21196 28644
rect 21252 28588 21262 28644
rect 21410 28476 21420 28532
rect 21476 28476 21868 28532
rect 21924 28476 21934 28532
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 0 27636 800 27664
rect 0 27580 4172 27636
rect 4228 27580 4238 27636
rect 14690 27580 14700 27636
rect 14756 27580 16044 27636
rect 16100 27580 16110 27636
rect 16370 27580 16380 27636
rect 16436 27580 17388 27636
rect 17444 27580 17454 27636
rect 0 27552 800 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 21522 27132 21532 27188
rect 21588 27132 24108 27188
rect 24164 27132 25004 27188
rect 25060 27132 25070 27188
rect 21634 27020 21644 27076
rect 21700 27020 22988 27076
rect 23044 27020 23054 27076
rect 15698 26908 15708 26964
rect 15764 26908 16940 26964
rect 16996 26908 18284 26964
rect 18340 26908 18956 26964
rect 19012 26908 19022 26964
rect 23090 26908 23100 26964
rect 23156 26908 23772 26964
rect 23828 26908 23838 26964
rect 23986 26908 23996 26964
rect 24052 26908 24668 26964
rect 24724 26908 24734 26964
rect 18610 26796 18620 26852
rect 18676 26796 21420 26852
rect 21476 26796 21486 26852
rect 25330 26796 25340 26852
rect 25396 26796 26460 26852
rect 26516 26796 28588 26852
rect 28644 26796 28654 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 17266 26236 17276 26292
rect 17332 26236 18172 26292
rect 18228 26236 20188 26292
rect 20244 26236 20254 26292
rect 19618 26124 19628 26180
rect 19684 26124 21084 26180
rect 21140 26124 21150 26180
rect 24434 26012 24444 26068
rect 24500 26012 25340 26068
rect 25396 26012 25406 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 16146 25564 16156 25620
rect 16212 25564 17388 25620
rect 17444 25564 17454 25620
rect 4274 25452 4284 25508
rect 4340 25452 15484 25508
rect 15540 25452 15550 25508
rect 22530 25452 22540 25508
rect 22596 25452 23660 25508
rect 23716 25452 23726 25508
rect 17938 25340 17948 25396
rect 18004 25340 18732 25396
rect 18788 25340 19292 25396
rect 19348 25340 19358 25396
rect 20402 25340 20412 25396
rect 20468 25340 21196 25396
rect 21252 25340 21868 25396
rect 21924 25340 21934 25396
rect 17154 25228 17164 25284
rect 17220 25228 17724 25284
rect 17780 25228 18620 25284
rect 18676 25228 18686 25284
rect 21074 25228 21084 25284
rect 21140 25228 21756 25284
rect 21812 25228 21822 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 0 24948 800 24976
rect 0 24892 1932 24948
rect 1988 24892 1998 24948
rect 0 24864 800 24892
rect 4274 24668 4284 24724
rect 4340 24668 14812 24724
rect 14868 24668 14878 24724
rect 15138 24556 15148 24612
rect 15204 24556 16268 24612
rect 16324 24556 16940 24612
rect 16996 24556 17500 24612
rect 17556 24556 17566 24612
rect 1922 24444 1932 24500
rect 1988 24444 1998 24500
rect 0 24276 800 24304
rect 1932 24276 1988 24444
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 0 24220 1988 24276
rect 0 24192 800 24220
rect 14354 23996 14364 24052
rect 14420 23996 17052 24052
rect 17108 23996 17118 24052
rect 4274 23884 4284 23940
rect 4340 23884 12236 23940
rect 12292 23884 15036 23940
rect 15092 23884 15708 23940
rect 15764 23884 15774 23940
rect 16818 23884 16828 23940
rect 16884 23884 21532 23940
rect 21588 23884 21598 23940
rect 19618 23772 19628 23828
rect 19684 23772 25116 23828
rect 25172 23772 25182 23828
rect 26450 23660 26460 23716
rect 26516 23660 28140 23716
rect 28196 23660 28206 23716
rect 0 23604 800 23632
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 18274 23436 18284 23492
rect 18340 23436 18956 23492
rect 19012 23436 19022 23492
rect 20402 23436 20412 23492
rect 20468 23436 21420 23492
rect 21476 23436 23884 23492
rect 23940 23436 23950 23492
rect 16594 23324 16604 23380
rect 16660 23324 17388 23380
rect 17444 23324 17454 23380
rect 18834 23324 18844 23380
rect 18900 23324 19516 23380
rect 19572 23324 19582 23380
rect 20178 23324 20188 23380
rect 20244 23324 21308 23380
rect 21364 23324 21374 23380
rect 18498 23212 18508 23268
rect 18564 23212 20300 23268
rect 20356 23212 20366 23268
rect 4274 23100 4284 23156
rect 4340 23100 11452 23156
rect 11508 23100 14140 23156
rect 14196 23100 14206 23156
rect 16930 23100 16940 23156
rect 16996 23100 18060 23156
rect 18116 23100 19964 23156
rect 20020 23100 20030 23156
rect 21074 23100 21084 23156
rect 21140 23100 23660 23156
rect 23716 23100 25340 23156
rect 25396 23100 25406 23156
rect 31892 23100 37660 23156
rect 37716 23100 37726 23156
rect 31892 23044 31948 23100
rect 20514 22988 20524 23044
rect 20580 22988 21644 23044
rect 21700 22988 21710 23044
rect 28130 22988 28140 23044
rect 28196 22988 31948 23044
rect 0 22932 800 22960
rect 41200 22932 42000 22960
rect 0 22876 1932 22932
rect 1988 22876 1998 22932
rect 13682 22876 13692 22932
rect 13748 22876 14812 22932
rect 14868 22876 14878 22932
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 0 22848 800 22876
rect 41200 22848 42000 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 14914 22540 14924 22596
rect 14980 22540 14990 22596
rect 14924 22036 14980 22540
rect 27794 22428 27804 22484
rect 27860 22428 28588 22484
rect 28644 22428 31948 22484
rect 31892 22372 31948 22428
rect 17490 22316 17500 22372
rect 17556 22316 19572 22372
rect 31892 22316 37660 22372
rect 37716 22316 37726 22372
rect 17714 22204 17724 22260
rect 17780 22204 19292 22260
rect 19348 22204 19358 22260
rect 19516 22148 19572 22316
rect 41200 22260 42000 22288
rect 22082 22204 22092 22260
rect 22148 22204 22316 22260
rect 22372 22204 26124 22260
rect 26180 22204 26190 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 41200 22176 42000 22204
rect 15586 22092 15596 22148
rect 15652 22092 17164 22148
rect 17220 22092 18508 22148
rect 18564 22092 18574 22148
rect 19506 22092 19516 22148
rect 19572 22092 20300 22148
rect 20356 22092 20366 22148
rect 22194 22092 22204 22148
rect 22260 22092 23660 22148
rect 23716 22092 23726 22148
rect 14914 21980 14924 22036
rect 14980 21980 14990 22036
rect 15474 21980 15484 22036
rect 15540 21980 18732 22036
rect 18788 21980 18798 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 15026 21756 15036 21812
rect 15092 21756 18844 21812
rect 18900 21756 18910 21812
rect 14802 21644 14812 21700
rect 14868 21644 21252 21700
rect 25666 21644 25676 21700
rect 25732 21644 26572 21700
rect 26628 21644 26638 21700
rect 0 21588 800 21616
rect 21196 21588 21252 21644
rect 0 21532 1932 21588
rect 1988 21532 1998 21588
rect 4274 21532 4284 21588
rect 4340 21532 11340 21588
rect 11396 21532 14140 21588
rect 14196 21532 14206 21588
rect 17602 21532 17612 21588
rect 17668 21532 19404 21588
rect 19460 21532 19470 21588
rect 21186 21532 21196 21588
rect 21252 21532 21262 21588
rect 23874 21532 23884 21588
rect 23940 21532 25900 21588
rect 25956 21532 25966 21588
rect 26450 21532 26460 21588
rect 26516 21532 27692 21588
rect 27748 21532 27758 21588
rect 0 21504 800 21532
rect 17612 21476 17668 21532
rect 4162 21420 4172 21476
rect 4228 21420 17668 21476
rect 17826 21420 17836 21476
rect 17892 21420 18396 21476
rect 18452 21420 18462 21476
rect 13682 21308 13692 21364
rect 13748 21308 14700 21364
rect 14756 21308 14766 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 41200 20916 42000 20944
rect 39890 20860 39900 20916
rect 39956 20860 42000 20916
rect 41200 20832 42000 20860
rect 14018 20748 14028 20804
rect 14084 20748 14924 20804
rect 14980 20748 15484 20804
rect 15540 20748 15550 20804
rect 20066 20748 20076 20804
rect 20132 20748 22876 20804
rect 22932 20748 22942 20804
rect 14242 20636 14252 20692
rect 14308 20636 15708 20692
rect 15764 20636 17276 20692
rect 17332 20636 17342 20692
rect 19170 20636 19180 20692
rect 19236 20636 21532 20692
rect 21588 20636 22428 20692
rect 22484 20636 23996 20692
rect 24052 20636 24062 20692
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 41200 20244 42000 20272
rect 40002 20188 40012 20244
rect 40068 20188 42000 20244
rect 41200 20160 42000 20188
rect 16146 20076 16156 20132
rect 16212 20076 16716 20132
rect 16772 20076 17500 20132
rect 17556 20076 17566 20132
rect 21746 20076 21756 20132
rect 21812 20076 23548 20132
rect 23604 20076 24220 20132
rect 24276 20076 24286 20132
rect 25554 20076 25564 20132
rect 25620 20076 26236 20132
rect 26292 20076 26302 20132
rect 26852 20076 27244 20132
rect 27300 20076 27310 20132
rect 26852 20020 26908 20076
rect 17826 19964 17836 20020
rect 17892 19964 19068 20020
rect 19124 19964 19740 20020
rect 19796 19964 19806 20020
rect 20066 19964 20076 20020
rect 20132 19964 21868 20020
rect 21924 19964 21934 20020
rect 24434 19964 24444 20020
rect 24500 19964 25340 20020
rect 25396 19964 25406 20020
rect 25666 19964 25676 20020
rect 25732 19964 26908 20020
rect 27346 19964 27356 20020
rect 27412 19964 29260 20020
rect 29316 19964 29326 20020
rect 19506 19852 19516 19908
rect 19572 19852 23772 19908
rect 23828 19852 26348 19908
rect 26404 19852 26414 19908
rect 21410 19740 21420 19796
rect 21476 19740 24444 19796
rect 24500 19740 25228 19796
rect 25284 19740 25294 19796
rect 26226 19740 26236 19796
rect 26292 19740 37884 19796
rect 37940 19740 37950 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 41200 19488 42000 19516
rect 17714 19404 17724 19460
rect 17780 19404 18284 19460
rect 18340 19404 18844 19460
rect 18900 19404 18910 19460
rect 20626 19404 20636 19460
rect 20692 19404 21756 19460
rect 21812 19404 21822 19460
rect 18498 19180 18508 19236
rect 18564 19180 20748 19236
rect 20804 19180 20814 19236
rect 25218 19180 25228 19236
rect 25284 19180 27468 19236
rect 27524 19180 27534 19236
rect 29250 19180 29260 19236
rect 29316 19180 29932 19236
rect 29988 19180 29998 19236
rect 18610 19068 18620 19124
rect 18676 19068 18956 19124
rect 19012 19068 19964 19124
rect 20020 19068 21420 19124
rect 21476 19068 22092 19124
rect 22148 19068 22158 19124
rect 29474 19068 29484 19124
rect 29540 19068 37996 19124
rect 38052 19068 38062 19124
rect 15698 18956 15708 19012
rect 15764 18956 16268 19012
rect 16324 18956 18172 19012
rect 18228 18956 18238 19012
rect 18722 18956 18732 19012
rect 18788 18956 19516 19012
rect 19572 18956 20524 19012
rect 20580 18956 20590 19012
rect 26674 18956 26684 19012
rect 26740 18956 27804 19012
rect 27860 18956 27870 19012
rect 30146 18956 30156 19012
rect 30212 18956 37548 19012
rect 37604 18956 37614 19012
rect 41200 18900 42000 18928
rect 40002 18844 40012 18900
rect 40068 18844 42000 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 41200 18816 42000 18844
rect 18162 18620 18172 18676
rect 18228 18620 20636 18676
rect 20692 18620 20702 18676
rect 31892 18620 37660 18676
rect 37716 18620 37726 18676
rect 31892 18564 31948 18620
rect 15586 18508 15596 18564
rect 15652 18508 17500 18564
rect 17556 18508 20076 18564
rect 20132 18508 20142 18564
rect 20738 18508 20748 18564
rect 20804 18508 21644 18564
rect 21700 18508 21710 18564
rect 23314 18508 23324 18564
rect 23380 18508 25676 18564
rect 25732 18508 25742 18564
rect 28578 18508 28588 18564
rect 28644 18508 29596 18564
rect 29652 18508 31948 18564
rect 4274 18396 4284 18452
rect 4340 18396 9996 18452
rect 10052 18396 10062 18452
rect 12002 18396 12012 18452
rect 12068 18396 12796 18452
rect 12852 18396 12862 18452
rect 13020 18396 15484 18452
rect 15540 18396 15550 18452
rect 16706 18396 16716 18452
rect 16772 18396 18396 18452
rect 18452 18396 18462 18452
rect 29362 18396 29372 18452
rect 29428 18396 37660 18452
rect 37716 18396 37726 18452
rect 9996 18340 10052 18396
rect 13020 18340 13076 18396
rect 9996 18284 13076 18340
rect 14242 18284 14252 18340
rect 14308 18284 15596 18340
rect 15652 18284 15662 18340
rect 17602 18284 17612 18340
rect 17668 18284 19628 18340
rect 19684 18284 19694 18340
rect 20738 18284 20748 18340
rect 20804 18284 22092 18340
rect 22148 18284 22158 18340
rect 0 18228 800 18256
rect 41200 18228 42000 18256
rect 0 18172 1932 18228
rect 1988 18172 1998 18228
rect 14802 18172 14812 18228
rect 14868 18172 15820 18228
rect 15876 18172 16492 18228
rect 16548 18172 16558 18228
rect 16818 18172 16828 18228
rect 16884 18172 17948 18228
rect 18004 18172 18620 18228
rect 18676 18172 18686 18228
rect 18834 18172 18844 18228
rect 18900 18172 19404 18228
rect 19460 18172 19470 18228
rect 22306 18172 22316 18228
rect 22372 18172 24108 18228
rect 24164 18172 24174 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 0 18144 800 18172
rect 41200 18144 42000 18172
rect 20290 18060 20300 18116
rect 20356 18060 20748 18116
rect 20804 18060 20814 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 13906 17836 13916 17892
rect 13972 17836 16716 17892
rect 16772 17836 17724 17892
rect 17780 17836 21308 17892
rect 21364 17836 21374 17892
rect 12114 17724 12124 17780
rect 12180 17724 14028 17780
rect 14084 17724 14094 17780
rect 16370 17724 16380 17780
rect 16436 17724 17276 17780
rect 17332 17724 18172 17780
rect 18228 17724 18238 17780
rect 18834 17724 18844 17780
rect 18900 17724 19404 17780
rect 19460 17724 21420 17780
rect 21476 17724 21868 17780
rect 21924 17724 21934 17780
rect 12786 17612 12796 17668
rect 12852 17612 13580 17668
rect 13636 17612 15036 17668
rect 15092 17612 15102 17668
rect 16482 17612 16492 17668
rect 16548 17612 18060 17668
rect 18116 17612 18126 17668
rect 18274 17612 18284 17668
rect 18340 17612 19516 17668
rect 19572 17612 21980 17668
rect 22036 17612 22046 17668
rect 14354 17500 14364 17556
rect 14420 17500 16156 17556
rect 16212 17500 16222 17556
rect 21410 17500 21420 17556
rect 21476 17500 26572 17556
rect 26628 17500 26638 17556
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 19954 17052 19964 17108
rect 20020 17052 21532 17108
rect 21588 17052 21598 17108
rect 20300 16940 20636 16996
rect 20692 16940 20702 16996
rect 21970 16940 21980 16996
rect 22036 16940 23100 16996
rect 23156 16940 23436 16996
rect 23492 16940 23502 16996
rect 23874 16940 23884 16996
rect 23940 16940 25228 16996
rect 25284 16940 26012 16996
rect 26068 16940 26078 16996
rect 20300 16884 20356 16940
rect 41200 16884 42000 16912
rect 20178 16828 20188 16884
rect 20244 16828 20356 16884
rect 20514 16828 20524 16884
rect 20580 16828 22092 16884
rect 22148 16828 22158 16884
rect 22642 16828 22652 16884
rect 22708 16828 23660 16884
rect 23716 16828 23726 16884
rect 40002 16828 40012 16884
rect 40068 16828 42000 16884
rect 41200 16800 42000 16828
rect 28354 16716 28364 16772
rect 28420 16716 29260 16772
rect 29316 16716 37884 16772
rect 37940 16716 37950 16772
rect 25554 16604 25564 16660
rect 25620 16604 37660 16660
rect 37716 16604 37726 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 41200 16212 42000 16240
rect 40002 16156 40012 16212
rect 40068 16156 42000 16212
rect 41200 16128 42000 16156
rect 22530 15932 22540 15988
rect 22596 15932 24668 15988
rect 24724 15932 24734 15988
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 16818 15372 16828 15428
rect 16884 15372 20748 15428
rect 20804 15372 20814 15428
rect 18498 15260 18508 15316
rect 18564 15260 19180 15316
rect 19236 15260 20076 15316
rect 20132 15260 20412 15316
rect 20468 15260 20478 15316
rect 18050 15148 18060 15204
rect 18116 15148 19068 15204
rect 19124 15148 19740 15204
rect 19796 15148 19806 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 18946 14588 18956 14644
rect 19012 14588 19516 14644
rect 19572 14588 21308 14644
rect 21364 14588 21374 14644
rect 19954 14476 19964 14532
rect 20020 14476 21644 14532
rect 21700 14476 21710 14532
rect 15138 14252 15148 14308
rect 15204 14252 16156 14308
rect 16212 14252 16940 14308
rect 16996 14252 17500 14308
rect 17556 14252 17836 14308
rect 17892 14252 20748 14308
rect 20804 14252 20814 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 24210 4060 24220 4116
rect 24276 4060 26236 4116
rect 26292 4060 26302 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 23538 3612 23548 3668
rect 23604 3612 25564 3668
rect 25620 3612 25630 3668
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _094_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _095_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18480 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _096_
timestamp 1698175906
transform -1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _097_
timestamp 1698175906
transform -1 0 16800 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _098_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18032 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _099_
timestamp 1698175906
transform 1 0 19936 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21728 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _101_
timestamp 1698175906
transform -1 0 20608 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19600 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _103_
timestamp 1698175906
transform -1 0 19040 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_
timestamp 1698175906
transform -1 0 16128 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16912 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_
timestamp 1698175906
transform -1 0 18368 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _107_
timestamp 1698175906
transform 1 0 18368 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _108_
timestamp 1698175906
transform 1 0 19488 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _109_
timestamp 1698175906
transform -1 0 24304 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _110_
timestamp 1698175906
transform -1 0 20272 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _111_
timestamp 1698175906
transform 1 0 17136 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _112_
timestamp 1698175906
transform -1 0 20384 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_
timestamp 1698175906
transform -1 0 18032 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _114_
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _115_
timestamp 1698175906
transform 1 0 22848 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _116_
timestamp 1698175906
transform 1 0 18032 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _117_
timestamp 1698175906
transform 1 0 19936 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _118_
timestamp 1698175906
transform 1 0 20384 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20272 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform -1 0 19936 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22512 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698175906
transform 1 0 17808 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23296 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _125_
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _126_
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21280 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _128_
timestamp 1698175906
transform -1 0 24304 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _129_
timestamp 1698175906
transform -1 0 21056 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18704 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _131_
timestamp 1698175906
transform 1 0 19152 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _132_
timestamp 1698175906
transform 1 0 19824 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _133_
timestamp 1698175906
transform 1 0 21504 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _134_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20496 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19040 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _136_
timestamp 1698175906
transform -1 0 18816 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _137_
timestamp 1698175906
transform -1 0 18032 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16912 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _139_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19152 0 -1 18816
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _140_
timestamp 1698175906
transform -1 0 15456 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _141_
timestamp 1698175906
transform -1 0 15792 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _142_
timestamp 1698175906
transform -1 0 15344 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _143_
timestamp 1698175906
transform -1 0 13776 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _144_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21504 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _145_
timestamp 1698175906
transform 1 0 21952 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _146_
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _147_
timestamp 1698175906
transform -1 0 24640 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _148_
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _149_
timestamp 1698175906
transform -1 0 22176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _150_
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _151_
timestamp 1698175906
transform -1 0 26768 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _152_
timestamp 1698175906
transform 1 0 18256 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _153_
timestamp 1698175906
transform -1 0 20384 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _154_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24976 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _155_
timestamp 1698175906
transform -1 0 19040 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _156_
timestamp 1698175906
transform -1 0 17696 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _157_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20160 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _158_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _159_
timestamp 1698175906
transform -1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform 1 0 27328 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _161_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26208 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _162_
timestamp 1698175906
transform -1 0 28000 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _163_
timestamp 1698175906
transform -1 0 28000 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _164_
timestamp 1698175906
transform 1 0 20384 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _165_
timestamp 1698175906
transform 1 0 23408 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _166_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 26880 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _167_
timestamp 1698175906
transform 1 0 27104 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _168_
timestamp 1698175906
transform -1 0 27104 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _169_
timestamp 1698175906
transform -1 0 25872 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _170_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24640 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _171_
timestamp 1698175906
transform -1 0 18144 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _172_
timestamp 1698175906
transform -1 0 16352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _173_
timestamp 1698175906
transform 1 0 22064 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _174_
timestamp 1698175906
transform 1 0 22624 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _175_
timestamp 1698175906
transform -1 0 15904 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _176_
timestamp 1698175906
transform -1 0 14448 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _177_
timestamp 1698175906
transform -1 0 19264 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _178_
timestamp 1698175906
transform 1 0 13888 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _179_
timestamp 1698175906
transform 1 0 14560 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _180_
timestamp 1698175906
transform -1 0 21952 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _181_
timestamp 1698175906
transform 1 0 13888 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _182_
timestamp 1698175906
transform 1 0 14448 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _183_
timestamp 1698175906
transform -1 0 18144 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _184_
timestamp 1698175906
transform 1 0 15344 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _185_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16128 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _186_
timestamp 1698175906
transform 1 0 18256 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _187_
timestamp 1698175906
transform -1 0 19824 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _188_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18368 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _189_
timestamp 1698175906
transform 1 0 21616 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _190_
timestamp 1698175906
transform 1 0 22960 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _191_
timestamp 1698175906
transform 1 0 20832 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _192_
timestamp 1698175906
transform 1 0 15904 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _193_
timestamp 1698175906
transform 1 0 17584 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_
timestamp 1698175906
transform 1 0 13440 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1698175906
transform 1 0 11760 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _196_
timestamp 1698175906
transform 1 0 23408 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _197_
timestamp 1698175906
transform -1 0 22736 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _198_
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _199_
timestamp 1698175906
transform 1 0 15456 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _200_
timestamp 1698175906
transform 1 0 26208 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1698175906
transform 1 0 25536 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_
timestamp 1698175906
transform 1 0 25536 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform 1 0 23184 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform 1 0 13776 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform 1 0 21616 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform -1 0 13104 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform -1 0 14560 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform -1 0 14448 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform -1 0 15344 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 17360 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _211_
timestamp 1698175906
transform -1 0 15344 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _212_
timestamp 1698175906
transform 1 0 29680 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _213_
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _214_
timestamp 1698175906
transform 1 0 28896 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _215_
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _216_
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _217_
timestamp 1698175906
transform -1 0 16016 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__A1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21392 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__CLK
timestamp 1698175906
transform -1 0 18368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__CLK
timestamp 1698175906
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__CLK
timestamp 1698175906
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1698175906
transform 1 0 15008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__CLK
timestamp 1698175906
transform 1 0 18928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform 1 0 16912 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 13552 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 15344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 14672 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 16240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 17584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output22_I
timestamp 1698175906
transform 1 0 24304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 20944 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 22624 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout27
timestamp 1698175906
transform -1 0 29792 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 28000 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 31584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_139
timestamp 1698175906
transform 1 0 16912 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_147
timestamp 1698175906
transform 1 0 17808 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_151
timestamp 1698175906
transform 1 0 18256 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_158 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19040 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_144
timestamp 1698175906
transform 1 0 17472 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_174
timestamp 1698175906
transform 1 0 20832 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698175906
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_127
timestamp 1698175906
transform 1 0 15568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_129
timestamp 1698175906
transform 1 0 15792 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_171
timestamp 1698175906
transform 1 0 20496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_183
timestamp 1698175906
transform 1 0 21840 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_215
timestamp 1698175906
transform 1 0 25424 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_231
timestamp 1698175906
transform 1 0 27216 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_239
timestamp 1698175906
transform 1 0 28112 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698175906
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_146
timestamp 1698175906
transform 1 0 17696 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_163
timestamp 1698175906
transform 1 0 19600 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_165
timestamp 1698175906
transform 1 0 19824 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_176
timestamp 1698175906
transform 1 0 21056 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_180
timestamp 1698175906
transform 1 0 21504 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_139
timestamp 1698175906
transform 1 0 16912 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_155
timestamp 1698175906
transform 1 0 18704 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698175906
transform 1 0 20720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_222
timestamp 1698175906
transform 1 0 26208 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_238
timestamp 1698175906
transform 1 0 28000 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_104
timestamp 1698175906
transform 1 0 12992 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698175906
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_146
timestamp 1698175906
transform 1 0 17696 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_156
timestamp 1698175906
transform 1 0 18816 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_164
timestamp 1698175906
transform 1 0 19712 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_166
timestamp 1698175906
transform 1 0 19936 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_172
timestamp 1698175906
transform 1 0 20608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_174
timestamp 1698175906
transform 1 0 20832 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_189
timestamp 1698175906
transform 1 0 22512 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_205
timestamp 1698175906
transform 1 0 24304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_218
timestamp 1698175906
transform 1 0 25760 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_251
timestamp 1698175906
transform 1 0 29456 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_267
timestamp 1698175906
transform 1 0 31248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_275
timestamp 1698175906
transform 1 0 32144 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 36512 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 37408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_69
timestamp 1698175906
transform 1 0 9072 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_73
timestamp 1698175906
transform 1 0 9520 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_75
timestamp 1698175906
transform 1 0 9744 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_117
timestamp 1698175906
transform 1 0 14448 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_121
timestamp 1698175906
transform 1 0 14896 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_124
timestamp 1698175906
transform 1 0 15232 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_128
timestamp 1698175906
transform 1 0 15680 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_130
timestamp 1698175906
transform 1 0 15904 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_139
timestamp 1698175906
transform 1 0 16912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_159
timestamp 1698175906
transform 1 0 19152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698175906
transform 1 0 20608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_185
timestamp 1698175906
transform 1 0 22064 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_193
timestamp 1698175906
transform 1 0 22960 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_197
timestamp 1698175906
transform 1 0 23408 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_205
timestamp 1698175906
transform 1 0 24304 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_221
timestamp 1698175906
transform 1 0 26096 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_238
timestamp 1698175906
transform 1 0 28000 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_242
timestamp 1698175906
transform 1 0 28448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 4480 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 8064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_88
timestamp 1698175906
transform 1 0 11200 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_92
timestamp 1698175906
transform 1 0 11648 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_130
timestamp 1698175906
transform 1 0 15904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_155
timestamp 1698175906
transform 1 0 18704 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_193
timestamp 1698175906
transform 1 0 22960 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_245
timestamp 1698175906
transform 1 0 28784 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_252
timestamp 1698175906
transform 1 0 29568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_268
timestamp 1698175906
transform 1 0 31360 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698175906
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_115
timestamp 1698175906
transform 1 0 14224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_119
timestamp 1698175906
transform 1 0 14672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_138
timestamp 1698175906
transform 1 0 16800 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_149
timestamp 1698175906
transform 1 0 18032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_157
timestamp 1698175906
transform 1 0 18928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_159
timestamp 1698175906
transform 1 0 19152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_182
timestamp 1698175906
transform 1 0 21728 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_190
timestamp 1698175906
transform 1 0 22624 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_194
timestamp 1698175906
transform 1 0 23072 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_224
timestamp 1698175906
transform 1 0 26432 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_237
timestamp 1698175906
transform 1 0 27888 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_259
timestamp 1698175906
transform 1 0 30352 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_291
timestamp 1698175906
transform 1 0 33936 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_307
timestamp 1698175906
transform 1 0 35728 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_104
timestamp 1698175906
transform 1 0 12992 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_111
timestamp 1698175906
transform 1 0 13776 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_127
timestamp 1698175906
transform 1 0 15568 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_135
timestamp 1698175906
transform 1 0 16464 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_168
timestamp 1698175906
transform 1 0 20160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_187
timestamp 1698175906
transform 1 0 22288 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_195
timestamp 1698175906
transform 1 0 23184 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_208
timestamp 1698175906
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_219
timestamp 1698175906
transform 1 0 25872 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_235
timestamp 1698175906
transform 1 0 27664 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_243
timestamp 1698175906
transform 1 0 28560 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_247
timestamp 1698175906
transform 1 0 29008 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_254
timestamp 1698175906
transform 1 0 29792 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_270
timestamp 1698175906
transform 1 0 31584 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_111
timestamp 1698175906
transform 1 0 13776 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_240
timestamp 1698175906
transform 1 0 28224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_129
timestamp 1698175906
transform 1 0 15792 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_137
timestamp 1698175906
transform 1 0 16688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698175906
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_144
timestamp 1698175906
transform 1 0 17472 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_228
timestamp 1698175906
transform 1 0 26880 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_232
timestamp 1698175906
transform 1 0 27328 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_238
timestamp 1698175906
transform 1 0 28000 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_270
timestamp 1698175906
transform 1 0 31584 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 4480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_111
timestamp 1698175906
transform 1 0 13776 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_117
timestamp 1698175906
transform 1 0 14448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_121
timestamp 1698175906
transform 1 0 14896 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_137
timestamp 1698175906
transform 1 0 16688 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_145
timestamp 1698175906
transform 1 0 17584 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_158
timestamp 1698175906
transform 1 0 19040 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_170
timestamp 1698175906
transform 1 0 20384 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_179
timestamp 1698175906
transform 1 0 21392 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_186
timestamp 1698175906
transform 1 0 22176 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_194
timestamp 1698175906
transform 1 0 23072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_196
timestamp 1698175906
transform 1 0 23296 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_202
timestamp 1698175906
transform 1 0 23968 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_210
timestamp 1698175906
transform 1 0 24864 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_214
timestamp 1698175906
transform 1 0 25312 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 4480 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_88
timestamp 1698175906
transform 1 0 11200 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_123
timestamp 1698175906
transform 1 0 15120 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_127
timestamp 1698175906
transform 1 0 15568 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_135
timestamp 1698175906
transform 1 0 16464 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_150
timestamp 1698175906
transform 1 0 18144 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_203
timestamp 1698175906
transform 1 0 24080 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698175906
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_241
timestamp 1698175906
transform 1 0 28336 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698175906
transform 1 0 31920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_115
timestamp 1698175906
transform 1 0 14224 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_130
timestamp 1698175906
transform 1 0 15904 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698175906
transform 1 0 20608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_181
timestamp 1698175906
transform 1 0 21616 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_197
timestamp 1698175906
transform 1 0 23408 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_205
timestamp 1698175906
transform 1 0 24304 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_209
timestamp 1698175906
transform 1 0 24752 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_219
timestamp 1698175906
transform 1 0 25872 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_221
timestamp 1698175906
transform 1 0 26096 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_227
timestamp 1698175906
transform 1 0 26768 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 4480 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 8064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_88
timestamp 1698175906
transform 1 0 11200 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_131
timestamp 1698175906
transform 1 0 16016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_135
timestamp 1698175906
transform 1 0 16464 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_146
timestamp 1698175906
transform 1 0 17696 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_178
timestamp 1698175906
transform 1 0 21280 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_194
timestamp 1698175906
transform 1 0 23072 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_202
timestamp 1698175906
transform 1 0 23968 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698175906
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_150
timestamp 1698175906
transform 1 0 18144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_157
timestamp 1698175906
transform 1 0 18928 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_165
timestamp 1698175906
transform 1 0 19824 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698175906
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_186
timestamp 1698175906
transform 1 0 22176 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_194
timestamp 1698175906
transform 1 0 23072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_196
timestamp 1698175906
transform 1 0 23296 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_226
timestamp 1698175906
transform 1 0 26656 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698175906
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_104
timestamp 1698175906
transform 1 0 12992 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_108
timestamp 1698175906
transform 1 0 13440 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_110
timestamp 1698175906
transform 1 0 13664 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_148
timestamp 1698175906
transform 1 0 17920 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_158
timestamp 1698175906
transform 1 0 19040 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_191
timestamp 1698175906
transform 1 0 22736 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698175906
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_217
timestamp 1698175906
transform 1 0 25648 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_249
timestamp 1698175906
transform 1 0 29232 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_265
timestamp 1698175906
transform 1 0 31024 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_273
timestamp 1698175906
transform 1 0 31920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 32368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_123
timestamp 1698175906
transform 1 0 15120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_125
timestamp 1698175906
transform 1 0 15344 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_155
timestamp 1698175906
transform 1 0 18704 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_159
timestamp 1698175906
transform 1 0 19152 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_161
timestamp 1698175906
transform 1 0 19376 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_167
timestamp 1698175906
transform 1 0 20048 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_186
timestamp 1698175906
transform 1 0 22176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_190
timestamp 1698175906
transform 1 0 22624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_197
timestamp 1698175906
transform 1 0 23408 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_199
timestamp 1698175906
transform 1 0 23632 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_205
timestamp 1698175906
transform 1 0 24304 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_237
timestamp 1698175906
transform 1 0 27888 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_104
timestamp 1698175906
transform 1 0 12992 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_120
timestamp 1698175906
transform 1 0 14784 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_128
timestamp 1698175906
transform 1 0 15680 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_134
timestamp 1698175906
transform 1 0 16352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_138
timestamp 1698175906
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_146
timestamp 1698175906
transform 1 0 17696 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_182
timestamp 1698175906
transform 1 0 21728 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_214
timestamp 1698175906
transform 1 0 25312 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_230
timestamp 1698175906
transform 1 0 27104 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_238
timestamp 1698175906
transform 1 0 28000 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_242
timestamp 1698175906
transform 1 0 28448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698175906
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_165
timestamp 1698175906
transform 1 0 19824 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_173
timestamp 1698175906
transform 1 0 20720 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_203
timestamp 1698175906
transform 1 0 24080 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_207
timestamp 1698175906
transform 1 0 24528 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_239
timestamp 1698175906
transform 1 0 28112 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_243
timestamp 1698175906
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_150
timestamp 1698175906
transform 1 0 18144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_154
timestamp 1698175906
transform 1 0 18592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 28000 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 31584 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_266
timestamp 1698175906
transform 1 0 31136 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_270
timestamp 1698175906
transform 1 0 31584 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 4480 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 37520 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 4480 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 16912 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform -1 0 4480 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 18704 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 4480 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 37520 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 21616 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698175906
transform 1 0 21280 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 20160 41200 20272 42000 0 FreeSans 448 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 41200 18816 42000 18928 0 FreeSans 448 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 41200 16800 42000 16912 0 FreeSans 448 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 16800 41200 16912 42000 0 FreeSans 448 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 41200 20160 42000 20272 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 18816 41200 18928 42000 0 FreeSans 448 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 41200 16128 42000 16240 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 17472 41200 17584 42000 0 FreeSans 448 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 26208 41200 26320 42000 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 23520 41200 23632 42000 0 FreeSans 448 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 21504 41200 21616 42000 0 FreeSans 448 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 24864 41200 24976 42000 0 FreeSans 448 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 18312 23632 18312 23632 0 _000_
rlabel metal2 19992 27384 19992 27384 0 _001_
rlabel metal2 23128 27496 23128 27496 0 _002_
rlabel metal2 23912 16408 23912 16408 0 _003_
rlabel metal2 21784 22736 21784 22736 0 _004_
rlabel metal3 18816 15400 18816 15400 0 _005_
rlabel metal2 18536 13216 18536 13216 0 _006_
rlabel metal2 14392 17248 14392 17248 0 _007_
rlabel metal2 12712 19320 12712 19320 0 _008_
rlabel metal2 24136 25144 24136 25144 0 _009_
rlabel metal2 21840 26936 21840 26936 0 _010_
rlabel metal2 26040 23296 26040 23296 0 _011_
rlabel metal2 16408 27384 16408 27384 0 _012_
rlabel metal2 27160 17192 27160 17192 0 _013_
rlabel metal2 26488 22008 26488 22008 0 _014_
rlabel metal2 26488 19208 26488 19208 0 _015_
rlabel metal2 24136 19544 24136 19544 0 _016_
rlabel metal3 15400 27608 15400 27608 0 _017_
rlabel metal2 22568 15512 22568 15512 0 _018_
rlabel metal3 13104 17752 13104 17752 0 _019_
rlabel metal2 13608 22960 13608 22960 0 _020_
rlabel metal2 13496 21392 13496 21392 0 _021_
rlabel metal2 14392 24304 14392 24304 0 _022_
rlabel metal2 21784 25872 21784 25872 0 _023_
rlabel metal3 27076 20104 27076 20104 0 _024_
rlabel metal2 25480 23968 25480 23968 0 _025_
rlabel metal3 19656 18984 19656 18984 0 _026_
rlabel metal2 19432 23016 19432 23016 0 _027_
rlabel metal2 17584 27720 17584 27720 0 _028_
rlabel metal2 23800 19936 23800 19936 0 _029_
rlabel metal3 24024 17528 24024 17528 0 _030_
rlabel metal2 28280 17080 28280 17080 0 _031_
rlabel metal2 26712 18312 26712 18312 0 _032_
rlabel metal2 27440 17640 27440 17640 0 _033_
rlabel metal3 27104 21560 27104 21560 0 _034_
rlabel metal2 21784 20048 21784 20048 0 _035_
rlabel metal3 24920 21560 24920 21560 0 _036_
rlabel metal2 27048 19880 27048 19880 0 _037_
rlabel metal3 24920 19992 24920 19992 0 _038_
rlabel metal3 16800 25592 16800 25592 0 _039_
rlabel metal2 22456 15792 22456 15792 0 _040_
rlabel metal2 14280 18088 14280 18088 0 _041_
rlabel metal2 18984 22456 18984 22456 0 _042_
rlabel metal2 14392 22512 14392 22512 0 _043_
rlabel metal3 21224 21616 21224 21616 0 _044_
rlabel metal2 14448 20776 14448 20776 0 _045_
rlabel metal2 16632 23632 16632 23632 0 _046_
rlabel metal2 16016 23912 16016 23912 0 _047_
rlabel metal2 18536 22960 18536 22960 0 _048_
rlabel metal2 17976 17920 17976 17920 0 _049_
rlabel metal3 21784 19096 21784 19096 0 _050_
rlabel metal2 16856 19208 16856 19208 0 _051_
rlabel metal2 20664 17584 20664 17584 0 _052_
rlabel metal2 17416 25088 17416 25088 0 _053_
rlabel metal2 21560 27832 21560 27832 0 _054_
rlabel metal2 20216 28336 20216 28336 0 _055_
rlabel metal3 18872 15288 18872 15288 0 _056_
rlabel metal2 18424 22008 18424 22008 0 _057_
rlabel metal3 17080 22120 17080 22120 0 _058_
rlabel metal2 20160 17528 20160 17528 0 _059_
rlabel metal2 18872 19712 18872 19712 0 _060_
rlabel metal3 19040 23128 19040 23128 0 _061_
rlabel metal2 19376 26936 19376 26936 0 _062_
rlabel metal3 23464 26936 23464 26936 0 _063_
rlabel metal3 20048 26824 20048 26824 0 _064_
rlabel metal2 20104 19656 20104 19656 0 _065_
rlabel metal2 19768 19712 19768 19712 0 _066_
rlabel metal3 16856 20104 16856 20104 0 _067_
rlabel metal3 22344 27048 22344 27048 0 _068_
rlabel metal3 19656 19208 19656 19208 0 _069_
rlabel metal2 20496 19992 20496 19992 0 _070_
rlabel metal2 21392 19992 21392 19992 0 _071_
rlabel metal3 20832 14504 20832 14504 0 _072_
rlabel metal2 22120 18368 22120 18368 0 _073_
rlabel metal2 22008 16408 22008 16408 0 _074_
rlabel metal2 22680 16464 22680 16464 0 _075_
rlabel metal2 23128 16912 23128 16912 0 _076_
rlabel metal2 23800 17360 23800 17360 0 _077_
rlabel metal2 22008 18368 22008 18368 0 _078_
rlabel metal2 20552 17304 20552 17304 0 _079_
rlabel metal2 26152 22568 26152 22568 0 _080_
rlabel metal2 19656 14868 19656 14868 0 _081_
rlabel metal3 20776 23352 20776 23352 0 _082_
rlabel metal2 21672 22792 21672 22792 0 _083_
rlabel metal2 18872 13664 18872 13664 0 _084_
rlabel metal2 18088 17360 18088 17360 0 _085_
rlabel metal2 17752 18088 17752 18088 0 _086_
rlabel metal2 18424 22848 18424 22848 0 _087_
rlabel metal2 15512 21224 15512 21224 0 _088_
rlabel metal2 15288 21280 15288 21280 0 _089_
rlabel metal2 13608 20160 13608 20160 0 _090_
rlabel metal2 22232 21448 22232 21448 0 _091_
rlabel metal2 24024 20944 24024 20944 0 _092_
rlabel metal2 24472 25424 24472 25424 0 _093_
rlabel metal3 2478 27608 2478 27608 0 clk
rlabel metal2 22904 21112 22904 21112 0 clknet_0_clk
rlabel metal2 15736 26992 15736 26992 0 clknet_1_0__leaf_clk
rlabel metal2 22176 27832 22176 27832 0 clknet_1_1__leaf_clk
rlabel metal2 21336 14560 21336 14560 0 dut43.count\[0\]
rlabel metal2 20664 14364 20664 14364 0 dut43.count\[1\]
rlabel metal2 17304 17696 17304 17696 0 dut43.count\[2\]
rlabel metal2 15848 18704 15848 18704 0 dut43.count\[3\]
rlabel metal2 11480 23072 11480 23072 0 net1
rlabel metal2 27832 22064 27832 22064 0 net10
rlabel metal2 14840 24248 14840 24248 0 net11
rlabel metal2 15680 23800 15680 23800 0 net12
rlabel metal2 37576 19488 37576 19488 0 net13
rlabel metal3 33768 19096 33768 19096 0 net14
rlabel metal2 18592 27160 18592 27160 0 net15
rlabel metal2 24584 5964 24584 5964 0 net16
rlabel metal2 10024 18088 10024 18088 0 net17
rlabel metal2 28168 23352 28168 23352 0 net18
rlabel metal2 37688 16744 37688 16744 0 net19
rlabel metal2 20832 36456 20832 36456 0 net2
rlabel metal2 17752 32256 17752 32256 0 net20
rlabel metal2 28616 32424 28616 32424 0 net21
rlabel metal2 24360 34076 24360 34076 0 net22
rlabel metal2 15512 25200 15512 25200 0 net23
rlabel metal3 21672 28504 21672 28504 0 net24
rlabel metal2 24696 28112 24696 28112 0 net25
rlabel metal2 21280 31920 21280 31920 0 net26
rlabel metal2 29288 20048 29288 20048 0 net27
rlabel metal2 29400 18480 29400 18480 0 net3
rlabel metal2 28616 18424 28616 18424 0 net4
rlabel metal2 37912 20664 37912 20664 0 net5
rlabel metal2 28392 16464 28392 16464 0 net6
rlabel metal3 24584 16968 24584 16968 0 net7
rlabel metal2 11368 21504 11368 21504 0 net8
rlabel metal2 17080 27160 17080 27160 0 net9
rlabel metal3 1358 22904 1358 22904 0 segm[0]
rlabel metal2 20216 38962 20216 38962 0 segm[10]
rlabel metal3 40642 18200 40642 18200 0 segm[11]
rlabel metal2 40040 19096 40040 19096 0 segm[12]
rlabel metal2 39928 21168 39928 21168 0 segm[13]
rlabel metal2 40040 17304 40040 17304 0 segm[1]
rlabel metal2 24248 2422 24248 2422 0 segm[2]
rlabel metal3 1358 21560 1358 21560 0 segm[3]
rlabel metal2 16856 38962 16856 38962 0 segm[4]
rlabel metal2 40040 22344 40040 22344 0 segm[5]
rlabel metal3 1358 24248 1358 24248 0 segm[6]
rlabel metal3 1358 23576 1358 23576 0 segm[7]
rlabel metal2 40040 19656 40040 19656 0 segm[8]
rlabel metal2 40040 20552 40040 20552 0 segm[9]
rlabel metal3 19376 37464 19376 37464 0 sel[0]
rlabel metal2 23576 2198 23576 2198 0 sel[10]
rlabel metal3 1358 18200 1358 18200 0 sel[11]
rlabel metal3 40642 22904 40642 22904 0 sel[1]
rlabel metal2 40040 16408 40040 16408 0 sel[2]
rlabel metal2 17528 39746 17528 39746 0 sel[3]
rlabel metal2 26264 39746 26264 39746 0 sel[4]
rlabel metal2 23576 39746 23576 39746 0 sel[5]
rlabel metal3 1358 24920 1358 24920 0 sel[6]
rlabel metal2 21560 39354 21560 39354 0 sel[7]
rlabel metal2 24920 39354 24920 39354 0 sel[8]
rlabel metal2 22232 39746 22232 39746 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
