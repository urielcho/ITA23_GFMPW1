magic
tech gf180mcuD
magscale 1 5
timestamp 1699642151
<< obsm1 >>
rect 672 1538 20328 19238
<< metal2 >>
rect 8736 20600 8792 21000
rect 9744 20600 9800 21000
rect 10416 20600 10472 21000
rect 10752 20600 10808 21000
rect 11088 20600 11144 21000
rect 12096 20600 12152 21000
rect 3360 0 3416 400
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 10080 0 10136 400
rect 11424 0 11480 400
rect 12096 0 12152 400
rect 13104 0 13160 400
<< obsm2 >>
rect 966 20570 8706 20600
rect 8822 20570 9714 20600
rect 9830 20570 10386 20600
rect 10502 20570 10722 20600
rect 10838 20570 11058 20600
rect 11174 20570 12066 20600
rect 12182 20570 20146 20600
rect 966 430 20146 20570
rect 966 400 3330 430
rect 3446 400 8706 430
rect 8822 400 9042 430
rect 9158 400 10050 430
rect 10166 400 11394 430
rect 11510 400 12066 430
rect 12182 400 13074 430
rect 13190 400 20146 430
<< metal3 >>
rect 20600 17136 21000 17192
rect 0 13776 400 13832
rect 20600 13440 21000 13496
rect 20600 13104 21000 13160
rect 0 12768 400 12824
rect 0 12432 400 12488
rect 20600 12432 21000 12488
rect 20600 11424 21000 11480
rect 20600 11088 21000 11144
rect 20600 10416 21000 10472
rect 20600 10080 21000 10136
rect 20600 9408 21000 9464
rect 20600 8736 21000 8792
rect 20600 7728 21000 7784
<< obsm3 >>
rect 400 17222 20600 19222
rect 400 17106 20570 17222
rect 400 13862 20600 17106
rect 430 13746 20600 13862
rect 400 13526 20600 13746
rect 400 13410 20570 13526
rect 400 13190 20600 13410
rect 400 13074 20570 13190
rect 400 12854 20600 13074
rect 430 12738 20600 12854
rect 400 12518 20600 12738
rect 430 12402 20570 12518
rect 400 11510 20600 12402
rect 400 11394 20570 11510
rect 400 11174 20600 11394
rect 400 11058 20570 11174
rect 400 10502 20600 11058
rect 400 10386 20570 10502
rect 400 10166 20600 10386
rect 400 10050 20570 10166
rect 400 9494 20600 10050
rect 400 9378 20570 9494
rect 400 8822 20600 9378
rect 400 8706 20570 8822
rect 400 7814 20600 8706
rect 400 7698 20570 7814
rect 400 1554 20600 7698
<< metal4 >>
rect 2224 1538 2384 19238
rect 9904 1538 10064 19238
rect 17584 1538 17744 19238
<< obsm4 >>
rect 9254 7961 9874 11527
rect 10094 7961 10682 11527
<< labels >>
rlabel metal3 s 0 13776 400 13832 6 clk
port 1 nsew signal input
rlabel metal3 s 20600 17136 21000 17192 6 segm[0]
port 2 nsew signal output
rlabel metal2 s 12096 0 12152 400 6 segm[10]
port 3 nsew signal output
rlabel metal2 s 8736 0 8792 400 6 segm[11]
port 4 nsew signal output
rlabel metal2 s 10080 0 10136 400 6 segm[12]
port 5 nsew signal output
rlabel metal3 s 20600 12432 21000 12488 6 segm[13]
port 6 nsew signal output
rlabel metal2 s 11088 20600 11144 21000 6 segm[1]
port 7 nsew signal output
rlabel metal2 s 10416 20600 10472 21000 6 segm[2]
port 8 nsew signal output
rlabel metal3 s 20600 10416 21000 10472 6 segm[3]
port 9 nsew signal output
rlabel metal2 s 3360 0 3416 400 6 segm[4]
port 10 nsew signal output
rlabel metal2 s 9744 20600 9800 21000 6 segm[5]
port 11 nsew signal output
rlabel metal2 s 11424 0 11480 400 6 segm[6]
port 12 nsew signal output
rlabel metal3 s 20600 11424 21000 11480 6 segm[7]
port 13 nsew signal output
rlabel metal3 s 20600 13440 21000 13496 6 segm[8]
port 14 nsew signal output
rlabel metal3 s 20600 13104 21000 13160 6 segm[9]
port 15 nsew signal output
rlabel metal3 s 0 12432 400 12488 6 sel[0]
port 16 nsew signal output
rlabel metal2 s 9072 0 9128 400 6 sel[10]
port 17 nsew signal output
rlabel metal2 s 13104 0 13160 400 6 sel[11]
port 18 nsew signal output
rlabel metal2 s 8736 20600 8792 21000 6 sel[1]
port 19 nsew signal output
rlabel metal3 s 0 12768 400 12824 6 sel[2]
port 20 nsew signal output
rlabel metal3 s 20600 10080 21000 10136 6 sel[3]
port 21 nsew signal output
rlabel metal3 s 20600 11088 21000 11144 6 sel[4]
port 22 nsew signal output
rlabel metal2 s 10752 20600 10808 21000 6 sel[5]
port 23 nsew signal output
rlabel metal3 s 20600 7728 21000 7784 6 sel[6]
port 24 nsew signal output
rlabel metal3 s 20600 9408 21000 9464 6 sel[7]
port 25 nsew signal output
rlabel metal3 s 20600 8736 21000 8792 6 sel[8]
port 26 nsew signal output
rlabel metal2 s 12096 20600 12152 21000 6 sel[9]
port 27 nsew signal output
rlabel metal4 s 2224 1538 2384 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 19238 6 vss
port 29 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 21000 21000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 507566
string GDS_FILE /home/urielcho/Proyectos_caravel/ITA23_GFMPW1b/openlane/ita25/runs/23_11_10_12_47/results/signoff/ita25.magic.gds
string GDS_START 165096
<< end >>

