magic
tech gf180mcuD
magscale 1 10
timestamp 1699641913
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 18622 38274 18674 38286
rect 18622 38210 18674 38222
rect 24782 38274 24834 38286
rect 24782 38210 24834 38222
rect 22194 38110 22206 38162
rect 22258 38110 22270 38162
rect 17602 37998 17614 38050
rect 17666 37998 17678 38050
rect 23538 37998 23550 38050
rect 23602 37998 23614 38050
rect 27010 37998 27022 38050
rect 27074 37998 27086 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 19854 37490 19906 37502
rect 19854 37426 19906 37438
rect 22766 37490 22818 37502
rect 22766 37426 22818 37438
rect 26238 37490 26290 37502
rect 26238 37426 26290 37438
rect 19170 37214 19182 37266
rect 19234 37214 19246 37266
rect 22194 37214 22206 37266
rect 22258 37214 22270 37266
rect 25666 37214 25678 37266
rect 25730 37214 25742 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 22318 36706 22370 36718
rect 22318 36642 22370 36654
rect 26798 36706 26850 36718
rect 26798 36642 26850 36654
rect 21298 36430 21310 36482
rect 21362 36430 21374 36482
rect 26002 36430 26014 36482
rect 26066 36430 26078 36482
rect 25118 36370 25170 36382
rect 25118 36306 25170 36318
rect 1710 36258 1762 36270
rect 1710 36194 1762 36206
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 19170 28702 19182 28754
rect 19234 28702 19246 28754
rect 16258 28590 16270 28642
rect 16322 28590 16334 28642
rect 21422 28530 21474 28542
rect 17042 28478 17054 28530
rect 17106 28478 17118 28530
rect 21422 28466 21474 28478
rect 19630 28418 19682 28430
rect 19630 28354 19682 28366
rect 21310 28418 21362 28430
rect 21310 28354 21362 28366
rect 22654 28418 22706 28430
rect 22654 28354 22706 28366
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 17726 28082 17778 28094
rect 17726 28018 17778 28030
rect 18286 28082 18338 28094
rect 18286 28018 18338 28030
rect 18510 28082 18562 28094
rect 24446 28082 24498 28094
rect 23090 28030 23102 28082
rect 23154 28030 23166 28082
rect 18510 28018 18562 28030
rect 24446 28018 24498 28030
rect 16718 27970 16770 27982
rect 22766 27970 22818 27982
rect 20290 27918 20302 27970
rect 20354 27918 20366 27970
rect 16718 27906 16770 27918
rect 22766 27906 22818 27918
rect 23886 27970 23938 27982
rect 23886 27906 23938 27918
rect 16830 27858 16882 27870
rect 16830 27794 16882 27806
rect 17614 27858 17666 27870
rect 17614 27794 17666 27806
rect 18622 27858 18674 27870
rect 23662 27858 23714 27870
rect 19506 27806 19518 27858
rect 19570 27806 19582 27858
rect 18622 27794 18674 27806
rect 23662 27794 23714 27806
rect 23998 27858 24050 27870
rect 23998 27794 24050 27806
rect 24334 27858 24386 27870
rect 24334 27794 24386 27806
rect 22418 27694 22430 27746
rect 22482 27694 22494 27746
rect 16718 27634 16770 27646
rect 16718 27570 16770 27582
rect 17726 27634 17778 27646
rect 17726 27570 17778 27582
rect 24446 27634 24498 27646
rect 24446 27570 24498 27582
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 21646 27186 21698 27198
rect 17826 27134 17838 27186
rect 17890 27134 17902 27186
rect 23650 27134 23662 27186
rect 23714 27134 23726 27186
rect 25778 27134 25790 27186
rect 25842 27134 25854 27186
rect 21646 27122 21698 27134
rect 21422 27074 21474 27086
rect 14914 27022 14926 27074
rect 14978 27022 14990 27074
rect 21422 27010 21474 27022
rect 21758 27074 21810 27086
rect 21970 27022 21982 27074
rect 22034 27022 22046 27074
rect 22866 27022 22878 27074
rect 22930 27022 22942 27074
rect 21758 27010 21810 27022
rect 21534 26962 21586 26974
rect 15698 26910 15710 26962
rect 15762 26910 15774 26962
rect 21534 26898 21586 26910
rect 18286 26850 18338 26862
rect 18286 26786 18338 26798
rect 22542 26850 22594 26862
rect 22542 26786 22594 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 16382 26514 16434 26526
rect 23550 26514 23602 26526
rect 21746 26462 21758 26514
rect 21810 26462 21822 26514
rect 16382 26450 16434 26462
rect 23550 26450 23602 26462
rect 16606 26402 16658 26414
rect 16606 26338 16658 26350
rect 16718 26402 16770 26414
rect 16718 26338 16770 26350
rect 22654 26402 22706 26414
rect 23438 26402 23490 26414
rect 22866 26350 22878 26402
rect 22930 26399 22942 26402
rect 23202 26399 23214 26402
rect 22930 26353 23214 26399
rect 22930 26350 22942 26353
rect 23202 26350 23214 26353
rect 23266 26350 23278 26402
rect 22654 26338 22706 26350
rect 23438 26338 23490 26350
rect 22094 26290 22146 26302
rect 4274 26238 4286 26290
rect 4338 26238 4350 26290
rect 14018 26238 14030 26290
rect 14082 26238 14094 26290
rect 22094 26226 22146 26238
rect 23662 26290 23714 26302
rect 23662 26226 23714 26238
rect 24110 26290 24162 26302
rect 24110 26226 24162 26238
rect 14478 26178 14530 26190
rect 11106 26126 11118 26178
rect 11170 26126 11182 26178
rect 13234 26126 13246 26178
rect 13298 26126 13310 26178
rect 14478 26114 14530 26126
rect 20638 26178 20690 26190
rect 22754 26126 22766 26178
rect 22818 26126 22830 26178
rect 20638 26114 20690 26126
rect 1934 26066 1986 26078
rect 1934 26002 1986 26014
rect 22430 26066 22482 26078
rect 22430 26002 22482 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 14366 25618 14418 25630
rect 2034 25566 2046 25618
rect 2098 25566 2110 25618
rect 14366 25554 14418 25566
rect 15374 25618 15426 25630
rect 15374 25554 15426 25566
rect 15934 25618 15986 25630
rect 20402 25566 20414 25618
rect 20466 25566 20478 25618
rect 23874 25566 23886 25618
rect 23938 25566 23950 25618
rect 26002 25566 26014 25618
rect 26066 25566 26078 25618
rect 15934 25554 15986 25566
rect 14478 25506 14530 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 14478 25442 14530 25454
rect 14814 25506 14866 25518
rect 14814 25442 14866 25454
rect 15038 25506 15090 25518
rect 15038 25442 15090 25454
rect 15710 25506 15762 25518
rect 17490 25454 17502 25506
rect 17554 25454 17566 25506
rect 23090 25454 23102 25506
rect 23154 25454 23166 25506
rect 15710 25442 15762 25454
rect 16158 25394 16210 25406
rect 16158 25330 16210 25342
rect 16382 25394 16434 25406
rect 21870 25394 21922 25406
rect 18274 25342 18286 25394
rect 18338 25342 18350 25394
rect 16382 25330 16434 25342
rect 21870 25330 21922 25342
rect 22206 25394 22258 25406
rect 22206 25330 22258 25342
rect 22430 25394 22482 25406
rect 22430 25330 22482 25342
rect 21534 25282 21586 25294
rect 21534 25218 21586 25230
rect 22094 25282 22146 25294
rect 22094 25218 22146 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 18174 24946 18226 24958
rect 18174 24882 18226 24894
rect 25342 24946 25394 24958
rect 25342 24882 25394 24894
rect 16046 24834 16098 24846
rect 16046 24770 16098 24782
rect 18510 24834 18562 24846
rect 25230 24834 25282 24846
rect 21522 24782 21534 24834
rect 21586 24782 21598 24834
rect 18510 24770 18562 24782
rect 25230 24770 25282 24782
rect 25566 24834 25618 24846
rect 26450 24782 26462 24834
rect 26514 24782 26526 24834
rect 25566 24770 25618 24782
rect 16270 24722 16322 24734
rect 15586 24670 15598 24722
rect 15650 24670 15662 24722
rect 16270 24658 16322 24670
rect 16494 24722 16546 24734
rect 16494 24658 16546 24670
rect 17838 24722 17890 24734
rect 17838 24658 17890 24670
rect 18286 24722 18338 24734
rect 25678 24722 25730 24734
rect 19170 24670 19182 24722
rect 19234 24670 19246 24722
rect 26226 24670 26238 24722
rect 26290 24670 26302 24722
rect 37650 24670 37662 24722
rect 37714 24670 37726 24722
rect 18286 24658 18338 24670
rect 25678 24658 25730 24670
rect 16158 24610 16210 24622
rect 12786 24558 12798 24610
rect 12850 24558 12862 24610
rect 14914 24558 14926 24610
rect 14978 24558 14990 24610
rect 16158 24546 16210 24558
rect 40014 24498 40066 24510
rect 40014 24434 40066 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 15374 24162 15426 24174
rect 15374 24098 15426 24110
rect 16942 24162 16994 24174
rect 16942 24098 16994 24110
rect 15038 24050 15090 24062
rect 15038 23986 15090 23998
rect 19854 24050 19906 24062
rect 40014 24050 40066 24062
rect 22642 23998 22654 24050
rect 22706 23998 22718 24050
rect 24770 23998 24782 24050
rect 24834 23998 24846 24050
rect 19854 23986 19906 23998
rect 40014 23986 40066 23998
rect 15262 23938 15314 23950
rect 17278 23938 17330 23950
rect 15586 23886 15598 23938
rect 15650 23886 15662 23938
rect 15262 23874 15314 23886
rect 17278 23874 17330 23886
rect 19966 23938 20018 23950
rect 21858 23886 21870 23938
rect 21922 23886 21934 23938
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 19966 23874 20018 23886
rect 14926 23826 14978 23838
rect 14926 23762 14978 23774
rect 17502 23826 17554 23838
rect 17502 23762 17554 23774
rect 21310 23826 21362 23838
rect 21310 23762 21362 23774
rect 16158 23714 16210 23726
rect 16158 23650 16210 23662
rect 19742 23714 19794 23726
rect 19742 23650 19794 23662
rect 20190 23714 20242 23726
rect 20190 23650 20242 23662
rect 21422 23714 21474 23726
rect 21422 23650 21474 23662
rect 21646 23714 21698 23726
rect 21646 23650 21698 23662
rect 25230 23714 25282 23726
rect 25230 23650 25282 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 24334 23378 24386 23390
rect 24334 23314 24386 23326
rect 17490 23214 17502 23266
rect 17554 23214 17566 23266
rect 17838 23154 17890 23166
rect 11442 23102 11454 23154
rect 11506 23102 11518 23154
rect 18722 23102 18734 23154
rect 18786 23102 18798 23154
rect 19506 23102 19518 23154
rect 19570 23102 19582 23154
rect 21074 23102 21086 23154
rect 21138 23102 21150 23154
rect 25778 23102 25790 23154
rect 25842 23102 25854 23154
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 17838 23090 17890 23102
rect 14702 23042 14754 23054
rect 25454 23042 25506 23054
rect 12114 22990 12126 23042
rect 12178 22990 12190 23042
rect 14242 22990 14254 23042
rect 14306 22990 14318 23042
rect 19394 22990 19406 23042
rect 19458 22990 19470 23042
rect 21746 22990 21758 23042
rect 21810 22990 21822 23042
rect 23874 22990 23886 23042
rect 23938 22990 23950 23042
rect 26562 22990 26574 23042
rect 26626 22990 26638 23042
rect 28690 22990 28702 23042
rect 28754 22990 28766 23042
rect 14702 22978 14754 22990
rect 25454 22978 25506 22990
rect 40014 22930 40066 22942
rect 19730 22878 19742 22930
rect 19794 22878 19806 22930
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 21534 22594 21586 22606
rect 21534 22530 21586 22542
rect 26574 22594 26626 22606
rect 26574 22530 26626 22542
rect 14702 22482 14754 22494
rect 14702 22418 14754 22430
rect 16718 22482 16770 22494
rect 21758 22482 21810 22494
rect 23102 22482 23154 22494
rect 17378 22430 17390 22482
rect 17442 22430 17454 22482
rect 21970 22430 21982 22482
rect 22034 22430 22046 22482
rect 16718 22418 16770 22430
rect 21758 22418 21810 22430
rect 23102 22418 23154 22430
rect 40014 22482 40066 22494
rect 40014 22418 40066 22430
rect 14814 22370 14866 22382
rect 14814 22306 14866 22318
rect 15262 22370 15314 22382
rect 15262 22306 15314 22318
rect 15598 22370 15650 22382
rect 15598 22306 15650 22318
rect 16158 22370 16210 22382
rect 19294 22370 19346 22382
rect 17826 22318 17838 22370
rect 17890 22318 17902 22370
rect 16158 22306 16210 22318
rect 19294 22306 19346 22318
rect 19630 22370 19682 22382
rect 19630 22306 19682 22318
rect 20078 22370 20130 22382
rect 20078 22306 20130 22318
rect 20414 22370 20466 22382
rect 20414 22306 20466 22318
rect 21310 22370 21362 22382
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 21310 22306 21362 22318
rect 17278 22258 17330 22270
rect 17278 22194 17330 22206
rect 17390 22258 17442 22270
rect 17390 22194 17442 22206
rect 21982 22258 22034 22270
rect 21982 22194 22034 22206
rect 26574 22258 26626 22270
rect 26574 22194 26626 22206
rect 26686 22258 26738 22270
rect 26686 22194 26738 22206
rect 27134 22258 27186 22270
rect 27134 22194 27186 22206
rect 27358 22258 27410 22270
rect 27358 22194 27410 22206
rect 27470 22258 27522 22270
rect 27470 22194 27522 22206
rect 14590 22146 14642 22158
rect 14590 22082 14642 22094
rect 15710 22146 15762 22158
rect 15710 22082 15762 22094
rect 15934 22146 15986 22158
rect 15934 22082 15986 22094
rect 17054 22146 17106 22158
rect 17054 22082 17106 22094
rect 19406 22146 19458 22158
rect 19406 22082 19458 22094
rect 20190 22146 20242 22158
rect 20190 22082 20242 22094
rect 22206 22146 22258 22158
rect 22206 22082 22258 22094
rect 22990 22146 23042 22158
rect 22990 22082 23042 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 17390 21810 17442 21822
rect 13794 21758 13806 21810
rect 13858 21758 13870 21810
rect 17390 21746 17442 21758
rect 15374 21698 15426 21710
rect 15374 21634 15426 21646
rect 15822 21698 15874 21710
rect 17714 21646 17726 21698
rect 17778 21646 17790 21698
rect 15822 21634 15874 21646
rect 13470 21586 13522 21598
rect 18174 21586 18226 21598
rect 25342 21586 25394 21598
rect 4274 21534 4286 21586
rect 4338 21534 4350 21586
rect 16258 21534 16270 21586
rect 16322 21534 16334 21586
rect 18498 21534 18510 21586
rect 18562 21534 18574 21586
rect 25666 21534 25678 21586
rect 25730 21534 25742 21586
rect 13470 21522 13522 21534
rect 18174 21522 18226 21534
rect 25342 21522 25394 21534
rect 13134 21474 13186 21486
rect 15474 21422 15486 21474
rect 15538 21422 15550 21474
rect 16594 21422 16606 21474
rect 16658 21422 16670 21474
rect 20514 21422 20526 21474
rect 20578 21422 20590 21474
rect 26450 21422 26462 21474
rect 26514 21422 26526 21474
rect 28578 21422 28590 21474
rect 28642 21422 28654 21474
rect 13134 21410 13186 21422
rect 1934 21362 1986 21374
rect 1934 21298 1986 21310
rect 15150 21362 15202 21374
rect 15150 21298 15202 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 26350 21026 26402 21038
rect 13682 20974 13694 21026
rect 13746 20974 13758 21026
rect 17490 20974 17502 21026
rect 17554 20974 17566 21026
rect 26350 20962 26402 20974
rect 16606 20914 16658 20926
rect 9986 20862 9998 20914
rect 10050 20862 10062 20914
rect 16606 20850 16658 20862
rect 16942 20914 16994 20926
rect 16942 20850 16994 20862
rect 18286 20914 18338 20926
rect 18286 20850 18338 20862
rect 22206 20914 22258 20926
rect 22206 20850 22258 20862
rect 13918 20802 13970 20814
rect 17166 20802 17218 20814
rect 22654 20802 22706 20814
rect 12898 20750 12910 20802
rect 12962 20750 12974 20802
rect 13682 20750 13694 20802
rect 13746 20750 13758 20802
rect 16146 20750 16158 20802
rect 16210 20750 16222 20802
rect 21970 20750 21982 20802
rect 22034 20750 22046 20802
rect 13918 20738 13970 20750
rect 17166 20738 17218 20750
rect 22654 20738 22706 20750
rect 25342 20802 25394 20814
rect 25342 20738 25394 20750
rect 27358 20802 27410 20814
rect 27358 20738 27410 20750
rect 14254 20690 14306 20702
rect 12114 20638 12126 20690
rect 12178 20638 12190 20690
rect 14254 20626 14306 20638
rect 22318 20690 22370 20702
rect 22318 20626 22370 20638
rect 22990 20690 23042 20702
rect 22990 20626 23042 20638
rect 26350 20690 26402 20702
rect 26350 20626 26402 20638
rect 26462 20690 26514 20702
rect 26462 20626 26514 20638
rect 27022 20690 27074 20702
rect 27022 20626 27074 20638
rect 27246 20690 27298 20702
rect 27246 20626 27298 20638
rect 13470 20578 13522 20590
rect 13470 20514 13522 20526
rect 18398 20578 18450 20590
rect 18398 20514 18450 20526
rect 22766 20578 22818 20590
rect 25666 20526 25678 20578
rect 25730 20526 25742 20578
rect 22766 20514 22818 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 13470 20242 13522 20254
rect 13470 20178 13522 20190
rect 14030 20242 14082 20254
rect 22990 20242 23042 20254
rect 21634 20190 21646 20242
rect 21698 20190 21710 20242
rect 14030 20178 14082 20190
rect 22990 20178 23042 20190
rect 19294 20130 19346 20142
rect 20302 20130 20354 20142
rect 16146 20078 16158 20130
rect 16210 20078 16222 20130
rect 19618 20078 19630 20130
rect 19682 20078 19694 20130
rect 19954 20078 19966 20130
rect 20018 20078 20030 20130
rect 21074 20078 21086 20130
rect 21138 20078 21150 20130
rect 19294 20066 19346 20078
rect 20302 20066 20354 20078
rect 13582 20018 13634 20030
rect 22542 20018 22594 20030
rect 4274 19966 4286 20018
rect 4338 19966 4350 20018
rect 13234 19966 13246 20018
rect 13298 19966 13310 20018
rect 15922 19966 15934 20018
rect 15986 19966 15998 20018
rect 20626 19966 20638 20018
rect 20690 19966 20702 20018
rect 21522 19966 21534 20018
rect 21586 19966 21598 20018
rect 13582 19954 13634 19966
rect 22542 19954 22594 19966
rect 22766 20018 22818 20030
rect 22766 19954 22818 19966
rect 22654 19906 22706 19918
rect 22654 19842 22706 19854
rect 1934 19794 1986 19806
rect 1934 19730 1986 19742
rect 13918 19794 13970 19806
rect 13918 19730 13970 19742
rect 14254 19794 14306 19806
rect 14254 19730 14306 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 17502 19458 17554 19470
rect 17502 19394 17554 19406
rect 21422 19458 21474 19470
rect 21422 19394 21474 19406
rect 19966 19346 20018 19358
rect 40014 19346 40066 19358
rect 9986 19294 9998 19346
rect 10050 19294 10062 19346
rect 12114 19294 12126 19346
rect 12178 19294 12190 19346
rect 22530 19294 22542 19346
rect 22594 19294 22606 19346
rect 24658 19294 24670 19346
rect 24722 19294 24734 19346
rect 19966 19282 20018 19294
rect 40014 19282 40066 19294
rect 16382 19234 16434 19246
rect 12898 19182 12910 19234
rect 12962 19182 12974 19234
rect 15586 19182 15598 19234
rect 15650 19182 15662 19234
rect 16382 19170 16434 19182
rect 16494 19234 16546 19246
rect 18734 19234 18786 19246
rect 16818 19182 16830 19234
rect 16882 19182 16894 19234
rect 17154 19182 17166 19234
rect 17218 19182 17230 19234
rect 16494 19170 16546 19182
rect 18734 19170 18786 19182
rect 19742 19234 19794 19246
rect 19742 19170 19794 19182
rect 20078 19234 20130 19246
rect 27470 19234 27522 19246
rect 22082 19182 22094 19234
rect 22146 19182 22158 19234
rect 25442 19182 25454 19234
rect 25506 19182 25518 19234
rect 26898 19182 26910 19234
rect 26962 19182 26974 19234
rect 20078 19170 20130 19182
rect 27470 19170 27522 19182
rect 27694 19234 27746 19246
rect 27694 19170 27746 19182
rect 28254 19234 28306 19246
rect 28254 19170 28306 19182
rect 28366 19234 28418 19246
rect 37650 19182 37662 19234
rect 37714 19182 37726 19234
rect 28366 19170 28418 19182
rect 16270 19122 16322 19134
rect 15810 19070 15822 19122
rect 15874 19070 15886 19122
rect 16270 19058 16322 19070
rect 17838 19122 17890 19134
rect 17838 19058 17890 19070
rect 20302 19122 20354 19134
rect 20302 19058 20354 19070
rect 21534 19122 21586 19134
rect 21534 19058 21586 19070
rect 26238 19122 26290 19134
rect 26238 19058 26290 19070
rect 27246 19122 27298 19134
rect 27246 19058 27298 19070
rect 13582 19010 13634 19022
rect 13582 18946 13634 18958
rect 16606 19010 16658 19022
rect 16606 18946 16658 18958
rect 17390 19010 17442 19022
rect 19070 19010 19122 19022
rect 18162 18958 18174 19010
rect 18226 18958 18238 19010
rect 17390 18946 17442 18958
rect 19070 18946 19122 18958
rect 19294 19010 19346 19022
rect 19294 18946 19346 18958
rect 19406 19010 19458 19022
rect 19406 18946 19458 18958
rect 19854 19010 19906 19022
rect 19854 18946 19906 18958
rect 21870 19010 21922 19022
rect 21870 18946 21922 18958
rect 25902 19010 25954 19022
rect 25902 18946 25954 18958
rect 26462 19010 26514 19022
rect 26462 18946 26514 18958
rect 26574 19010 26626 19022
rect 26574 18946 26626 18958
rect 26686 19010 26738 19022
rect 26686 18946 26738 18958
rect 27582 19010 27634 19022
rect 27582 18946 27634 18958
rect 27806 19010 27858 19022
rect 27806 18946 27858 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 15822 18674 15874 18686
rect 14242 18622 14254 18674
rect 14306 18622 14318 18674
rect 15822 18610 15874 18622
rect 23102 18674 23154 18686
rect 23102 18610 23154 18622
rect 16046 18562 16098 18574
rect 19406 18562 19458 18574
rect 23326 18562 23378 18574
rect 14354 18510 14366 18562
rect 14418 18510 14430 18562
rect 16258 18510 16270 18562
rect 16322 18510 16334 18562
rect 20850 18510 20862 18562
rect 20914 18510 20926 18562
rect 21858 18510 21870 18562
rect 21922 18510 21934 18562
rect 16046 18498 16098 18510
rect 19406 18498 19458 18510
rect 23326 18498 23378 18510
rect 14926 18450 14978 18462
rect 14242 18398 14254 18450
rect 14306 18398 14318 18450
rect 14926 18386 14978 18398
rect 15374 18450 15426 18462
rect 15374 18386 15426 18398
rect 16494 18450 16546 18462
rect 19742 18450 19794 18462
rect 16594 18398 16606 18450
rect 16658 18398 16670 18450
rect 17714 18398 17726 18450
rect 17778 18398 17790 18450
rect 17938 18398 17950 18450
rect 18002 18398 18014 18450
rect 16494 18386 16546 18398
rect 19742 18386 19794 18398
rect 19966 18450 20018 18462
rect 20962 18398 20974 18450
rect 21026 18398 21038 18450
rect 21634 18398 21646 18450
rect 21698 18398 21710 18450
rect 22978 18398 22990 18450
rect 23042 18398 23054 18450
rect 23650 18398 23662 18450
rect 23714 18398 23726 18450
rect 26002 18398 26014 18450
rect 26066 18398 26078 18450
rect 26786 18398 26798 18450
rect 26850 18398 26862 18450
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 19966 18386 20018 18398
rect 16158 18338 16210 18350
rect 19518 18338 19570 18350
rect 17826 18286 17838 18338
rect 17890 18286 17902 18338
rect 16158 18274 16210 18286
rect 19518 18274 19570 18286
rect 23438 18338 23490 18350
rect 23438 18274 23490 18286
rect 25678 18338 25730 18350
rect 28914 18286 28926 18338
rect 28978 18286 28990 18338
rect 25678 18274 25730 18286
rect 15150 18226 15202 18238
rect 40014 18226 40066 18238
rect 17490 18174 17502 18226
rect 17554 18174 17566 18226
rect 15150 18162 15202 18174
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 22990 17890 23042 17902
rect 22990 17826 23042 17838
rect 15598 17778 15650 17790
rect 15598 17714 15650 17726
rect 18062 17778 18114 17790
rect 18062 17714 18114 17726
rect 21422 17778 21474 17790
rect 23314 17726 23326 17778
rect 23378 17726 23390 17778
rect 26450 17726 26462 17778
rect 26514 17726 26526 17778
rect 28578 17726 28590 17778
rect 28642 17726 28654 17778
rect 21422 17714 21474 17726
rect 20750 17666 20802 17678
rect 22654 17666 22706 17678
rect 16258 17614 16270 17666
rect 16322 17614 16334 17666
rect 19730 17614 19742 17666
rect 19794 17614 19806 17666
rect 21858 17614 21870 17666
rect 21922 17614 21934 17666
rect 20750 17602 20802 17614
rect 22654 17602 22706 17614
rect 23550 17666 23602 17678
rect 25666 17614 25678 17666
rect 25730 17614 25742 17666
rect 23550 17602 23602 17614
rect 14366 17554 14418 17566
rect 14366 17490 14418 17502
rect 16830 17554 16882 17566
rect 16830 17490 16882 17502
rect 24110 17554 24162 17566
rect 24110 17490 24162 17502
rect 14478 17442 14530 17454
rect 14478 17378 14530 17390
rect 15038 17442 15090 17454
rect 15038 17378 15090 17390
rect 16382 17442 16434 17454
rect 23214 17442 23266 17454
rect 19506 17390 19518 17442
rect 19570 17390 19582 17442
rect 20402 17390 20414 17442
rect 20466 17390 20478 17442
rect 22306 17390 22318 17442
rect 22370 17390 22382 17442
rect 16382 17378 16434 17390
rect 23214 17378 23266 17390
rect 23886 17442 23938 17454
rect 23886 17378 23938 17390
rect 24222 17442 24274 17454
rect 24222 17378 24274 17390
rect 25342 17442 25394 17454
rect 25342 17378 25394 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 15374 17106 15426 17118
rect 14466 17054 14478 17106
rect 14530 17054 14542 17106
rect 15374 17042 15426 17054
rect 27918 17106 27970 17118
rect 27918 17042 27970 17054
rect 18734 16994 18786 17006
rect 11218 16942 11230 16994
rect 11282 16942 11294 16994
rect 15698 16942 15710 16994
rect 15762 16942 15774 16994
rect 18734 16930 18786 16942
rect 28030 16994 28082 17006
rect 28030 16930 28082 16942
rect 17726 16882 17778 16894
rect 18510 16882 18562 16894
rect 10546 16830 10558 16882
rect 10610 16830 10622 16882
rect 14242 16830 14254 16882
rect 14306 16830 14318 16882
rect 16034 16830 16046 16882
rect 16098 16830 16110 16882
rect 18050 16830 18062 16882
rect 18114 16830 18126 16882
rect 19170 16830 19182 16882
rect 19234 16830 19246 16882
rect 17726 16818 17778 16830
rect 18510 16818 18562 16830
rect 13806 16770 13858 16782
rect 13346 16718 13358 16770
rect 13410 16718 13422 16770
rect 13806 16706 13858 16718
rect 16270 16770 16322 16782
rect 16270 16706 16322 16718
rect 16382 16770 16434 16782
rect 16382 16706 16434 16718
rect 18622 16770 18674 16782
rect 21858 16718 21870 16770
rect 21922 16718 21934 16770
rect 18622 16706 18674 16718
rect 18286 16658 18338 16670
rect 18286 16594 18338 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 15598 16322 15650 16334
rect 15598 16258 15650 16270
rect 17614 16322 17666 16334
rect 17614 16258 17666 16270
rect 18846 16210 18898 16222
rect 23326 16210 23378 16222
rect 20066 16158 20078 16210
rect 20130 16158 20142 16210
rect 24434 16158 24446 16210
rect 24498 16158 24510 16210
rect 26562 16158 26574 16210
rect 26626 16158 26638 16210
rect 18846 16146 18898 16158
rect 23326 16146 23378 16158
rect 14366 16098 14418 16110
rect 14130 16046 14142 16098
rect 14194 16046 14206 16098
rect 14366 16034 14418 16046
rect 17166 16098 17218 16110
rect 19854 16098 19906 16110
rect 17378 16046 17390 16098
rect 17442 16046 17454 16098
rect 17938 16046 17950 16098
rect 18002 16046 18014 16098
rect 18386 16046 18398 16098
rect 18450 16046 18462 16098
rect 19618 16046 19630 16098
rect 19682 16046 19694 16098
rect 20290 16046 20302 16098
rect 20354 16046 20366 16098
rect 23762 16046 23774 16098
rect 23826 16046 23838 16098
rect 17166 16034 17218 16046
rect 19854 16034 19906 16046
rect 12574 15986 12626 15998
rect 12574 15922 12626 15934
rect 12910 15986 12962 15998
rect 12910 15922 12962 15934
rect 13470 15986 13522 15998
rect 15486 15986 15538 15998
rect 14802 15934 14814 15986
rect 14866 15934 14878 15986
rect 13470 15922 13522 15934
rect 15486 15922 15538 15934
rect 15150 15874 15202 15886
rect 15150 15810 15202 15822
rect 17278 15874 17330 15886
rect 17278 15810 17330 15822
rect 20078 15874 20130 15886
rect 20078 15810 20130 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 24110 15538 24162 15550
rect 24110 15474 24162 15486
rect 24334 15538 24386 15550
rect 24334 15474 24386 15486
rect 19854 15426 19906 15438
rect 12338 15374 12350 15426
rect 12402 15374 12414 15426
rect 18946 15374 18958 15426
rect 19010 15374 19022 15426
rect 19854 15362 19906 15374
rect 20078 15426 20130 15438
rect 20078 15362 20130 15374
rect 22766 15426 22818 15438
rect 22766 15362 22818 15374
rect 23998 15426 24050 15438
rect 23998 15362 24050 15374
rect 22430 15314 22482 15326
rect 11666 15262 11678 15314
rect 11730 15262 11742 15314
rect 18722 15262 18734 15314
rect 18786 15262 18798 15314
rect 22430 15250 22482 15262
rect 22542 15314 22594 15326
rect 22542 15250 22594 15262
rect 22990 15314 23042 15326
rect 22990 15250 23042 15262
rect 14926 15202 14978 15214
rect 14466 15150 14478 15202
rect 14530 15150 14542 15202
rect 14926 15138 14978 15150
rect 19742 15090 19794 15102
rect 19742 15026 19794 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 17278 14754 17330 14766
rect 17278 14690 17330 14702
rect 22766 14754 22818 14766
rect 22766 14690 22818 14702
rect 17502 14642 17554 14654
rect 22542 14642 22594 14654
rect 18610 14590 18622 14642
rect 18674 14590 18686 14642
rect 20738 14590 20750 14642
rect 20802 14590 20814 14642
rect 17502 14578 17554 14590
rect 22542 14578 22594 14590
rect 23662 14642 23714 14654
rect 23662 14578 23714 14590
rect 17054 14530 17106 14542
rect 21982 14530 22034 14542
rect 17938 14478 17950 14530
rect 18002 14478 18014 14530
rect 17054 14466 17106 14478
rect 21982 14466 22034 14478
rect 22318 14530 22370 14542
rect 22318 14466 22370 14478
rect 22878 14530 22930 14542
rect 22878 14466 22930 14478
rect 23326 14530 23378 14542
rect 23326 14466 23378 14478
rect 23438 14530 23490 14542
rect 23438 14466 23490 14478
rect 23998 14530 24050 14542
rect 23998 14466 24050 14478
rect 23886 14418 23938 14430
rect 21634 14366 21646 14418
rect 21698 14366 21710 14418
rect 23886 14354 23938 14366
rect 16606 14306 16658 14318
rect 16606 14242 16658 14254
rect 22430 14306 22482 14318
rect 22430 14242 22482 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 19070 13970 19122 13982
rect 17378 13918 17390 13970
rect 17442 13918 17454 13970
rect 19070 13906 19122 13918
rect 20974 13970 21026 13982
rect 20974 13906 21026 13918
rect 15934 13858 15986 13870
rect 15934 13794 15986 13806
rect 16270 13858 16322 13870
rect 16270 13794 16322 13806
rect 19854 13858 19906 13870
rect 25230 13858 25282 13870
rect 22530 13806 22542 13858
rect 22594 13806 22606 13858
rect 19854 13794 19906 13806
rect 25230 13794 25282 13806
rect 17726 13746 17778 13758
rect 19170 13694 19182 13746
rect 19234 13694 19246 13746
rect 19618 13694 19630 13746
rect 19682 13694 19694 13746
rect 21746 13694 21758 13746
rect 21810 13694 21822 13746
rect 17726 13682 17778 13694
rect 17950 13634 18002 13646
rect 25342 13634 25394 13646
rect 24658 13582 24670 13634
rect 24722 13582 24734 13634
rect 17950 13570 18002 13582
rect 25342 13570 25394 13582
rect 25790 13634 25842 13646
rect 25790 13570 25842 13582
rect 19282 13470 19294 13522
rect 19346 13470 19358 13522
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 21422 13074 21474 13086
rect 15138 13022 15150 13074
rect 15202 13022 15214 13074
rect 17266 13022 17278 13074
rect 17330 13022 17342 13074
rect 18386 13022 18398 13074
rect 18450 13022 18462 13074
rect 20514 13022 20526 13074
rect 20578 13022 20590 13074
rect 22642 13022 22654 13074
rect 22706 13022 22718 13074
rect 24770 13022 24782 13074
rect 24834 13022 24846 13074
rect 21422 13010 21474 13022
rect 25230 12962 25282 12974
rect 14466 12910 14478 12962
rect 14530 12910 14542 12962
rect 17714 12910 17726 12962
rect 17778 12910 17790 12962
rect 21858 12910 21870 12962
rect 21922 12910 21934 12962
rect 25230 12898 25282 12910
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 17614 12402 17666 12414
rect 17614 12338 17666 12350
rect 19854 12402 19906 12414
rect 19854 12338 19906 12350
rect 19966 12290 20018 12302
rect 19966 12226 20018 12238
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 26126 5234 26178 5246
rect 26126 5170 26178 5182
rect 25554 5070 25566 5122
rect 25618 5070 25630 5122
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 20402 4286 20414 4338
rect 20466 4286 20478 4338
rect 25442 4286 25454 4338
rect 25506 4286 25518 4338
rect 21422 4114 21474 4126
rect 21422 4050 21474 4062
rect 26238 4114 26290 4126
rect 26238 4050 26290 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 18622 3666 18674 3678
rect 18622 3602 18674 3614
rect 22094 3666 22146 3678
rect 22094 3602 22146 3614
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 17714 3502 17726 3554
rect 17778 3502 17790 3554
rect 21074 3502 21086 3554
rect 21138 3502 21150 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 18622 38222 18674 38274
rect 24782 38222 24834 38274
rect 22206 38110 22258 38162
rect 17614 37998 17666 38050
rect 23550 37998 23602 38050
rect 27022 37998 27074 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 19854 37438 19906 37490
rect 22766 37438 22818 37490
rect 26238 37438 26290 37490
rect 19182 37214 19234 37266
rect 22206 37214 22258 37266
rect 25678 37214 25730 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 22318 36654 22370 36706
rect 26798 36654 26850 36706
rect 21310 36430 21362 36482
rect 26014 36430 26066 36482
rect 25118 36318 25170 36370
rect 1710 36206 1762 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19182 28702 19234 28754
rect 16270 28590 16322 28642
rect 17054 28478 17106 28530
rect 21422 28478 21474 28530
rect 19630 28366 19682 28418
rect 21310 28366 21362 28418
rect 22654 28366 22706 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 17726 28030 17778 28082
rect 18286 28030 18338 28082
rect 18510 28030 18562 28082
rect 23102 28030 23154 28082
rect 24446 28030 24498 28082
rect 16718 27918 16770 27970
rect 20302 27918 20354 27970
rect 22766 27918 22818 27970
rect 23886 27918 23938 27970
rect 16830 27806 16882 27858
rect 17614 27806 17666 27858
rect 18622 27806 18674 27858
rect 19518 27806 19570 27858
rect 23662 27806 23714 27858
rect 23998 27806 24050 27858
rect 24334 27806 24386 27858
rect 22430 27694 22482 27746
rect 16718 27582 16770 27634
rect 17726 27582 17778 27634
rect 24446 27582 24498 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 17838 27134 17890 27186
rect 21646 27134 21698 27186
rect 23662 27134 23714 27186
rect 25790 27134 25842 27186
rect 14926 27022 14978 27074
rect 21422 27022 21474 27074
rect 21758 27022 21810 27074
rect 21982 27022 22034 27074
rect 22878 27022 22930 27074
rect 15710 26910 15762 26962
rect 21534 26910 21586 26962
rect 18286 26798 18338 26850
rect 22542 26798 22594 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 16382 26462 16434 26514
rect 21758 26462 21810 26514
rect 23550 26462 23602 26514
rect 16606 26350 16658 26402
rect 16718 26350 16770 26402
rect 22654 26350 22706 26402
rect 22878 26350 22930 26402
rect 23214 26350 23266 26402
rect 23438 26350 23490 26402
rect 4286 26238 4338 26290
rect 14030 26238 14082 26290
rect 22094 26238 22146 26290
rect 23662 26238 23714 26290
rect 24110 26238 24162 26290
rect 11118 26126 11170 26178
rect 13246 26126 13298 26178
rect 14478 26126 14530 26178
rect 20638 26126 20690 26178
rect 22766 26126 22818 26178
rect 1934 26014 1986 26066
rect 22430 26014 22482 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 2046 25566 2098 25618
rect 14366 25566 14418 25618
rect 15374 25566 15426 25618
rect 15934 25566 15986 25618
rect 20414 25566 20466 25618
rect 23886 25566 23938 25618
rect 26014 25566 26066 25618
rect 4286 25454 4338 25506
rect 14478 25454 14530 25506
rect 14814 25454 14866 25506
rect 15038 25454 15090 25506
rect 15710 25454 15762 25506
rect 17502 25454 17554 25506
rect 23102 25454 23154 25506
rect 16158 25342 16210 25394
rect 16382 25342 16434 25394
rect 18286 25342 18338 25394
rect 21870 25342 21922 25394
rect 22206 25342 22258 25394
rect 22430 25342 22482 25394
rect 21534 25230 21586 25282
rect 22094 25230 22146 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 18174 24894 18226 24946
rect 25342 24894 25394 24946
rect 16046 24782 16098 24834
rect 18510 24782 18562 24834
rect 21534 24782 21586 24834
rect 25230 24782 25282 24834
rect 25566 24782 25618 24834
rect 26462 24782 26514 24834
rect 15598 24670 15650 24722
rect 16270 24670 16322 24722
rect 16494 24670 16546 24722
rect 17838 24670 17890 24722
rect 18286 24670 18338 24722
rect 19182 24670 19234 24722
rect 25678 24670 25730 24722
rect 26238 24670 26290 24722
rect 37662 24670 37714 24722
rect 12798 24558 12850 24610
rect 14926 24558 14978 24610
rect 16158 24558 16210 24610
rect 40014 24446 40066 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 15374 24110 15426 24162
rect 16942 24110 16994 24162
rect 15038 23998 15090 24050
rect 19854 23998 19906 24050
rect 22654 23998 22706 24050
rect 24782 23998 24834 24050
rect 40014 23998 40066 24050
rect 15262 23886 15314 23938
rect 15598 23886 15650 23938
rect 17278 23886 17330 23938
rect 19966 23886 20018 23938
rect 21870 23886 21922 23938
rect 37662 23886 37714 23938
rect 14926 23774 14978 23826
rect 17502 23774 17554 23826
rect 21310 23774 21362 23826
rect 16158 23662 16210 23714
rect 19742 23662 19794 23714
rect 20190 23662 20242 23714
rect 21422 23662 21474 23714
rect 21646 23662 21698 23714
rect 25230 23662 25282 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 24334 23326 24386 23378
rect 17502 23214 17554 23266
rect 11454 23102 11506 23154
rect 17838 23102 17890 23154
rect 18734 23102 18786 23154
rect 19518 23102 19570 23154
rect 21086 23102 21138 23154
rect 25790 23102 25842 23154
rect 37662 23102 37714 23154
rect 12126 22990 12178 23042
rect 14254 22990 14306 23042
rect 14702 22990 14754 23042
rect 19406 22990 19458 23042
rect 21758 22990 21810 23042
rect 23886 22990 23938 23042
rect 25454 22990 25506 23042
rect 26574 22990 26626 23042
rect 28702 22990 28754 23042
rect 19742 22878 19794 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 21534 22542 21586 22594
rect 26574 22542 26626 22594
rect 14702 22430 14754 22482
rect 16718 22430 16770 22482
rect 17390 22430 17442 22482
rect 21758 22430 21810 22482
rect 21982 22430 22034 22482
rect 23102 22430 23154 22482
rect 40014 22430 40066 22482
rect 14814 22318 14866 22370
rect 15262 22318 15314 22370
rect 15598 22318 15650 22370
rect 16158 22318 16210 22370
rect 17838 22318 17890 22370
rect 19294 22318 19346 22370
rect 19630 22318 19682 22370
rect 20078 22318 20130 22370
rect 20414 22318 20466 22370
rect 21310 22318 21362 22370
rect 37662 22318 37714 22370
rect 17278 22206 17330 22258
rect 17390 22206 17442 22258
rect 21982 22206 22034 22258
rect 26574 22206 26626 22258
rect 26686 22206 26738 22258
rect 27134 22206 27186 22258
rect 27358 22206 27410 22258
rect 27470 22206 27522 22258
rect 14590 22094 14642 22146
rect 15710 22094 15762 22146
rect 15934 22094 15986 22146
rect 17054 22094 17106 22146
rect 19406 22094 19458 22146
rect 20190 22094 20242 22146
rect 22206 22094 22258 22146
rect 22990 22094 23042 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 13806 21758 13858 21810
rect 17390 21758 17442 21810
rect 15374 21646 15426 21698
rect 15822 21646 15874 21698
rect 17726 21646 17778 21698
rect 4286 21534 4338 21586
rect 13470 21534 13522 21586
rect 16270 21534 16322 21586
rect 18174 21534 18226 21586
rect 18510 21534 18562 21586
rect 25342 21534 25394 21586
rect 25678 21534 25730 21586
rect 13134 21422 13186 21474
rect 15486 21422 15538 21474
rect 16606 21422 16658 21474
rect 20526 21422 20578 21474
rect 26462 21422 26514 21474
rect 28590 21422 28642 21474
rect 1934 21310 1986 21362
rect 15150 21310 15202 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 13694 20974 13746 21026
rect 17502 20974 17554 21026
rect 26350 20974 26402 21026
rect 9998 20862 10050 20914
rect 16606 20862 16658 20914
rect 16942 20862 16994 20914
rect 18286 20862 18338 20914
rect 22206 20862 22258 20914
rect 12910 20750 12962 20802
rect 13694 20750 13746 20802
rect 13918 20750 13970 20802
rect 16158 20750 16210 20802
rect 17166 20750 17218 20802
rect 21982 20750 22034 20802
rect 22654 20750 22706 20802
rect 25342 20750 25394 20802
rect 27358 20750 27410 20802
rect 12126 20638 12178 20690
rect 14254 20638 14306 20690
rect 22318 20638 22370 20690
rect 22990 20638 23042 20690
rect 26350 20638 26402 20690
rect 26462 20638 26514 20690
rect 27022 20638 27074 20690
rect 27246 20638 27298 20690
rect 13470 20526 13522 20578
rect 18398 20526 18450 20578
rect 22766 20526 22818 20578
rect 25678 20526 25730 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 13470 20190 13522 20242
rect 14030 20190 14082 20242
rect 21646 20190 21698 20242
rect 22990 20190 23042 20242
rect 16158 20078 16210 20130
rect 19294 20078 19346 20130
rect 19630 20078 19682 20130
rect 19966 20078 20018 20130
rect 20302 20078 20354 20130
rect 21086 20078 21138 20130
rect 4286 19966 4338 20018
rect 13246 19966 13298 20018
rect 13582 19966 13634 20018
rect 15934 19966 15986 20018
rect 20638 19966 20690 20018
rect 21534 19966 21586 20018
rect 22542 19966 22594 20018
rect 22766 19966 22818 20018
rect 22654 19854 22706 19906
rect 1934 19742 1986 19794
rect 13918 19742 13970 19794
rect 14254 19742 14306 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 17502 19406 17554 19458
rect 21422 19406 21474 19458
rect 9998 19294 10050 19346
rect 12126 19294 12178 19346
rect 19966 19294 20018 19346
rect 22542 19294 22594 19346
rect 24670 19294 24722 19346
rect 40014 19294 40066 19346
rect 12910 19182 12962 19234
rect 15598 19182 15650 19234
rect 16382 19182 16434 19234
rect 16494 19182 16546 19234
rect 16830 19182 16882 19234
rect 17166 19182 17218 19234
rect 18734 19182 18786 19234
rect 19742 19182 19794 19234
rect 20078 19182 20130 19234
rect 22094 19182 22146 19234
rect 25454 19182 25506 19234
rect 26910 19182 26962 19234
rect 27470 19182 27522 19234
rect 27694 19182 27746 19234
rect 28254 19182 28306 19234
rect 28366 19182 28418 19234
rect 37662 19182 37714 19234
rect 15822 19070 15874 19122
rect 16270 19070 16322 19122
rect 17838 19070 17890 19122
rect 20302 19070 20354 19122
rect 21534 19070 21586 19122
rect 26238 19070 26290 19122
rect 27246 19070 27298 19122
rect 13582 18958 13634 19010
rect 16606 18958 16658 19010
rect 17390 18958 17442 19010
rect 18174 18958 18226 19010
rect 19070 18958 19122 19010
rect 19294 18958 19346 19010
rect 19406 18958 19458 19010
rect 19854 18958 19906 19010
rect 21870 18958 21922 19010
rect 25902 18958 25954 19010
rect 26462 18958 26514 19010
rect 26574 18958 26626 19010
rect 26686 18958 26738 19010
rect 27582 18958 27634 19010
rect 27806 18958 27858 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 14254 18622 14306 18674
rect 15822 18622 15874 18674
rect 23102 18622 23154 18674
rect 14366 18510 14418 18562
rect 16046 18510 16098 18562
rect 16270 18510 16322 18562
rect 19406 18510 19458 18562
rect 20862 18510 20914 18562
rect 21870 18510 21922 18562
rect 23326 18510 23378 18562
rect 14254 18398 14306 18450
rect 14926 18398 14978 18450
rect 15374 18398 15426 18450
rect 16494 18398 16546 18450
rect 16606 18398 16658 18450
rect 17726 18398 17778 18450
rect 17950 18398 18002 18450
rect 19742 18398 19794 18450
rect 19966 18398 20018 18450
rect 20974 18398 21026 18450
rect 21646 18398 21698 18450
rect 22990 18398 23042 18450
rect 23662 18398 23714 18450
rect 26014 18398 26066 18450
rect 26798 18398 26850 18450
rect 37662 18398 37714 18450
rect 16158 18286 16210 18338
rect 17838 18286 17890 18338
rect 19518 18286 19570 18338
rect 23438 18286 23490 18338
rect 25678 18286 25730 18338
rect 28926 18286 28978 18338
rect 15150 18174 15202 18226
rect 17502 18174 17554 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 22990 17838 23042 17890
rect 15598 17726 15650 17778
rect 18062 17726 18114 17778
rect 21422 17726 21474 17778
rect 23326 17726 23378 17778
rect 26462 17726 26514 17778
rect 28590 17726 28642 17778
rect 16270 17614 16322 17666
rect 19742 17614 19794 17666
rect 20750 17614 20802 17666
rect 21870 17614 21922 17666
rect 22654 17614 22706 17666
rect 23550 17614 23602 17666
rect 25678 17614 25730 17666
rect 14366 17502 14418 17554
rect 16830 17502 16882 17554
rect 24110 17502 24162 17554
rect 14478 17390 14530 17442
rect 15038 17390 15090 17442
rect 16382 17390 16434 17442
rect 19518 17390 19570 17442
rect 20414 17390 20466 17442
rect 22318 17390 22370 17442
rect 23214 17390 23266 17442
rect 23886 17390 23938 17442
rect 24222 17390 24274 17442
rect 25342 17390 25394 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 14478 17054 14530 17106
rect 15374 17054 15426 17106
rect 27918 17054 27970 17106
rect 11230 16942 11282 16994
rect 15710 16942 15762 16994
rect 18734 16942 18786 16994
rect 28030 16942 28082 16994
rect 10558 16830 10610 16882
rect 14254 16830 14306 16882
rect 16046 16830 16098 16882
rect 17726 16830 17778 16882
rect 18062 16830 18114 16882
rect 18510 16830 18562 16882
rect 19182 16830 19234 16882
rect 13358 16718 13410 16770
rect 13806 16718 13858 16770
rect 16270 16718 16322 16770
rect 16382 16718 16434 16770
rect 18622 16718 18674 16770
rect 21870 16718 21922 16770
rect 18286 16606 18338 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 15598 16270 15650 16322
rect 17614 16270 17666 16322
rect 18846 16158 18898 16210
rect 20078 16158 20130 16210
rect 23326 16158 23378 16210
rect 24446 16158 24498 16210
rect 26574 16158 26626 16210
rect 14142 16046 14194 16098
rect 14366 16046 14418 16098
rect 17166 16046 17218 16098
rect 17390 16046 17442 16098
rect 17950 16046 18002 16098
rect 18398 16046 18450 16098
rect 19630 16046 19682 16098
rect 19854 16046 19906 16098
rect 20302 16046 20354 16098
rect 23774 16046 23826 16098
rect 12574 15934 12626 15986
rect 12910 15934 12962 15986
rect 13470 15934 13522 15986
rect 14814 15934 14866 15986
rect 15486 15934 15538 15986
rect 15150 15822 15202 15874
rect 17278 15822 17330 15874
rect 20078 15822 20130 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 24110 15486 24162 15538
rect 24334 15486 24386 15538
rect 12350 15374 12402 15426
rect 18958 15374 19010 15426
rect 19854 15374 19906 15426
rect 20078 15374 20130 15426
rect 22766 15374 22818 15426
rect 23998 15374 24050 15426
rect 11678 15262 11730 15314
rect 18734 15262 18786 15314
rect 22430 15262 22482 15314
rect 22542 15262 22594 15314
rect 22990 15262 23042 15314
rect 14478 15150 14530 15202
rect 14926 15150 14978 15202
rect 19742 15038 19794 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 17278 14702 17330 14754
rect 22766 14702 22818 14754
rect 17502 14590 17554 14642
rect 18622 14590 18674 14642
rect 20750 14590 20802 14642
rect 22542 14590 22594 14642
rect 23662 14590 23714 14642
rect 17054 14478 17106 14530
rect 17950 14478 18002 14530
rect 21982 14478 22034 14530
rect 22318 14478 22370 14530
rect 22878 14478 22930 14530
rect 23326 14478 23378 14530
rect 23438 14478 23490 14530
rect 23998 14478 24050 14530
rect 21646 14366 21698 14418
rect 23886 14366 23938 14418
rect 16606 14254 16658 14306
rect 22430 14254 22482 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 17390 13918 17442 13970
rect 19070 13918 19122 13970
rect 20974 13918 21026 13970
rect 15934 13806 15986 13858
rect 16270 13806 16322 13858
rect 19854 13806 19906 13858
rect 22542 13806 22594 13858
rect 25230 13806 25282 13858
rect 17726 13694 17778 13746
rect 19182 13694 19234 13746
rect 19630 13694 19682 13746
rect 21758 13694 21810 13746
rect 17950 13582 18002 13634
rect 24670 13582 24722 13634
rect 25342 13582 25394 13634
rect 25790 13582 25842 13634
rect 19294 13470 19346 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 15150 13022 15202 13074
rect 17278 13022 17330 13074
rect 18398 13022 18450 13074
rect 20526 13022 20578 13074
rect 21422 13022 21474 13074
rect 22654 13022 22706 13074
rect 24782 13022 24834 13074
rect 14478 12910 14530 12962
rect 17726 12910 17778 12962
rect 21870 12910 21922 12962
rect 25230 12910 25282 12962
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 17614 12350 17666 12402
rect 19854 12350 19906 12402
rect 19966 12238 20018 12290
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 26126 5182 26178 5234
rect 25566 5070 25618 5122
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 20414 4286 20466 4338
rect 25454 4286 25506 4338
rect 21422 4062 21474 4114
rect 26238 4062 26290 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18622 3614 18674 3666
rect 22094 3614 22146 3666
rect 25566 3614 25618 3666
rect 17726 3502 17778 3554
rect 21086 3502 21138 3554
rect 24558 3502 24610 3554
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 17472 41200 17584 42000
rect 18816 41200 18928 42000
rect 20160 41200 20272 42000
rect 21504 41200 21616 42000
rect 22176 41200 22288 42000
rect 23520 41200 23632 42000
rect 24192 41200 24304 42000
rect 24864 41200 24976 42000
rect 25536 41200 25648 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 17500 38276 17556 41200
rect 17500 38210 17556 38220
rect 18620 38276 18676 38286
rect 18620 38182 18676 38220
rect 17612 38050 17668 38062
rect 17612 37998 17614 38050
rect 17666 37998 17668 38050
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 1708 36258 1764 36270
rect 1708 36206 1710 36258
rect 1762 36206 1764 36258
rect 1708 35700 1764 36206
rect 1708 35634 1764 35644
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 17612 31948 17668 37998
rect 18844 37492 18900 41200
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 18844 37426 18900 37436
rect 19852 37492 19908 37502
rect 19852 37398 19908 37436
rect 17500 31892 17668 31948
rect 19180 37266 19236 37278
rect 19180 37214 19182 37266
rect 19234 37214 19236 37266
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 16268 28642 16324 28654
rect 16268 28590 16270 28642
rect 16322 28590 16324 28642
rect 4172 27636 4228 27646
rect 1932 26066 1988 26078
rect 1932 26014 1934 26066
rect 1986 26014 1988 26066
rect 1932 25620 1988 26014
rect 1932 25554 1988 25564
rect 2044 25618 2100 25630
rect 2044 25566 2046 25618
rect 2098 25566 2100 25618
rect 2044 24948 2100 25566
rect 2044 24882 2100 24892
rect 4172 21476 4228 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 14924 27188 14980 27198
rect 14924 27074 14980 27132
rect 16268 27188 16324 28590
rect 17052 28530 17108 28542
rect 17052 28478 17054 28530
rect 17106 28478 17108 28530
rect 16716 27972 16772 27982
rect 16716 27878 16772 27916
rect 16828 27860 16884 27870
rect 16828 27766 16884 27804
rect 16268 27122 16324 27132
rect 16716 27634 16772 27646
rect 16716 27582 16718 27634
rect 16770 27582 16772 27634
rect 14924 27022 14926 27074
rect 14978 27022 14980 27074
rect 4284 26292 4340 26302
rect 4284 26198 4340 26236
rect 14028 26290 14084 26302
rect 14028 26238 14030 26290
rect 14082 26238 14084 26290
rect 11116 26180 11172 26190
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 11116 25620 11172 26124
rect 13244 26180 13300 26190
rect 14028 26180 14084 26238
rect 14476 26180 14532 26190
rect 14028 26178 14532 26180
rect 14028 26126 14478 26178
rect 14530 26126 14532 26178
rect 14028 26124 14532 26126
rect 13244 26086 13300 26124
rect 14476 25732 14532 26124
rect 14924 25732 14980 27022
rect 15708 26964 15764 26974
rect 15708 26962 16436 26964
rect 15708 26910 15710 26962
rect 15762 26910 16436 26962
rect 15708 26908 16436 26910
rect 15708 26898 15764 26908
rect 16380 26514 16436 26908
rect 16380 26462 16382 26514
rect 16434 26462 16436 26514
rect 16380 26450 16436 26462
rect 16604 26404 16660 26414
rect 16492 26402 16660 26404
rect 16492 26350 16606 26402
rect 16658 26350 16660 26402
rect 16492 26348 16660 26350
rect 14476 25676 14980 25732
rect 11116 25554 11172 25564
rect 14364 25620 14420 25630
rect 14364 25526 14420 25564
rect 4284 25508 4340 25518
rect 4284 25414 4340 25452
rect 12796 25508 12852 25518
rect 12796 24724 12852 25452
rect 14476 25508 14532 25518
rect 14812 25508 14868 25518
rect 14476 25506 14868 25508
rect 14476 25454 14478 25506
rect 14530 25454 14814 25506
rect 14866 25454 14868 25506
rect 14476 25452 14868 25454
rect 14476 25442 14532 25452
rect 14812 25442 14868 25452
rect 14924 25284 14980 25676
rect 15932 26180 15988 26190
rect 15372 25620 15428 25630
rect 15372 25618 15764 25620
rect 15372 25566 15374 25618
rect 15426 25566 15764 25618
rect 15372 25564 15764 25566
rect 15372 25554 15428 25564
rect 14924 25218 14980 25228
rect 15036 25506 15092 25518
rect 15036 25454 15038 25506
rect 15090 25454 15092 25506
rect 12796 24610 12852 24668
rect 12796 24558 12798 24610
rect 12850 24558 12852 24610
rect 12796 24546 12852 24558
rect 14924 24610 14980 24622
rect 14924 24558 14926 24610
rect 14978 24558 14980 24610
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 14924 24052 14980 24558
rect 15036 24276 15092 25454
rect 15708 25506 15764 25564
rect 15932 25618 15988 26124
rect 16492 25620 16548 26348
rect 16604 26338 16660 26348
rect 16716 26402 16772 27582
rect 17052 27636 17108 28478
rect 17500 27972 17556 31892
rect 19180 28756 19236 37214
rect 20188 36708 20244 41200
rect 21532 37492 21588 41200
rect 22204 38162 22260 41200
rect 23548 38276 23604 41200
rect 23548 38210 23604 38220
rect 22204 38110 22206 38162
rect 22258 38110 22260 38162
rect 22204 38098 22260 38110
rect 23548 38050 23604 38062
rect 23548 37998 23550 38050
rect 23602 37998 23604 38050
rect 21532 37426 21588 37436
rect 22764 37492 22820 37502
rect 22764 37398 22820 37436
rect 20188 36642 20244 36652
rect 22204 37266 22260 37278
rect 22204 37214 22206 37266
rect 22258 37214 22260 37266
rect 21308 36482 21364 36494
rect 21308 36430 21310 36482
rect 21362 36430 21364 36482
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 21308 31948 21364 36430
rect 20412 31892 21364 31948
rect 22204 31948 22260 37214
rect 22316 36708 22372 36718
rect 22316 36614 22372 36652
rect 22204 31892 22484 31948
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 18508 28754 19236 28756
rect 18508 28702 19182 28754
rect 19234 28702 19236 28754
rect 18508 28700 19236 28702
rect 17724 28084 17780 28094
rect 18284 28084 18340 28094
rect 17724 28082 18340 28084
rect 17724 28030 17726 28082
rect 17778 28030 18286 28082
rect 18338 28030 18340 28082
rect 17724 28028 18340 28030
rect 17724 28018 17780 28028
rect 18284 28018 18340 28028
rect 18508 28082 18564 28700
rect 19180 28690 19236 28700
rect 18508 28030 18510 28082
rect 18562 28030 18564 28082
rect 18508 28018 18564 28030
rect 19628 28418 19684 28430
rect 19628 28366 19630 28418
rect 19682 28366 19684 28418
rect 17500 27748 17556 27916
rect 17500 27682 17556 27692
rect 17612 27858 17668 27870
rect 17612 27806 17614 27858
rect 17666 27806 17668 27858
rect 17052 27570 17108 27580
rect 17612 26908 17668 27806
rect 18620 27860 18676 27870
rect 18620 27766 18676 27804
rect 19516 27860 19572 27870
rect 19628 27860 19684 28366
rect 20300 28420 20356 28430
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20300 27970 20356 28364
rect 20300 27918 20302 27970
rect 20354 27918 20356 27970
rect 20300 27906 20356 27918
rect 19516 27858 19684 27860
rect 19516 27806 19518 27858
rect 19570 27806 19684 27858
rect 19516 27804 19684 27806
rect 17836 27748 17892 27758
rect 17724 27636 17780 27646
rect 17724 27542 17780 27580
rect 17836 27186 17892 27692
rect 17836 27134 17838 27186
rect 17890 27134 17892 27186
rect 17836 27122 17892 27134
rect 16716 26350 16718 26402
rect 16770 26350 16772 26402
rect 16716 26338 16772 26350
rect 17388 26852 17668 26908
rect 18284 26964 18340 26974
rect 18284 26852 18340 26908
rect 19516 26964 19572 27804
rect 19516 26898 19572 26908
rect 15932 25566 15934 25618
rect 15986 25566 15988 25618
rect 15932 25554 15988 25566
rect 16044 25564 16772 25620
rect 15708 25454 15710 25506
rect 15762 25454 15764 25506
rect 15708 25442 15764 25454
rect 15484 25284 15540 25294
rect 15484 24724 15540 25228
rect 16044 24834 16100 25564
rect 16156 25394 16212 25406
rect 16156 25342 16158 25394
rect 16210 25342 16212 25394
rect 16156 25172 16212 25342
rect 16380 25396 16436 25406
rect 16380 25394 16660 25396
rect 16380 25342 16382 25394
rect 16434 25342 16660 25394
rect 16380 25340 16660 25342
rect 16380 25330 16436 25340
rect 16156 25106 16212 25116
rect 16044 24782 16046 24834
rect 16098 24782 16100 24834
rect 16044 24770 16100 24782
rect 15596 24724 15652 24734
rect 15484 24722 15652 24724
rect 15484 24670 15598 24722
rect 15650 24670 15652 24722
rect 15484 24668 15652 24670
rect 15036 24220 15428 24276
rect 15372 24164 15428 24220
rect 15372 24070 15428 24108
rect 15036 24052 15092 24062
rect 14924 24050 15092 24052
rect 14924 23998 15038 24050
rect 15090 23998 15092 24050
rect 14924 23996 15092 23998
rect 15036 23986 15092 23996
rect 15260 23938 15316 23950
rect 15260 23886 15262 23938
rect 15314 23886 15316 23938
rect 14924 23826 14980 23838
rect 14924 23774 14926 23826
rect 14978 23774 14980 23826
rect 11452 23154 11508 23166
rect 11452 23102 11454 23154
rect 11506 23102 11508 23154
rect 11452 23044 11508 23102
rect 11452 22978 11508 22988
rect 12124 23042 12180 23054
rect 12124 22990 12126 23042
rect 12178 22990 12180 23042
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 12124 22484 12180 22990
rect 12124 22418 12180 22428
rect 13132 23044 13188 23054
rect 4284 21588 4340 21598
rect 4284 21494 4340 21532
rect 9996 21588 10052 21598
rect 4172 21410 4228 21420
rect 1932 21362 1988 21374
rect 1932 21310 1934 21362
rect 1986 21310 1988 21362
rect 1932 20916 1988 21310
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 1932 20850 1988 20860
rect 9996 20916 10052 21532
rect 9996 20822 10052 20860
rect 13132 21474 13188 22988
rect 14252 23042 14308 23054
rect 14252 22990 14254 23042
rect 14306 22990 14308 23042
rect 14140 22372 14196 22382
rect 13804 22316 14140 22372
rect 13804 21812 13860 22316
rect 14140 22306 14196 22316
rect 13804 21810 13972 21812
rect 13804 21758 13806 21810
rect 13858 21758 13972 21810
rect 13804 21756 13972 21758
rect 13804 21746 13860 21756
rect 13468 21588 13524 21598
rect 13132 21422 13134 21474
rect 13186 21422 13188 21474
rect 12908 20804 12964 20814
rect 13132 20804 13188 21422
rect 13356 21586 13524 21588
rect 13356 21534 13470 21586
rect 13522 21534 13524 21586
rect 13356 21532 13524 21534
rect 12908 20802 13188 20804
rect 12908 20750 12910 20802
rect 12962 20750 13188 20802
rect 12908 20748 13188 20750
rect 13244 20916 13300 20926
rect 12908 20738 12964 20748
rect 12124 20690 12180 20702
rect 12124 20638 12126 20690
rect 12178 20638 12180 20690
rect 12124 20580 12180 20638
rect 12124 20514 12180 20524
rect 4284 20020 4340 20030
rect 4284 19926 4340 19964
rect 9996 20020 10052 20030
rect 1932 19796 1988 19806
rect 1932 19702 1988 19740
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 9996 19348 10052 19964
rect 13244 20018 13300 20860
rect 13244 19966 13246 20018
rect 13298 19966 13300 20018
rect 13244 19954 13300 19966
rect 13356 20020 13412 21532
rect 13468 21522 13524 21532
rect 13692 21028 13748 21038
rect 13580 21026 13748 21028
rect 13580 20974 13694 21026
rect 13746 20974 13748 21026
rect 13580 20972 13748 20974
rect 13468 20580 13524 20590
rect 13468 20486 13524 20524
rect 13468 20244 13524 20254
rect 13580 20244 13636 20972
rect 13692 20962 13748 20972
rect 13468 20242 13636 20244
rect 13468 20190 13470 20242
rect 13522 20190 13636 20242
rect 13468 20188 13636 20190
rect 13692 20802 13748 20814
rect 13692 20750 13694 20802
rect 13746 20750 13748 20802
rect 13468 20178 13524 20188
rect 13580 20020 13636 20030
rect 13356 20018 13636 20020
rect 13356 19966 13582 20018
rect 13634 19966 13636 20018
rect 13356 19964 13636 19966
rect 13580 19908 13636 19964
rect 13580 19842 13636 19852
rect 9996 19254 10052 19292
rect 12124 19796 12180 19806
rect 12124 19346 12180 19740
rect 13692 19572 13748 20750
rect 13916 20804 13972 21756
rect 14252 21700 14308 22990
rect 14700 23044 14756 23054
rect 14700 22950 14756 22988
rect 14700 22484 14756 22494
rect 14700 22390 14756 22428
rect 14812 22372 14868 22382
rect 14924 22372 14980 23774
rect 15260 23828 15316 23886
rect 15372 23828 15428 23838
rect 15260 23772 15372 23828
rect 14868 22316 14980 22372
rect 15260 22370 15316 22382
rect 15260 22318 15262 22370
rect 15314 22318 15316 22370
rect 14812 22278 14868 22316
rect 14252 21634 14308 21644
rect 14588 22146 14644 22158
rect 14588 22094 14590 22146
rect 14642 22094 14644 22146
rect 14588 21588 14644 22094
rect 15260 22148 15316 22318
rect 15260 22082 15316 22092
rect 15372 21924 15428 23772
rect 15484 23380 15540 24668
rect 15596 24658 15652 24668
rect 16268 24724 16324 24734
rect 16268 24630 16324 24668
rect 16492 24722 16548 24734
rect 16492 24670 16494 24722
rect 16546 24670 16548 24722
rect 16156 24610 16212 24622
rect 16156 24558 16158 24610
rect 16210 24558 16212 24610
rect 16156 24276 16212 24558
rect 15596 24220 16212 24276
rect 15596 23938 15652 24220
rect 15596 23886 15598 23938
rect 15650 23886 15652 23938
rect 15596 23874 15652 23886
rect 15484 23314 15540 23324
rect 16156 23714 16212 23726
rect 16156 23662 16158 23714
rect 16210 23662 16212 23714
rect 16156 23380 16212 23662
rect 16156 23314 16212 23324
rect 15596 22372 15652 22382
rect 16156 22372 16212 22382
rect 15260 21868 15428 21924
rect 15484 22370 16212 22372
rect 15484 22318 15598 22370
rect 15650 22318 16158 22370
rect 16210 22318 16212 22370
rect 15484 22316 16212 22318
rect 14588 21522 14644 21532
rect 15148 21700 15204 21710
rect 15148 21362 15204 21644
rect 15148 21310 15150 21362
rect 15202 21310 15204 21362
rect 15148 20916 15204 21310
rect 15148 20850 15204 20860
rect 13916 20802 14084 20804
rect 13916 20750 13918 20802
rect 13970 20750 14084 20802
rect 13916 20748 14084 20750
rect 13916 20738 13972 20748
rect 14028 20242 14084 20748
rect 14028 20190 14030 20242
rect 14082 20190 14084 20242
rect 14028 20178 14084 20190
rect 14252 20690 14308 20702
rect 14252 20638 14254 20690
rect 14306 20638 14308 20690
rect 14252 20188 14308 20638
rect 14140 20132 14308 20188
rect 13916 19796 13972 19806
rect 13916 19702 13972 19740
rect 13692 19506 13748 19516
rect 12124 19294 12126 19346
rect 12178 19294 12180 19346
rect 12124 19282 12180 19294
rect 12908 19236 12964 19246
rect 12908 19142 12964 19180
rect 13580 19236 13636 19246
rect 13580 19010 13636 19180
rect 13580 18958 13582 19010
rect 13634 18958 13636 19010
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 11228 17444 11284 17454
rect 11228 16994 11284 17388
rect 11228 16942 11230 16994
rect 11282 16942 11284 16994
rect 11228 16930 11284 16942
rect 10556 16882 10612 16894
rect 10556 16830 10558 16882
rect 10610 16830 10612 16882
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 10556 15204 10612 16830
rect 13468 16884 13524 16894
rect 13356 16772 13412 16782
rect 13468 16772 13524 16828
rect 13356 16770 13524 16772
rect 13356 16718 13358 16770
rect 13410 16718 13524 16770
rect 13356 16716 13524 16718
rect 13580 16772 13636 18958
rect 14140 18676 14196 20132
rect 14252 20066 14308 20076
rect 15260 20132 15316 21868
rect 15372 21698 15428 21710
rect 15372 21646 15374 21698
rect 15426 21646 15428 21698
rect 15372 21252 15428 21646
rect 15484 21474 15540 22316
rect 15596 22306 15652 22316
rect 16156 22306 16212 22316
rect 15708 22146 15764 22158
rect 15708 22094 15710 22146
rect 15762 22094 15764 22146
rect 15708 21812 15764 22094
rect 15932 22148 15988 22158
rect 15932 22054 15988 22092
rect 15708 21746 15764 21756
rect 15820 22036 15876 22046
rect 15820 21698 15876 21980
rect 15820 21646 15822 21698
rect 15874 21646 15876 21698
rect 15820 21634 15876 21646
rect 15484 21422 15486 21474
rect 15538 21422 15540 21474
rect 15484 21410 15540 21422
rect 16268 21586 16324 21598
rect 16268 21534 16270 21586
rect 16322 21534 16324 21586
rect 16268 21252 16324 21534
rect 15372 21196 16324 21252
rect 15260 20066 15316 20076
rect 14252 19794 14308 19806
rect 14252 19742 14254 19794
rect 14306 19742 14308 19794
rect 14252 19236 14308 19742
rect 14252 19170 14308 19180
rect 15596 19234 15652 19246
rect 15596 19182 15598 19234
rect 15650 19182 15652 19234
rect 14252 18676 14308 18686
rect 14140 18674 14308 18676
rect 14140 18622 14254 18674
rect 14306 18622 14308 18674
rect 14140 18620 14308 18622
rect 14252 18610 14308 18620
rect 14364 18562 14420 18574
rect 14364 18510 14366 18562
rect 14418 18510 14420 18562
rect 14252 18450 14308 18462
rect 14252 18398 14254 18450
rect 14306 18398 14308 18450
rect 14252 18228 14308 18398
rect 14252 18162 14308 18172
rect 14364 18452 14420 18510
rect 14924 18452 14980 18462
rect 14364 18450 14980 18452
rect 14364 18398 14926 18450
rect 14978 18398 14980 18450
rect 14364 18396 14980 18398
rect 14364 17554 14420 18396
rect 14924 18386 14980 18396
rect 15372 18452 15428 18462
rect 15596 18452 15652 19182
rect 15820 19124 15876 21196
rect 16492 21140 16548 24670
rect 16604 23940 16660 25340
rect 16716 24948 16772 25564
rect 17276 25172 17332 25182
rect 16716 24892 16996 24948
rect 16940 24162 16996 24892
rect 16940 24110 16942 24162
rect 16994 24110 16996 24162
rect 16940 24098 16996 24110
rect 16716 23940 16772 23950
rect 16604 23884 16716 23940
rect 16716 22482 16772 23884
rect 17276 23938 17332 25116
rect 17276 23886 17278 23938
rect 17330 23886 17332 23938
rect 17276 23268 17332 23886
rect 16716 22430 16718 22482
rect 16770 22430 16772 22482
rect 16716 22418 16772 22430
rect 16940 23212 17276 23268
rect 16940 22148 16996 23212
rect 17276 23174 17332 23212
rect 17276 23044 17332 23054
rect 17164 22484 17220 22494
rect 16716 22092 16996 22148
rect 17052 22146 17108 22158
rect 17052 22094 17054 22146
rect 17106 22094 17108 22146
rect 16268 21084 16548 21140
rect 16604 21474 16660 21486
rect 16604 21422 16606 21474
rect 16658 21422 16660 21474
rect 16156 20916 16212 20926
rect 15932 20804 15988 20814
rect 15932 20020 15988 20748
rect 16156 20802 16212 20860
rect 16156 20750 16158 20802
rect 16210 20750 16212 20802
rect 16156 20738 16212 20750
rect 16156 20132 16212 20142
rect 16156 20038 16212 20076
rect 15932 20018 16100 20020
rect 15932 19966 15934 20018
rect 15986 19966 16100 20018
rect 15932 19964 16100 19966
rect 15932 19954 15988 19964
rect 15932 19124 15988 19134
rect 15820 19122 15932 19124
rect 15820 19070 15822 19122
rect 15874 19070 15932 19122
rect 15820 19068 15932 19070
rect 15820 19058 15876 19068
rect 15820 18900 15876 18910
rect 15820 18674 15876 18844
rect 15820 18622 15822 18674
rect 15874 18622 15876 18674
rect 15820 18610 15876 18622
rect 15932 18564 15988 19068
rect 16044 18788 16100 19964
rect 16268 19908 16324 21084
rect 16156 19852 16324 19908
rect 16604 20914 16660 21422
rect 16604 20862 16606 20914
rect 16658 20862 16660 20914
rect 16156 18900 16212 19852
rect 16604 19460 16660 20862
rect 16604 19394 16660 19404
rect 16380 19348 16436 19358
rect 16380 19234 16436 19292
rect 16380 19182 16382 19234
rect 16434 19182 16436 19234
rect 16380 19170 16436 19182
rect 16492 19236 16548 19274
rect 16492 19170 16548 19180
rect 16268 19122 16324 19134
rect 16268 19070 16270 19122
rect 16322 19070 16324 19122
rect 16268 19012 16324 19070
rect 16492 19012 16548 19022
rect 16268 18956 16492 19012
rect 16492 18946 16548 18956
rect 16604 19010 16660 19022
rect 16604 18958 16606 19010
rect 16658 18958 16660 19010
rect 16156 18844 16436 18900
rect 16044 18732 16324 18788
rect 16044 18564 16100 18574
rect 15932 18562 16100 18564
rect 15932 18510 16046 18562
rect 16098 18510 16100 18562
rect 15932 18508 16100 18510
rect 16044 18498 16100 18508
rect 16268 18562 16324 18732
rect 16268 18510 16270 18562
rect 16322 18510 16324 18562
rect 15372 18450 15652 18452
rect 15372 18398 15374 18450
rect 15426 18398 15652 18450
rect 15372 18396 15652 18398
rect 15372 18386 15428 18396
rect 15036 18228 15092 18238
rect 15148 18228 15204 18238
rect 15092 18226 15204 18228
rect 15092 18174 15150 18226
rect 15202 18174 15204 18226
rect 15092 18172 15204 18174
rect 14364 17502 14366 17554
rect 14418 17502 14420 17554
rect 14364 17108 14420 17502
rect 14476 17892 14532 17902
rect 14476 17444 14532 17836
rect 14476 17350 14532 17388
rect 15036 17442 15092 18172
rect 15148 18162 15204 18172
rect 15596 18116 15652 18396
rect 16156 18340 16212 18350
rect 16156 18246 16212 18284
rect 15596 18050 15652 18060
rect 15596 17780 15652 17790
rect 15596 17686 15652 17724
rect 16268 17780 16324 18510
rect 16268 17666 16324 17724
rect 16268 17614 16270 17666
rect 16322 17614 16324 17666
rect 16268 17602 16324 17614
rect 15036 17390 15038 17442
rect 15090 17390 15092 17442
rect 14476 17108 14532 17118
rect 14364 17052 14476 17108
rect 14476 17014 14532 17052
rect 14252 16884 14308 16894
rect 14140 16828 14252 16884
rect 13804 16772 13860 16782
rect 13580 16770 13860 16772
rect 13580 16718 13806 16770
rect 13858 16718 13860 16770
rect 13580 16716 13860 16718
rect 13356 16706 13412 16716
rect 12572 16100 12628 16110
rect 12572 15988 12628 16044
rect 12348 15986 12628 15988
rect 12348 15934 12574 15986
rect 12626 15934 12628 15986
rect 12348 15932 12628 15934
rect 12348 15426 12404 15932
rect 12572 15922 12628 15932
rect 12908 15988 12964 15998
rect 13468 15988 13524 15998
rect 12908 15986 13524 15988
rect 12908 15934 12910 15986
rect 12962 15934 13470 15986
rect 13522 15934 13524 15986
rect 12908 15932 13524 15934
rect 12908 15922 12964 15932
rect 13468 15922 13524 15932
rect 12348 15374 12350 15426
rect 12402 15374 12404 15426
rect 12348 15362 12404 15374
rect 10556 15138 10612 15148
rect 11676 15314 11732 15326
rect 11676 15262 11678 15314
rect 11730 15262 11732 15314
rect 11676 15204 11732 15262
rect 11676 15138 11732 15148
rect 13804 15204 13860 16716
rect 14140 16098 14196 16828
rect 14252 16790 14308 16828
rect 14140 16046 14142 16098
rect 14194 16046 14196 16098
rect 14140 16034 14196 16046
rect 14364 16100 14420 16110
rect 15036 16100 15092 17390
rect 16380 17444 16436 18844
rect 16604 18676 16660 18958
rect 16716 18900 16772 22092
rect 16940 21924 16996 21934
rect 16828 21868 16940 21924
rect 16828 20916 16884 21868
rect 16940 21858 16996 21868
rect 17052 21364 17108 22094
rect 17164 21924 17220 22428
rect 17276 22258 17332 22988
rect 17388 22482 17444 26852
rect 18172 26850 18340 26852
rect 18172 26798 18286 26850
rect 18338 26798 18340 26850
rect 18172 26796 18340 26798
rect 17500 25506 17556 25518
rect 17500 25454 17502 25506
rect 17554 25454 17556 25506
rect 17500 25284 17556 25454
rect 17500 25218 17556 25228
rect 18172 25284 18228 26796
rect 18284 26758 18340 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20412 25618 20468 31892
rect 21420 28532 21476 28542
rect 21420 28530 21700 28532
rect 21420 28478 21422 28530
rect 21474 28478 21700 28530
rect 21420 28476 21700 28478
rect 21420 28466 21476 28476
rect 21308 28420 21364 28430
rect 21308 28326 21364 28364
rect 21644 27186 21700 28476
rect 21644 27134 21646 27186
rect 21698 27134 21700 27186
rect 21644 27122 21700 27134
rect 21756 27972 21812 27982
rect 21420 27074 21476 27086
rect 21420 27022 21422 27074
rect 21474 27022 21476 27074
rect 20412 25566 20414 25618
rect 20466 25566 20468 25618
rect 18172 25218 18228 25228
rect 18284 25394 18340 25406
rect 18284 25342 18286 25394
rect 18338 25342 18340 25394
rect 18172 24948 18228 24958
rect 18284 24948 18340 25342
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 18172 24946 18340 24948
rect 18172 24894 18174 24946
rect 18226 24894 18340 24946
rect 18172 24892 18340 24894
rect 19068 24892 19908 24948
rect 18172 24882 18228 24892
rect 18508 24836 18564 24846
rect 19068 24836 19124 24892
rect 18508 24834 19124 24836
rect 18508 24782 18510 24834
rect 18562 24782 19124 24834
rect 18508 24780 19124 24782
rect 18508 24770 18564 24780
rect 17836 24724 17892 24734
rect 17612 24722 17892 24724
rect 17612 24670 17838 24722
rect 17890 24670 17892 24722
rect 17612 24668 17892 24670
rect 17612 24164 17668 24668
rect 17836 24658 17892 24668
rect 18284 24722 18340 24734
rect 18284 24670 18286 24722
rect 18338 24670 18340 24722
rect 17500 23826 17556 23838
rect 17500 23774 17502 23826
rect 17554 23774 17556 23826
rect 17500 23266 17556 23774
rect 17500 23214 17502 23266
rect 17554 23214 17556 23266
rect 17500 23044 17556 23214
rect 17500 22978 17556 22988
rect 17388 22430 17390 22482
rect 17442 22430 17444 22482
rect 17388 22418 17444 22430
rect 17276 22206 17278 22258
rect 17330 22206 17332 22258
rect 17276 22194 17332 22206
rect 17388 22258 17444 22270
rect 17388 22206 17390 22258
rect 17442 22206 17444 22258
rect 17388 22036 17444 22206
rect 17612 22036 17668 24108
rect 18284 23716 18340 24670
rect 18284 23650 18340 23660
rect 19180 24722 19236 24734
rect 19180 24670 19182 24722
rect 19234 24670 19236 24722
rect 18732 23268 18788 23278
rect 17836 23156 17892 23166
rect 17836 23154 18116 23156
rect 17836 23102 17838 23154
rect 17890 23102 18116 23154
rect 17836 23100 18116 23102
rect 17836 23090 17892 23100
rect 17444 21980 17668 22036
rect 17836 22370 17892 22382
rect 17836 22318 17838 22370
rect 17890 22318 17892 22370
rect 17388 21970 17444 21980
rect 17164 21858 17220 21868
rect 17388 21812 17444 21822
rect 17444 21756 17556 21812
rect 17388 21718 17444 21756
rect 17052 21308 17332 21364
rect 16940 20916 16996 20926
rect 16828 20914 16996 20916
rect 16828 20862 16942 20914
rect 16994 20862 16996 20914
rect 16828 20860 16996 20862
rect 16828 19348 16884 19358
rect 16828 19234 16884 19292
rect 16828 19182 16830 19234
rect 16882 19182 16884 19234
rect 16828 19170 16884 19182
rect 16716 18834 16772 18844
rect 16604 18610 16660 18620
rect 16492 18452 16548 18462
rect 16492 17668 16548 18396
rect 16604 18450 16660 18462
rect 16604 18398 16606 18450
rect 16658 18398 16660 18450
rect 16604 17892 16660 18398
rect 16604 17826 16660 17836
rect 16492 17612 16884 17668
rect 16828 17554 16884 17612
rect 16828 17502 16830 17554
rect 16882 17502 16884 17554
rect 16828 17490 16884 17502
rect 16380 17350 16436 17388
rect 15372 17108 15428 17118
rect 15372 17014 15428 17052
rect 15596 16996 15652 17006
rect 15596 16322 15652 16940
rect 15708 16994 15764 17006
rect 15708 16942 15710 16994
rect 15762 16942 15764 16994
rect 15708 16660 15764 16942
rect 16380 16996 16436 17006
rect 16044 16884 16100 16922
rect 16044 16818 16100 16828
rect 16268 16772 16324 16782
rect 16268 16678 16324 16716
rect 16380 16770 16436 16940
rect 16380 16718 16382 16770
rect 16434 16718 16436 16770
rect 16380 16706 16436 16718
rect 15708 16594 15764 16604
rect 16940 16660 16996 20860
rect 17164 20804 17220 20814
rect 17164 20710 17220 20748
rect 17164 19234 17220 19246
rect 17164 19182 17166 19234
rect 17218 19182 17220 19234
rect 17164 17892 17220 19182
rect 17164 17826 17220 17836
rect 16940 16594 16996 16604
rect 15596 16270 15598 16322
rect 15650 16270 15652 16322
rect 15596 16258 15652 16270
rect 14364 16098 15092 16100
rect 14364 16046 14366 16098
rect 14418 16046 15092 16098
rect 14364 16044 15092 16046
rect 17164 16100 17220 16110
rect 17276 16100 17332 21308
rect 17500 21026 17556 21756
rect 17724 21698 17780 21710
rect 17724 21646 17726 21698
rect 17778 21646 17780 21698
rect 17724 21588 17780 21646
rect 17724 21522 17780 21532
rect 17500 20974 17502 21026
rect 17554 20974 17556 21026
rect 17500 20962 17556 20974
rect 17500 20132 17556 20142
rect 17500 19458 17556 20076
rect 17836 20020 17892 22318
rect 18060 21252 18116 23100
rect 18732 23154 18788 23212
rect 18732 23102 18734 23154
rect 18786 23102 18788 23154
rect 18732 23090 18788 23102
rect 18844 21924 18900 21934
rect 18172 21588 18228 21598
rect 18508 21588 18564 21598
rect 18172 21586 18564 21588
rect 18172 21534 18174 21586
rect 18226 21534 18510 21586
rect 18562 21534 18564 21586
rect 18172 21532 18564 21534
rect 18172 21476 18228 21532
rect 18508 21522 18564 21532
rect 18172 21410 18228 21420
rect 18060 21196 18340 21252
rect 18284 20916 18340 21196
rect 18284 20822 18340 20860
rect 18396 20578 18452 20590
rect 18396 20526 18398 20578
rect 18450 20526 18452 20578
rect 18396 20132 18452 20526
rect 18396 20066 18452 20076
rect 17836 19954 17892 19964
rect 18732 19908 18788 19918
rect 17612 19572 17668 19582
rect 17668 19516 17780 19572
rect 17612 19506 17668 19516
rect 17500 19406 17502 19458
rect 17554 19406 17556 19458
rect 17500 19394 17556 19406
rect 17388 19010 17444 19022
rect 17388 18958 17390 19010
rect 17442 18958 17444 19010
rect 17388 18676 17444 18958
rect 17388 18610 17444 18620
rect 17724 18450 17780 19516
rect 18508 19460 18564 19470
rect 17836 19124 17892 19134
rect 17836 19030 17892 19068
rect 18172 19010 18228 19022
rect 18172 18958 18174 19010
rect 18226 18958 18228 19010
rect 18172 18900 18228 18958
rect 18172 18834 18228 18844
rect 17724 18398 17726 18450
rect 17778 18398 17780 18450
rect 17724 18386 17780 18398
rect 17836 18452 17892 18462
rect 17612 18340 17668 18350
rect 17500 18226 17556 18238
rect 17500 18174 17502 18226
rect 17554 18174 17556 18226
rect 17220 16044 17332 16100
rect 17388 16884 17444 16894
rect 17388 16098 17444 16828
rect 17388 16046 17390 16098
rect 17442 16046 17444 16098
rect 14364 16034 14420 16044
rect 14812 15986 14868 16044
rect 17164 16006 17220 16044
rect 17388 16034 17444 16046
rect 14812 15934 14814 15986
rect 14866 15934 14868 15986
rect 14812 15922 14868 15934
rect 15484 15986 15540 15998
rect 15484 15934 15486 15986
rect 15538 15934 15540 15986
rect 15148 15876 15204 15886
rect 15484 15876 15540 15934
rect 15148 15874 15540 15876
rect 15148 15822 15150 15874
rect 15202 15822 15540 15874
rect 15148 15820 15540 15822
rect 17276 15874 17332 15886
rect 17276 15822 17278 15874
rect 17330 15822 17332 15874
rect 13804 15138 13860 15148
rect 14476 15540 14532 15550
rect 14476 15202 14532 15484
rect 15036 15540 15092 15550
rect 15148 15540 15204 15820
rect 15092 15484 15204 15540
rect 15036 15474 15092 15484
rect 14476 15150 14478 15202
rect 14530 15150 14532 15202
rect 14476 15138 14532 15150
rect 14924 15204 14980 15214
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 14476 12964 14532 12974
rect 14476 12870 14532 12908
rect 14924 12964 14980 15148
rect 17276 14754 17332 15822
rect 17500 15148 17556 18174
rect 17612 16322 17668 18284
rect 17836 18338 17892 18396
rect 17836 18286 17838 18338
rect 17890 18286 17892 18338
rect 17836 18274 17892 18286
rect 17948 18450 18004 18462
rect 17948 18398 17950 18450
rect 18002 18398 18004 18450
rect 17948 18340 18004 18398
rect 17836 16996 17892 17006
rect 17948 16996 18004 18284
rect 18060 17892 18116 17902
rect 18060 17778 18116 17836
rect 18060 17726 18062 17778
rect 18114 17726 18116 17778
rect 18060 17714 18116 17726
rect 17892 16940 18004 16996
rect 18508 17444 18564 19404
rect 18732 19234 18788 19852
rect 18732 19182 18734 19234
rect 18786 19182 18788 19234
rect 18732 19170 18788 19182
rect 18844 19012 18900 21868
rect 18956 21588 19012 21598
rect 18956 19236 19012 21532
rect 18956 19170 19012 19180
rect 19180 21476 19236 24670
rect 19852 24050 19908 24892
rect 19852 23998 19854 24050
rect 19906 23998 19908 24050
rect 19852 23986 19908 23998
rect 19964 23940 20020 23950
rect 20412 23940 20468 25566
rect 20636 26964 20692 26974
rect 20636 26178 20692 26908
rect 20636 26126 20638 26178
rect 20690 26126 20692 26178
rect 20636 25284 20692 26126
rect 20636 25218 20692 25228
rect 19964 23938 20468 23940
rect 19964 23886 19966 23938
rect 20018 23886 20468 23938
rect 19964 23884 20468 23886
rect 21308 25060 21364 25070
rect 21308 23940 21364 25004
rect 19964 23874 20020 23884
rect 21308 23826 21364 23884
rect 21308 23774 21310 23826
rect 21362 23774 21364 23826
rect 19740 23716 19796 23726
rect 19628 23714 19796 23716
rect 19628 23662 19742 23714
rect 19794 23662 19796 23714
rect 19628 23660 19796 23662
rect 19628 23268 19684 23660
rect 19740 23650 19796 23660
rect 20188 23716 20244 23726
rect 20188 23714 20356 23716
rect 20188 23662 20190 23714
rect 20242 23662 20356 23714
rect 20188 23660 20356 23662
rect 20188 23650 20244 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19740 23268 19796 23278
rect 19628 23212 19740 23268
rect 19516 23154 19572 23166
rect 19516 23102 19518 23154
rect 19570 23102 19572 23154
rect 19404 23044 19460 23054
rect 19292 22372 19348 22382
rect 19404 22372 19460 22988
rect 19292 22370 19460 22372
rect 19292 22318 19294 22370
rect 19346 22318 19460 22370
rect 19292 22316 19460 22318
rect 19292 22306 19348 22316
rect 19404 22148 19460 22158
rect 19516 22148 19572 23102
rect 19628 22370 19684 23212
rect 19740 23202 19796 23212
rect 19628 22318 19630 22370
rect 19682 22318 19684 22370
rect 19628 22306 19684 22318
rect 19740 22930 19796 22942
rect 19740 22878 19742 22930
rect 19794 22878 19796 22930
rect 19740 22372 19796 22878
rect 20188 22596 20244 22606
rect 19740 22306 19796 22316
rect 20076 22540 20188 22596
rect 20076 22370 20132 22540
rect 20188 22530 20244 22540
rect 20076 22318 20078 22370
rect 20130 22318 20132 22370
rect 20076 22306 20132 22318
rect 20300 22260 20356 23660
rect 21308 23604 21364 23774
rect 21308 23538 21364 23548
rect 21420 23716 21476 27022
rect 21756 27074 21812 27916
rect 22428 27972 22484 31892
rect 23548 28532 23604 37998
rect 24220 37492 24276 41200
rect 24892 38724 24948 41200
rect 24892 38668 25172 38724
rect 24780 38276 24836 38286
rect 24780 38182 24836 38220
rect 24220 37426 24276 37436
rect 25116 36370 25172 38668
rect 25564 36708 25620 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 27020 38050 27076 38062
rect 27020 37998 27022 38050
rect 27074 37998 27076 38050
rect 26236 37492 26292 37502
rect 26236 37398 26292 37436
rect 25676 37268 25732 37278
rect 25676 37266 25844 37268
rect 25676 37214 25678 37266
rect 25730 37214 25844 37266
rect 25676 37212 25844 37214
rect 25676 37202 25732 37212
rect 25564 36642 25620 36652
rect 25116 36318 25118 36370
rect 25170 36318 25172 36370
rect 25116 36306 25172 36318
rect 23100 28476 23604 28532
rect 21980 27860 22036 27870
rect 21980 27076 22036 27804
rect 22428 27746 22484 27916
rect 22428 27694 22430 27746
rect 22482 27694 22484 27746
rect 22428 27682 22484 27694
rect 22652 28418 22708 28430
rect 22652 28366 22654 28418
rect 22706 28366 22708 28418
rect 21756 27022 21758 27074
rect 21810 27022 21812 27074
rect 21756 27010 21812 27022
rect 21868 27074 22036 27076
rect 21868 27022 21982 27074
rect 22034 27022 22036 27074
rect 21868 27020 22036 27022
rect 21532 26964 21588 26974
rect 21868 26908 21924 27020
rect 21980 27010 22036 27020
rect 22652 26908 22708 28366
rect 23100 28082 23156 28476
rect 23100 28030 23102 28082
rect 23154 28030 23156 28082
rect 23100 28018 23156 28030
rect 24444 28084 24500 28094
rect 24444 27990 24500 28028
rect 25788 28084 25844 37212
rect 26796 36708 26852 36718
rect 26796 36614 26852 36652
rect 22764 27972 22820 27982
rect 22764 27878 22820 27916
rect 23884 27970 23940 27982
rect 23884 27918 23886 27970
rect 23938 27918 23940 27970
rect 23660 27858 23716 27870
rect 23660 27806 23662 27858
rect 23714 27806 23716 27858
rect 23660 27186 23716 27806
rect 23660 27134 23662 27186
rect 23714 27134 23716 27186
rect 23660 27122 23716 27134
rect 22876 27074 22932 27086
rect 22876 27022 22878 27074
rect 22930 27022 22932 27074
rect 22876 26908 22932 27022
rect 21532 26870 21588 26908
rect 21756 26852 21924 26908
rect 22540 26852 22932 26908
rect 22988 26964 23044 26974
rect 21756 26514 21812 26852
rect 21756 26462 21758 26514
rect 21810 26462 21812 26514
rect 21756 26450 21812 26462
rect 22540 26850 22596 26852
rect 22540 26798 22542 26850
rect 22594 26798 22596 26850
rect 22092 26292 22148 26302
rect 22092 26198 22148 26236
rect 22428 26068 22484 26078
rect 21980 26066 22484 26068
rect 21980 26014 22430 26066
rect 22482 26014 22484 26066
rect 21980 26012 22484 26014
rect 21868 25394 21924 25406
rect 21868 25342 21870 25394
rect 21922 25342 21924 25394
rect 21532 25284 21588 25294
rect 21532 24836 21588 25228
rect 21756 25060 21812 25070
rect 21868 25060 21924 25342
rect 21812 25004 21924 25060
rect 21756 24994 21812 25004
rect 21532 24834 21924 24836
rect 21532 24782 21534 24834
rect 21586 24782 21924 24834
rect 21532 24780 21924 24782
rect 21532 24770 21588 24780
rect 21084 23380 21140 23390
rect 21084 23154 21140 23324
rect 21084 23102 21086 23154
rect 21138 23102 21140 23154
rect 21084 23090 21140 23102
rect 20412 22372 20468 22382
rect 21308 22372 21364 22382
rect 20412 22370 21364 22372
rect 20412 22318 20414 22370
rect 20466 22318 21310 22370
rect 21362 22318 21364 22370
rect 20412 22316 21364 22318
rect 20412 22306 20468 22316
rect 21308 22306 21364 22316
rect 20300 22194 20356 22204
rect 19460 22092 19572 22148
rect 20188 22148 20244 22158
rect 19404 21924 19460 22092
rect 20188 22054 20244 22092
rect 21420 22036 21476 23660
rect 21532 24612 21588 24622
rect 21532 23828 21588 24556
rect 21868 23938 21924 24780
rect 21868 23886 21870 23938
rect 21922 23886 21924 23938
rect 21868 23874 21924 23886
rect 21532 22594 21588 23772
rect 21644 23716 21700 23726
rect 21644 23622 21700 23660
rect 21980 23268 22036 26012
rect 22428 26002 22484 26012
rect 22204 25394 22260 25406
rect 22204 25342 22206 25394
rect 22258 25342 22260 25394
rect 22092 25282 22148 25294
rect 22092 25230 22094 25282
rect 22146 25230 22148 25282
rect 22092 24500 22148 25230
rect 22204 24724 22260 25342
rect 22428 25394 22484 25406
rect 22428 25342 22430 25394
rect 22482 25342 22484 25394
rect 22428 24948 22484 25342
rect 22540 25284 22596 26798
rect 22652 26404 22708 26414
rect 22652 26310 22708 26348
rect 22876 26402 22932 26414
rect 22876 26350 22878 26402
rect 22930 26350 22932 26402
rect 22764 26180 22820 26190
rect 22876 26180 22932 26350
rect 22764 26178 22932 26180
rect 22764 26126 22766 26178
rect 22818 26126 22932 26178
rect 22764 26124 22932 26126
rect 22764 26114 22820 26124
rect 22540 25218 22596 25228
rect 22428 24882 22484 24892
rect 22204 24658 22260 24668
rect 22092 24444 22708 24500
rect 22652 24050 22708 24444
rect 22652 23998 22654 24050
rect 22706 23998 22708 24050
rect 22652 23986 22708 23998
rect 21980 23156 22036 23212
rect 21980 23100 22148 23156
rect 21756 23044 21812 23054
rect 21756 23042 22036 23044
rect 21756 22990 21758 23042
rect 21810 22990 22036 23042
rect 21756 22988 22036 22990
rect 21756 22978 21812 22988
rect 21532 22542 21534 22594
rect 21586 22542 21588 22594
rect 21532 22530 21588 22542
rect 21756 22484 21812 22494
rect 21756 22390 21812 22428
rect 21980 22482 22036 22988
rect 21980 22430 21982 22482
rect 22034 22430 22036 22482
rect 21980 22418 22036 22430
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 21196 21980 21476 22036
rect 21868 22372 21924 22382
rect 21868 22036 21924 22316
rect 21980 22260 22036 22270
rect 22092 22260 22148 23100
rect 22988 22372 23044 26908
rect 23548 26516 23604 26526
rect 23548 26514 23828 26516
rect 23548 26462 23550 26514
rect 23602 26462 23828 26514
rect 23548 26460 23828 26462
rect 23548 26450 23604 26460
rect 23212 26404 23268 26414
rect 23436 26404 23492 26414
rect 23212 26402 23492 26404
rect 23212 26350 23214 26402
rect 23266 26350 23438 26402
rect 23490 26350 23492 26402
rect 23212 26348 23492 26350
rect 23212 26338 23268 26348
rect 23436 26338 23492 26348
rect 23660 26290 23716 26302
rect 23660 26238 23662 26290
rect 23714 26238 23716 26290
rect 23324 25956 23380 25966
rect 23100 25506 23156 25518
rect 23100 25454 23102 25506
rect 23154 25454 23156 25506
rect 23100 25284 23156 25454
rect 23100 25218 23156 25228
rect 23212 23604 23268 23614
rect 23100 22932 23156 22942
rect 23100 22482 23156 22876
rect 23100 22430 23102 22482
rect 23154 22430 23156 22482
rect 23100 22418 23156 22430
rect 21980 22258 22148 22260
rect 21980 22206 21982 22258
rect 22034 22206 22148 22258
rect 21980 22204 22148 22206
rect 22876 22316 23044 22372
rect 21980 22194 22036 22204
rect 22204 22148 22260 22158
rect 22540 22148 22596 22158
rect 22204 22146 22540 22148
rect 22204 22094 22206 22146
rect 22258 22094 22540 22146
rect 22204 22092 22540 22094
rect 22204 22082 22260 22092
rect 22540 22082 22596 22092
rect 21868 21980 22148 22036
rect 19404 21858 19460 21868
rect 18508 17108 18564 17388
rect 17836 16930 17892 16940
rect 17724 16882 17780 16894
rect 17724 16830 17726 16882
rect 17778 16830 17780 16882
rect 17724 16772 17780 16830
rect 18060 16884 18116 16894
rect 18060 16790 18116 16828
rect 18508 16882 18564 17052
rect 18732 18956 18900 19012
rect 19068 19010 19124 19022
rect 19068 18958 19070 19010
rect 19122 18958 19124 19010
rect 18732 16996 18788 18956
rect 19068 18900 19124 18958
rect 19068 18834 19124 18844
rect 18732 16902 18788 16940
rect 18844 18228 18900 18238
rect 18508 16830 18510 16882
rect 18562 16830 18564 16882
rect 18508 16818 18564 16830
rect 17724 16706 17780 16716
rect 18396 16772 18452 16782
rect 18284 16660 18340 16670
rect 18284 16566 18340 16604
rect 17612 16270 17614 16322
rect 17666 16270 17668 16322
rect 17612 16258 17668 16270
rect 17948 16098 18004 16110
rect 17948 16046 17950 16098
rect 18002 16046 18004 16098
rect 17948 15428 18004 16046
rect 18396 16098 18452 16716
rect 18396 16046 18398 16098
rect 18450 16046 18452 16098
rect 18396 16034 18452 16046
rect 18620 16770 18676 16782
rect 18620 16718 18622 16770
rect 18674 16718 18676 16770
rect 18620 15988 18676 16718
rect 17948 15362 18004 15372
rect 18508 15932 18676 15988
rect 18732 16660 18788 16670
rect 17276 14702 17278 14754
rect 17330 14702 17332 14754
rect 17276 14690 17332 14702
rect 17388 15092 17556 15148
rect 17724 15316 17780 15326
rect 17388 14644 17444 15092
rect 17500 14644 17556 14654
rect 17388 14588 17500 14644
rect 17500 14550 17556 14588
rect 17052 14532 17108 14542
rect 17052 14530 17444 14532
rect 17052 14478 17054 14530
rect 17106 14478 17444 14530
rect 17052 14476 17444 14478
rect 17052 14466 17108 14476
rect 16604 14308 16660 14318
rect 16268 14306 16660 14308
rect 16268 14254 16606 14306
rect 16658 14254 16660 14306
rect 16268 14252 16660 14254
rect 15932 13860 15988 13870
rect 15148 13858 15988 13860
rect 15148 13806 15934 13858
rect 15986 13806 15988 13858
rect 15148 13804 15988 13806
rect 15148 13074 15204 13804
rect 15932 13794 15988 13804
rect 16268 13858 16324 14252
rect 16604 14242 16660 14252
rect 17388 13970 17444 14476
rect 17388 13918 17390 13970
rect 17442 13918 17444 13970
rect 17388 13906 17444 13918
rect 16268 13806 16270 13858
rect 16322 13806 16324 13858
rect 16268 13794 16324 13806
rect 17724 13746 17780 15260
rect 17948 14530 18004 14542
rect 17948 14478 17950 14530
rect 18002 14478 18004 14530
rect 17948 13972 18004 14478
rect 18508 14420 18564 15932
rect 18732 15316 18788 16604
rect 18844 16210 18900 18172
rect 19180 16882 19236 21420
rect 20524 21476 20580 21486
rect 20524 21382 20580 21420
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19292 20132 19348 20142
rect 19628 20132 19684 20170
rect 19348 20076 19572 20132
rect 19292 20038 19348 20076
rect 19292 19010 19348 19022
rect 19292 18958 19294 19010
rect 19346 18958 19348 19010
rect 19292 18340 19348 18958
rect 19404 19012 19460 19022
rect 19404 18918 19460 18956
rect 19404 18564 19460 18574
rect 19516 18564 19572 20076
rect 19628 20066 19684 20076
rect 19964 20130 20020 20142
rect 19964 20078 19966 20130
rect 20018 20078 20020 20130
rect 19964 19908 20020 20078
rect 20300 20132 20356 20142
rect 20300 20038 20356 20076
rect 21084 20132 21140 20142
rect 21084 20038 21140 20076
rect 20636 20020 20692 20030
rect 20636 19926 20692 19964
rect 19964 19842 20020 19852
rect 19964 19684 20020 19694
rect 19740 19460 19796 19470
rect 19740 19234 19796 19404
rect 19964 19346 20020 19628
rect 19964 19294 19966 19346
rect 20018 19294 20020 19346
rect 19964 19282 20020 19294
rect 19740 19182 19742 19234
rect 19794 19182 19796 19234
rect 19740 19170 19796 19182
rect 20076 19236 20132 19246
rect 20076 19142 20132 19180
rect 20300 19122 20356 19134
rect 20300 19070 20302 19122
rect 20354 19070 20356 19122
rect 19852 19012 19908 19022
rect 19404 18562 19572 18564
rect 19404 18510 19406 18562
rect 19458 18510 19572 18562
rect 19404 18508 19572 18510
rect 19628 19010 19908 19012
rect 19628 18958 19854 19010
rect 19906 18958 19908 19010
rect 19628 18956 19908 18958
rect 19628 18900 19684 18956
rect 19852 18946 19908 18956
rect 19404 18498 19460 18508
rect 19516 18340 19572 18350
rect 19292 18274 19348 18284
rect 19404 18338 19572 18340
rect 19404 18286 19518 18338
rect 19570 18286 19572 18338
rect 19404 18284 19572 18286
rect 19180 16830 19182 16882
rect 19234 16830 19236 16882
rect 19180 16818 19236 16830
rect 19404 16660 19460 18284
rect 19516 18274 19572 18284
rect 19516 17442 19572 17454
rect 19516 17390 19518 17442
rect 19570 17390 19572 17442
rect 19516 16996 19572 17390
rect 19516 16930 19572 16940
rect 19404 16594 19460 16604
rect 18844 16158 18846 16210
rect 18898 16158 18900 16210
rect 18844 16146 18900 16158
rect 19628 16098 19684 18844
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19740 18450 19796 18462
rect 19740 18398 19742 18450
rect 19794 18398 19796 18450
rect 19740 18340 19796 18398
rect 19964 18452 20020 18462
rect 19964 18358 20020 18396
rect 19740 18274 19796 18284
rect 19740 18116 19796 18126
rect 19740 17666 19796 18060
rect 19740 17614 19742 17666
rect 19794 17614 19796 17666
rect 19740 17602 19796 17614
rect 20300 17444 20356 19070
rect 20972 18676 21028 18686
rect 20860 18562 20916 18574
rect 20860 18510 20862 18562
rect 20914 18510 20916 18562
rect 20748 17668 20804 17678
rect 20748 17574 20804 17612
rect 20412 17444 20468 17454
rect 20860 17444 20916 18510
rect 20972 18450 21028 18620
rect 20972 18398 20974 18450
rect 21026 18398 21028 18450
rect 20972 18386 21028 18398
rect 21196 18228 21252 21980
rect 21980 20804 22036 20814
rect 21420 20802 22036 20804
rect 21420 20750 21982 20802
rect 22034 20750 22036 20802
rect 21420 20748 22036 20750
rect 21196 18162 21252 18172
rect 21308 19572 21364 19582
rect 21308 17780 21364 19516
rect 21420 19458 21476 20748
rect 21980 20738 22036 20748
rect 22092 20580 22148 21980
rect 22204 21028 22260 21038
rect 22204 20914 22260 20972
rect 22876 20916 22932 22316
rect 22988 22148 23044 22158
rect 22988 22054 23044 22092
rect 22204 20862 22206 20914
rect 22258 20862 22260 20914
rect 22204 20850 22260 20862
rect 22652 20860 22932 20916
rect 22652 20802 22708 20860
rect 22652 20750 22654 20802
rect 22706 20750 22708 20802
rect 22652 20738 22708 20750
rect 22316 20692 22372 20702
rect 22316 20690 22484 20692
rect 22316 20638 22318 20690
rect 22370 20638 22484 20690
rect 22316 20636 22484 20638
rect 22316 20626 22372 20636
rect 21980 20524 22148 20580
rect 21644 20244 21700 20254
rect 21644 20242 21812 20244
rect 21644 20190 21646 20242
rect 21698 20190 21812 20242
rect 21644 20188 21812 20190
rect 21644 20178 21700 20188
rect 21532 20018 21588 20030
rect 21532 19966 21534 20018
rect 21586 19966 21588 20018
rect 21532 19572 21588 19966
rect 21532 19506 21588 19516
rect 21420 19406 21422 19458
rect 21474 19406 21476 19458
rect 21420 18452 21476 19406
rect 21532 19124 21588 19134
rect 21532 19030 21588 19068
rect 21756 18564 21812 20188
rect 21868 19010 21924 19022
rect 21868 18958 21870 19010
rect 21922 18958 21924 19010
rect 21868 18788 21924 18958
rect 21980 18900 22036 20524
rect 22428 20132 22484 20636
rect 22764 20578 22820 20590
rect 22764 20526 22766 20578
rect 22818 20526 22820 20578
rect 22764 20468 22820 20526
rect 22092 19234 22148 19246
rect 22092 19182 22094 19234
rect 22146 19182 22148 19234
rect 22092 19124 22148 19182
rect 22092 19058 22148 19068
rect 21980 18844 22372 18900
rect 21868 18732 22260 18788
rect 21868 18564 21924 18574
rect 21756 18562 22148 18564
rect 21756 18510 21870 18562
rect 21922 18510 22148 18562
rect 21756 18508 22148 18510
rect 21868 18498 21924 18508
rect 21420 18228 21476 18396
rect 21644 18452 21700 18462
rect 21644 18358 21700 18396
rect 21420 18172 21924 18228
rect 21420 17780 21476 17790
rect 21308 17778 21476 17780
rect 21308 17726 21422 17778
rect 21474 17726 21476 17778
rect 21308 17724 21476 17726
rect 21420 17714 21476 17724
rect 21868 17666 21924 18172
rect 21868 17614 21870 17666
rect 21922 17614 21924 17666
rect 21868 17602 21924 17614
rect 20300 17442 20916 17444
rect 20300 17390 20414 17442
rect 20466 17390 20916 17442
rect 20300 17388 20916 17390
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 16046 19630 16098
rect 19682 16046 19684 16098
rect 19628 16034 19684 16046
rect 19852 17108 19908 17118
rect 19852 16098 19908 17052
rect 20412 16884 20468 17388
rect 20412 16818 20468 16828
rect 21868 16770 21924 16782
rect 21868 16718 21870 16770
rect 21922 16718 21924 16770
rect 19852 16046 19854 16098
rect 19906 16046 19908 16098
rect 19852 16034 19908 16046
rect 20076 16210 20132 16222
rect 20076 16158 20078 16210
rect 20130 16158 20132 16210
rect 20076 16100 20132 16158
rect 21868 16212 21924 16718
rect 20076 16044 20244 16100
rect 20076 15876 20132 15914
rect 20076 15810 20132 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20188 15540 20244 16044
rect 20076 15484 20244 15540
rect 20300 16098 20356 16110
rect 20300 16046 20302 16098
rect 20354 16046 20356 16098
rect 18956 15428 19012 15438
rect 18956 15334 19012 15372
rect 19852 15426 19908 15438
rect 19852 15374 19854 15426
rect 19906 15374 19908 15426
rect 18732 15222 18788 15260
rect 19740 15092 19796 15102
rect 18620 15090 19796 15092
rect 18620 15038 19742 15090
rect 19794 15038 19796 15090
rect 18620 15036 19796 15038
rect 18620 14642 18676 15036
rect 19740 15026 19796 15036
rect 18620 14590 18622 14642
rect 18674 14590 18676 14642
rect 18620 14578 18676 14590
rect 19852 14644 19908 15374
rect 20076 15426 20132 15484
rect 20076 15374 20078 15426
rect 20130 15374 20132 15426
rect 20076 15362 20132 15374
rect 20300 15428 20356 16046
rect 20300 15148 20356 15372
rect 18508 14364 19348 14420
rect 19180 14196 19236 14206
rect 19068 13972 19124 13982
rect 17724 13694 17726 13746
rect 17778 13694 17780 13746
rect 17724 13682 17780 13694
rect 17836 13916 17948 13972
rect 15148 13022 15150 13074
rect 15202 13022 15204 13074
rect 15148 13010 15204 13022
rect 17276 13074 17332 13086
rect 17276 13022 17278 13074
rect 17330 13022 17332 13074
rect 14924 12898 14980 12908
rect 17276 12180 17332 13022
rect 17724 12964 17780 12974
rect 17836 12964 17892 13916
rect 17948 13906 18004 13916
rect 18396 13970 19124 13972
rect 18396 13918 19070 13970
rect 19122 13918 19124 13970
rect 18396 13916 19124 13918
rect 17780 12908 17892 12964
rect 17948 13634 18004 13646
rect 17948 13582 17950 13634
rect 18002 13582 18004 13634
rect 17612 12404 17668 12414
rect 17724 12404 17780 12908
rect 17612 12402 17780 12404
rect 17612 12350 17614 12402
rect 17666 12350 17780 12402
rect 17612 12348 17780 12350
rect 17612 12338 17668 12348
rect 17948 12180 18004 13582
rect 18396 13074 18452 13916
rect 19068 13906 19124 13916
rect 19180 13746 19236 14140
rect 19180 13694 19182 13746
rect 19234 13694 19236 13746
rect 19180 13682 19236 13694
rect 19292 13522 19348 14364
rect 19740 14308 19796 14318
rect 19852 14308 19908 14588
rect 19796 14252 19908 14308
rect 20076 15092 20356 15148
rect 20748 15876 20804 15886
rect 20076 14308 20132 15092
rect 20748 14642 20804 15820
rect 20748 14590 20750 14642
rect 20802 14590 20804 14642
rect 20076 14252 20244 14308
rect 19740 14242 19796 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20188 13972 20244 14252
rect 19852 13916 20244 13972
rect 19852 13858 19908 13916
rect 19852 13806 19854 13858
rect 19906 13806 19908 13858
rect 19852 13794 19908 13806
rect 19292 13470 19294 13522
rect 19346 13470 19348 13522
rect 19292 13458 19348 13470
rect 19628 13746 19684 13758
rect 19628 13694 19630 13746
rect 19682 13694 19684 13746
rect 18396 13022 18398 13074
rect 18450 13022 18452 13074
rect 18396 13010 18452 13022
rect 19628 12404 19684 13694
rect 20524 13076 20580 13086
rect 20412 13074 20580 13076
rect 20412 13022 20526 13074
rect 20578 13022 20580 13074
rect 20412 13020 20580 13022
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19852 12404 19908 12414
rect 19628 12402 19908 12404
rect 19628 12350 19854 12402
rect 19906 12350 19908 12402
rect 19628 12348 19908 12350
rect 19852 12338 19908 12348
rect 19964 12292 20020 12302
rect 19964 12198 20020 12236
rect 20412 12292 20468 13020
rect 20524 13010 20580 13020
rect 17276 12124 18004 12180
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 17276 8428 17332 12124
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 17276 8372 17780 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 17500 3668 17556 3678
rect 17500 800 17556 3612
rect 17724 3554 17780 8372
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 20412 4338 20468 12236
rect 20748 8428 20804 14590
rect 21644 14644 21700 14654
rect 21644 14418 21700 14588
rect 21644 14366 21646 14418
rect 21698 14366 21700 14418
rect 21644 14354 21700 14366
rect 20972 13972 21028 13982
rect 20972 13878 21028 13916
rect 21756 13972 21812 13982
rect 21756 13748 21812 13916
rect 21868 13748 21924 16156
rect 22092 15148 22148 18508
rect 22204 18452 22260 18732
rect 22204 18116 22260 18396
rect 22204 18050 22260 18060
rect 22316 17892 22372 18844
rect 22428 18564 22484 20076
rect 22540 20412 22820 20468
rect 22540 20018 22596 20412
rect 22540 19966 22542 20018
rect 22594 19966 22596 20018
rect 22540 19684 22596 19966
rect 22764 20018 22820 20030
rect 22764 19966 22766 20018
rect 22818 19966 22820 20018
rect 22652 19908 22708 19918
rect 22652 19814 22708 19852
rect 22540 19628 22708 19684
rect 22540 19346 22596 19358
rect 22540 19294 22542 19346
rect 22594 19294 22596 19346
rect 22540 19124 22596 19294
rect 22652 19236 22708 19628
rect 22764 19572 22820 19966
rect 22764 19506 22820 19516
rect 22652 19170 22708 19180
rect 22876 19348 22932 20860
rect 22988 20692 23044 20702
rect 22988 20242 23044 20636
rect 22988 20190 22990 20242
rect 23042 20190 23044 20242
rect 22988 20178 23044 20190
rect 22540 19058 22596 19068
rect 22428 18498 22484 18508
rect 22204 17836 22372 17892
rect 22652 18340 22708 18350
rect 22204 17220 22260 17836
rect 22652 17668 22708 18284
rect 22876 17892 22932 19292
rect 23100 18676 23156 18686
rect 23100 18582 23156 18620
rect 22988 18452 23044 18462
rect 23212 18452 23268 23548
rect 23324 21028 23380 25900
rect 23660 24724 23716 26238
rect 23772 25620 23828 26460
rect 23884 26292 23940 27918
rect 23996 27858 24052 27870
rect 23996 27806 23998 27858
rect 24050 27806 24052 27858
rect 23996 27636 24052 27806
rect 24332 27860 24388 27870
rect 24332 27766 24388 27804
rect 24444 27636 24500 27646
rect 23996 27634 24500 27636
rect 23996 27582 24446 27634
rect 24498 27582 24500 27634
rect 23996 27580 24500 27582
rect 24444 27570 24500 27580
rect 25788 27186 25844 28028
rect 25788 27134 25790 27186
rect 25842 27134 25844 27186
rect 25788 27122 25844 27134
rect 26012 36482 26068 36494
rect 26012 36430 26014 36482
rect 26066 36430 26068 36482
rect 26012 26404 26068 36430
rect 24108 26292 24164 26302
rect 23884 26290 24164 26292
rect 23884 26238 24110 26290
rect 24162 26238 24164 26290
rect 23884 26236 24164 26238
rect 23884 25620 23940 25630
rect 23772 25618 23940 25620
rect 23772 25566 23886 25618
rect 23938 25566 23940 25618
rect 23772 25564 23940 25566
rect 23884 25554 23940 25564
rect 23660 22372 23716 24668
rect 24108 23716 24164 26236
rect 25228 26292 25284 26302
rect 24780 24836 24836 24846
rect 24780 24050 24836 24780
rect 25228 24834 25284 26236
rect 26012 25618 26068 26348
rect 26012 25566 26014 25618
rect 26066 25566 26068 25618
rect 26012 25554 26068 25566
rect 25340 24948 25396 24958
rect 25340 24854 25396 24892
rect 25564 24948 25620 24958
rect 25228 24782 25230 24834
rect 25282 24782 25284 24834
rect 25228 24770 25284 24782
rect 25564 24834 25620 24892
rect 25564 24782 25566 24834
rect 25618 24782 25620 24834
rect 25564 24770 25620 24782
rect 26236 24948 26292 24958
rect 25676 24724 25732 24734
rect 25676 24630 25732 24668
rect 26236 24722 26292 24892
rect 27020 24948 27076 37998
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 27020 24882 27076 24892
rect 26460 24836 26516 24846
rect 26460 24742 26516 24780
rect 26236 24670 26238 24722
rect 26290 24670 26292 24722
rect 26236 24658 26292 24670
rect 37660 24724 37716 24734
rect 37660 24630 37716 24668
rect 40012 24498 40068 24510
rect 40012 24446 40014 24498
rect 40066 24446 40068 24498
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 40012 24276 40068 24446
rect 40012 24210 40068 24220
rect 24780 23998 24782 24050
rect 24834 23998 24836 24050
rect 24780 23986 24836 23998
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 37660 23938 37716 23950
rect 37660 23886 37662 23938
rect 37714 23886 37716 23938
rect 23884 23042 23940 23054
rect 23884 22990 23886 23042
rect 23938 22990 23940 23042
rect 23884 22932 23940 22990
rect 23884 22866 23940 22876
rect 23660 22306 23716 22316
rect 23324 20962 23380 20972
rect 23324 18564 23380 18602
rect 23324 18498 23380 18508
rect 22988 18450 23268 18452
rect 22988 18398 22990 18450
rect 23042 18398 23268 18450
rect 22988 18396 23268 18398
rect 23660 18452 23716 18462
rect 22988 18386 23044 18396
rect 23660 18358 23716 18396
rect 23436 18340 23492 18350
rect 23436 18246 23492 18284
rect 22988 17892 23044 17902
rect 22652 17574 22708 17612
rect 22764 17890 23044 17892
rect 22764 17838 22990 17890
rect 23042 17838 23044 17890
rect 22764 17836 23044 17838
rect 22316 17444 22372 17454
rect 22764 17444 22820 17836
rect 22988 17826 23044 17836
rect 23324 17780 23380 17790
rect 23324 17778 23604 17780
rect 23324 17726 23326 17778
rect 23378 17726 23604 17778
rect 23324 17724 23604 17726
rect 23324 17714 23380 17724
rect 23548 17666 23604 17724
rect 23548 17614 23550 17666
rect 23602 17614 23604 17666
rect 23548 17602 23604 17614
rect 24108 17554 24164 23660
rect 25228 23714 25284 23726
rect 25228 23662 25230 23714
rect 25282 23662 25284 23714
rect 24332 23380 24388 23390
rect 24332 23286 24388 23324
rect 25228 23380 25284 23662
rect 37660 23492 37716 23886
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 37660 23426 37716 23436
rect 25228 23044 25284 23324
rect 27356 23268 27412 23278
rect 25788 23154 25844 23166
rect 25788 23102 25790 23154
rect 25842 23102 25844 23154
rect 25452 23044 25508 23054
rect 25788 23044 25844 23102
rect 25228 23042 25844 23044
rect 25228 22990 25454 23042
rect 25506 22990 25844 23042
rect 25228 22988 25844 22990
rect 26572 23042 26628 23054
rect 26572 22990 26574 23042
rect 26626 22990 26628 23042
rect 25340 21588 25396 21598
rect 25452 21588 25508 22988
rect 26572 22594 26628 22990
rect 26572 22542 26574 22594
rect 26626 22542 26628 22594
rect 26572 22530 26628 22542
rect 26572 22260 26628 22270
rect 26572 22166 26628 22204
rect 26684 22260 26740 22270
rect 27132 22260 27188 22270
rect 26684 22258 27188 22260
rect 26684 22206 26686 22258
rect 26738 22206 27134 22258
rect 27186 22206 27188 22258
rect 26684 22204 27188 22206
rect 26684 22194 26740 22204
rect 27132 22194 27188 22204
rect 27356 22258 27412 23212
rect 28700 23268 28756 23278
rect 28700 23042 28756 23212
rect 37660 23156 37716 23166
rect 37660 23062 37716 23100
rect 28700 22990 28702 23042
rect 28754 22990 28756 23042
rect 28700 22978 28756 22990
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 37660 22370 37716 22382
rect 37660 22318 37662 22370
rect 37714 22318 37716 22370
rect 27356 22206 27358 22258
rect 27410 22206 27412 22258
rect 27356 22194 27412 22206
rect 27468 22258 27524 22270
rect 27468 22206 27470 22258
rect 27522 22206 27524 22258
rect 27244 21812 27300 21822
rect 25676 21588 25732 21598
rect 25340 21586 25732 21588
rect 25340 21534 25342 21586
rect 25394 21534 25678 21586
rect 25730 21534 25732 21586
rect 25340 21532 25732 21534
rect 25340 21522 25396 21532
rect 25676 21522 25732 21532
rect 26460 21476 26516 21486
rect 26348 21474 26516 21476
rect 26348 21422 26462 21474
rect 26514 21422 26516 21474
rect 26348 21420 26516 21422
rect 25340 21028 25396 21038
rect 25340 20802 25396 20972
rect 26348 21026 26404 21420
rect 26460 21410 26516 21420
rect 26348 20974 26350 21026
rect 26402 20974 26404 21026
rect 26348 20962 26404 20974
rect 25340 20750 25342 20802
rect 25394 20750 25396 20802
rect 25340 20738 25396 20750
rect 26348 20692 26404 20702
rect 26348 20598 26404 20636
rect 26460 20692 26516 20702
rect 27020 20692 27076 20702
rect 26460 20690 27076 20692
rect 26460 20638 26462 20690
rect 26514 20638 27022 20690
rect 27074 20638 27076 20690
rect 26460 20636 27076 20638
rect 26460 20626 26516 20636
rect 27020 20626 27076 20636
rect 27244 20690 27300 21756
rect 27244 20638 27246 20690
rect 27298 20638 27300 20690
rect 27244 20626 27300 20638
rect 27356 20804 27412 20814
rect 27468 20804 27524 22206
rect 28588 21812 28644 21822
rect 28588 21474 28644 21756
rect 37660 21812 37716 22318
rect 37660 21746 37716 21756
rect 40012 21588 40068 22430
rect 40012 21522 40068 21532
rect 28588 21422 28590 21474
rect 28642 21422 28644 21474
rect 28588 21410 28644 21422
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 27356 20802 27524 20804
rect 27356 20750 27358 20802
rect 27410 20750 27524 20802
rect 27356 20748 27524 20750
rect 25676 20580 25732 20590
rect 25676 20486 25732 20524
rect 26908 20468 26964 20478
rect 26908 20188 26964 20412
rect 27356 20188 27412 20748
rect 26908 20132 27412 20188
rect 24668 19908 24724 19918
rect 24668 19346 24724 19852
rect 24668 19294 24670 19346
rect 24722 19294 24724 19346
rect 24668 19282 24724 19294
rect 25452 19234 25508 19246
rect 25452 19182 25454 19234
rect 25506 19182 25508 19234
rect 25452 18340 25508 19182
rect 26908 19234 26964 20132
rect 26908 19182 26910 19234
rect 26962 19182 26964 19234
rect 26236 19124 26292 19134
rect 25900 19010 25956 19022
rect 25900 18958 25902 19010
rect 25954 18958 25956 19010
rect 25676 18340 25732 18350
rect 25900 18340 25956 18958
rect 26236 18676 26292 19068
rect 26460 19012 26516 19022
rect 26460 18918 26516 18956
rect 26572 19010 26628 19022
rect 26572 18958 26574 19010
rect 26626 18958 26628 19010
rect 26236 18610 26292 18620
rect 26012 18450 26068 18462
rect 26012 18398 26014 18450
rect 26066 18398 26068 18450
rect 26012 18340 26068 18398
rect 25452 18338 26068 18340
rect 25452 18286 25678 18338
rect 25730 18286 26068 18338
rect 25452 18284 26068 18286
rect 24108 17502 24110 17554
rect 24162 17502 24164 17554
rect 24108 17490 24164 17502
rect 25676 17666 25732 18284
rect 26460 17780 26516 17790
rect 26572 17780 26628 18958
rect 26460 17778 26628 17780
rect 26460 17726 26462 17778
rect 26514 17726 26628 17778
rect 26460 17724 26628 17726
rect 26684 19010 26740 19022
rect 26684 18958 26686 19010
rect 26738 18958 26740 19010
rect 26460 17714 26516 17724
rect 25676 17614 25678 17666
rect 25730 17614 25732 17666
rect 22316 17442 22820 17444
rect 22316 17390 22318 17442
rect 22370 17390 22820 17442
rect 22316 17388 22820 17390
rect 23212 17442 23268 17454
rect 23212 17390 23214 17442
rect 23266 17390 23268 17442
rect 22316 17378 22372 17388
rect 22204 17164 22932 17220
rect 22316 16548 22372 16558
rect 22316 15540 22372 16492
rect 22316 15484 22820 15540
rect 21980 15092 22036 15102
rect 22092 15092 22260 15148
rect 21980 14532 22036 15036
rect 21980 14438 22036 14476
rect 22204 14532 22260 15092
rect 22204 14466 22260 14476
rect 22316 14530 22372 15484
rect 22764 15426 22820 15484
rect 22764 15374 22766 15426
rect 22818 15374 22820 15426
rect 22764 15362 22820 15374
rect 22428 15314 22484 15326
rect 22428 15262 22430 15314
rect 22482 15262 22484 15314
rect 22428 15148 22484 15262
rect 22540 15316 22596 15326
rect 22540 15314 22708 15316
rect 22540 15262 22542 15314
rect 22594 15262 22708 15314
rect 22540 15260 22708 15262
rect 22540 15250 22596 15260
rect 22428 15092 22596 15148
rect 22540 14644 22596 15092
rect 22540 14550 22596 14588
rect 22316 14478 22318 14530
rect 22370 14478 22372 14530
rect 22316 14466 22372 14478
rect 22428 14308 22484 14318
rect 22428 14306 22596 14308
rect 22428 14254 22430 14306
rect 22482 14254 22596 14306
rect 22428 14252 22596 14254
rect 22428 14242 22484 14252
rect 22540 13858 22596 14252
rect 22540 13806 22542 13858
rect 22594 13806 22596 13858
rect 22540 13794 22596 13806
rect 21756 13746 21924 13748
rect 21756 13694 21758 13746
rect 21810 13694 21924 13746
rect 21756 13692 21924 13694
rect 21756 13682 21812 13692
rect 21420 13076 21476 13086
rect 21868 13076 21924 13692
rect 21420 13074 21924 13076
rect 21420 13022 21422 13074
rect 21474 13022 21924 13074
rect 21420 13020 21924 13022
rect 21420 13010 21476 13020
rect 21868 12964 21924 13020
rect 22652 13074 22708 15260
rect 22764 14756 22820 14766
rect 22876 14756 22932 17164
rect 22764 14754 22932 14756
rect 22764 14702 22766 14754
rect 22818 14702 22932 14754
rect 22764 14700 22932 14702
rect 22988 15314 23044 15326
rect 22988 15262 22990 15314
rect 23042 15262 23044 15314
rect 22764 14690 22820 14700
rect 22988 14644 23044 15262
rect 23212 15092 23268 17390
rect 23884 17444 23940 17454
rect 24220 17444 24276 17454
rect 25340 17444 25396 17454
rect 25676 17444 25732 17614
rect 23884 17442 24052 17444
rect 23884 17390 23886 17442
rect 23938 17390 24052 17442
rect 23884 17388 24052 17390
rect 23884 17378 23940 17388
rect 23996 16324 24052 17388
rect 24220 17442 24500 17444
rect 24220 17390 24222 17442
rect 24274 17390 24500 17442
rect 24220 17388 24500 17390
rect 24220 17378 24276 17388
rect 23996 16268 24388 16324
rect 23324 16212 23380 16222
rect 23324 16118 23380 16156
rect 23772 16212 23828 16222
rect 23772 16098 23828 16156
rect 23772 16046 23774 16098
rect 23826 16046 23828 16098
rect 23772 16034 23828 16046
rect 24108 15540 24164 15550
rect 24108 15446 24164 15484
rect 24332 15538 24388 16268
rect 24444 16210 24500 17388
rect 24444 16158 24446 16210
rect 24498 16158 24500 16210
rect 24444 16146 24500 16158
rect 25340 17442 25732 17444
rect 25340 17390 25342 17442
rect 25394 17390 25732 17442
rect 25340 17388 25732 17390
rect 25340 16212 25396 17388
rect 26684 17108 26740 18958
rect 26908 19012 26964 19182
rect 27468 19684 27524 19694
rect 27468 19234 27524 19628
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 40012 19346 40068 19358
rect 40012 19294 40014 19346
rect 40066 19294 40068 19346
rect 27468 19182 27470 19234
rect 27522 19182 27524 19234
rect 27468 19170 27524 19182
rect 27692 19236 27748 19246
rect 28252 19236 28308 19246
rect 27692 19234 28308 19236
rect 27692 19182 27694 19234
rect 27746 19182 28254 19234
rect 28306 19182 28308 19234
rect 27692 19180 28308 19182
rect 27692 19170 27748 19180
rect 28252 19170 28308 19180
rect 28364 19236 28420 19246
rect 28364 19142 28420 19180
rect 28924 19236 28980 19246
rect 27244 19124 27300 19134
rect 27244 19030 27300 19068
rect 27132 19012 27188 19022
rect 26908 18956 27132 19012
rect 27132 18946 27188 18956
rect 27580 19010 27636 19022
rect 27580 18958 27582 19010
rect 27634 18958 27636 19010
rect 26796 18564 26852 18574
rect 26796 18450 26852 18508
rect 27580 18564 27636 18958
rect 27804 19012 27860 19022
rect 27804 18918 27860 18956
rect 27580 18498 27636 18508
rect 26796 18398 26798 18450
rect 26850 18398 26852 18450
rect 26796 18386 26852 18398
rect 28588 18452 28644 18462
rect 28588 17780 28644 18396
rect 28924 18338 28980 19180
rect 37660 19236 37716 19246
rect 37660 19142 37716 19180
rect 40012 18900 40068 19294
rect 40012 18834 40068 18844
rect 37660 18452 37716 18462
rect 37660 18358 37716 18396
rect 28924 18286 28926 18338
rect 28978 18286 28980 18338
rect 28924 18274 28980 18286
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 28028 17778 28644 17780
rect 28028 17726 28590 17778
rect 28642 17726 28644 17778
rect 28028 17724 28644 17726
rect 26684 17042 26740 17052
rect 27916 17108 27972 17118
rect 27916 17014 27972 17052
rect 28028 16994 28084 17724
rect 28588 17714 28644 17724
rect 28028 16942 28030 16994
rect 28082 16942 28084 16994
rect 28028 16930 28084 16942
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 25340 16146 25396 16156
rect 25564 16212 25620 16222
rect 24332 15486 24334 15538
rect 24386 15486 24388 15538
rect 24332 15474 24388 15486
rect 25564 15540 25620 16156
rect 26572 16212 26628 16222
rect 26572 16118 26628 16156
rect 23996 15428 24052 15438
rect 23996 15334 24052 15372
rect 25564 15148 25620 15484
rect 23212 15026 23268 15036
rect 23996 15092 24052 15102
rect 22988 14578 23044 14588
rect 23660 14644 23716 14654
rect 23660 14550 23716 14588
rect 22876 14532 22932 14542
rect 22876 14438 22932 14476
rect 23324 14530 23380 14542
rect 23324 14478 23326 14530
rect 23378 14478 23380 14530
rect 23324 13860 23380 14478
rect 23436 14532 23492 14542
rect 23436 14438 23492 14476
rect 23996 14530 24052 15036
rect 23996 14478 23998 14530
rect 24050 14478 24052 14530
rect 23996 14466 24052 14478
rect 25452 15092 25620 15148
rect 23324 13794 23380 13804
rect 23884 14418 23940 14430
rect 23884 14366 23886 14418
rect 23938 14366 23940 14418
rect 22652 13022 22654 13074
rect 22706 13022 22708 13074
rect 22652 13010 22708 13022
rect 23884 13076 23940 14366
rect 25228 13860 25284 13898
rect 25228 13794 25284 13804
rect 24668 13636 24724 13646
rect 24668 13542 24724 13580
rect 25340 13636 25396 13646
rect 25340 13542 25396 13580
rect 24780 13076 24836 13086
rect 23884 13074 24836 13076
rect 23884 13022 24782 13074
rect 24834 13022 24836 13074
rect 23884 13020 24836 13022
rect 21868 12870 21924 12908
rect 24780 8428 24836 13020
rect 25228 12964 25284 13002
rect 25228 12898 25284 12908
rect 20748 8372 21140 8428
rect 20412 4286 20414 4338
rect 20466 4286 20468 4338
rect 20412 4274 20468 4286
rect 20188 4116 20244 4126
rect 18620 3668 18676 3678
rect 18620 3574 18676 3612
rect 17724 3502 17726 3554
rect 17778 3502 17780 3554
rect 17724 3490 17780 3502
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 800 20244 4060
rect 20860 3668 20916 3678
rect 20860 800 20916 3612
rect 21084 3554 21140 8372
rect 24556 8372 24836 8428
rect 21420 4116 21476 4126
rect 21420 4022 21476 4060
rect 24220 4116 24276 4126
rect 22092 3668 22148 3678
rect 22092 3574 22148 3612
rect 23548 3668 23604 3678
rect 21084 3502 21086 3554
rect 21138 3502 21140 3554
rect 21084 3490 21140 3502
rect 23548 800 23604 3612
rect 24220 800 24276 4060
rect 24556 3554 24612 8372
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 24892 5236 24948 5246
rect 24892 800 24948 5180
rect 25452 4338 25508 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 25564 13636 25620 13646
rect 25564 12740 25620 13580
rect 25788 13634 25844 13646
rect 25788 13582 25790 13634
rect 25842 13582 25844 13634
rect 25676 12964 25732 12974
rect 25788 12964 25844 13582
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 25732 12908 25844 12964
rect 25676 12898 25732 12908
rect 25564 12684 25732 12740
rect 25676 11844 25732 12684
rect 25564 11788 25732 11844
rect 35196 11788 35460 11798
rect 25564 5122 25620 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 26124 5236 26180 5246
rect 26124 5142 26180 5180
rect 25564 5070 25566 5122
rect 25618 5070 25620 5122
rect 25564 5058 25620 5070
rect 25452 4286 25454 4338
rect 25506 4286 25508 4338
rect 25452 4274 25508 4286
rect 26236 4116 26292 4126
rect 26236 4022 26292 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 17472 0 17584 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 24864 0 24976 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 17500 38220 17556 38276
rect 18620 38274 18676 38276
rect 18620 38222 18622 38274
rect 18622 38222 18674 38274
rect 18674 38222 18676 38274
rect 18620 38220 18676 38222
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 1708 35644 1764 35700
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 18844 37436 18900 37492
rect 19852 37490 19908 37492
rect 19852 37438 19854 37490
rect 19854 37438 19906 37490
rect 19906 37438 19908 37490
rect 19852 37436 19908 37438
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4172 27580 4228 27636
rect 1932 25564 1988 25620
rect 2044 24892 2100 24948
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 14924 27132 14980 27188
rect 16716 27970 16772 27972
rect 16716 27918 16718 27970
rect 16718 27918 16770 27970
rect 16770 27918 16772 27970
rect 16716 27916 16772 27918
rect 16828 27858 16884 27860
rect 16828 27806 16830 27858
rect 16830 27806 16882 27858
rect 16882 27806 16884 27858
rect 16828 27804 16884 27806
rect 16268 27132 16324 27188
rect 4284 26290 4340 26292
rect 4284 26238 4286 26290
rect 4286 26238 4338 26290
rect 4338 26238 4340 26290
rect 4284 26236 4340 26238
rect 11116 26178 11172 26180
rect 11116 26126 11118 26178
rect 11118 26126 11170 26178
rect 11170 26126 11172 26178
rect 11116 26124 11172 26126
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 13244 26178 13300 26180
rect 13244 26126 13246 26178
rect 13246 26126 13298 26178
rect 13298 26126 13300 26178
rect 13244 26124 13300 26126
rect 11116 25564 11172 25620
rect 14364 25618 14420 25620
rect 14364 25566 14366 25618
rect 14366 25566 14418 25618
rect 14418 25566 14420 25618
rect 14364 25564 14420 25566
rect 4284 25506 4340 25508
rect 4284 25454 4286 25506
rect 4286 25454 4338 25506
rect 4338 25454 4340 25506
rect 4284 25452 4340 25454
rect 12796 25452 12852 25508
rect 15932 26124 15988 26180
rect 14924 25228 14980 25284
rect 12796 24668 12852 24724
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 23548 38220 23604 38276
rect 21532 37436 21588 37492
rect 22764 37490 22820 37492
rect 22764 37438 22766 37490
rect 22766 37438 22818 37490
rect 22818 37438 22820 37490
rect 22764 37436 22820 37438
rect 20188 36652 20244 36708
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 22316 36706 22372 36708
rect 22316 36654 22318 36706
rect 22318 36654 22370 36706
rect 22370 36654 22372 36706
rect 22316 36652 22372 36654
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 17500 27916 17556 27972
rect 17500 27692 17556 27748
rect 17052 27580 17108 27636
rect 18620 27858 18676 27860
rect 18620 27806 18622 27858
rect 18622 27806 18674 27858
rect 18674 27806 18676 27858
rect 18620 27804 18676 27806
rect 20300 28364 20356 28420
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 17836 27692 17892 27748
rect 17724 27634 17780 27636
rect 17724 27582 17726 27634
rect 17726 27582 17778 27634
rect 17778 27582 17780 27634
rect 17724 27580 17780 27582
rect 18284 26908 18340 26964
rect 19516 26908 19572 26964
rect 15484 25228 15540 25284
rect 16156 25116 16212 25172
rect 15372 24162 15428 24164
rect 15372 24110 15374 24162
rect 15374 24110 15426 24162
rect 15426 24110 15428 24162
rect 15372 24108 15428 24110
rect 11452 22988 11508 23044
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 12124 22428 12180 22484
rect 13132 22988 13188 23044
rect 4284 21586 4340 21588
rect 4284 21534 4286 21586
rect 4286 21534 4338 21586
rect 4338 21534 4340 21586
rect 4284 21532 4340 21534
rect 9996 21532 10052 21588
rect 4172 21420 4228 21476
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 1932 20860 1988 20916
rect 9996 20914 10052 20916
rect 9996 20862 9998 20914
rect 9998 20862 10050 20914
rect 10050 20862 10052 20914
rect 9996 20860 10052 20862
rect 14140 22316 14196 22372
rect 13244 20860 13300 20916
rect 12124 20524 12180 20580
rect 4284 20018 4340 20020
rect 4284 19966 4286 20018
rect 4286 19966 4338 20018
rect 4338 19966 4340 20018
rect 4284 19964 4340 19966
rect 9996 19964 10052 20020
rect 1932 19794 1988 19796
rect 1932 19742 1934 19794
rect 1934 19742 1986 19794
rect 1986 19742 1988 19794
rect 1932 19740 1988 19742
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 13468 20578 13524 20580
rect 13468 20526 13470 20578
rect 13470 20526 13522 20578
rect 13522 20526 13524 20578
rect 13468 20524 13524 20526
rect 13580 19852 13636 19908
rect 9996 19346 10052 19348
rect 9996 19294 9998 19346
rect 9998 19294 10050 19346
rect 10050 19294 10052 19346
rect 9996 19292 10052 19294
rect 12124 19740 12180 19796
rect 14700 23042 14756 23044
rect 14700 22990 14702 23042
rect 14702 22990 14754 23042
rect 14754 22990 14756 23042
rect 14700 22988 14756 22990
rect 14700 22482 14756 22484
rect 14700 22430 14702 22482
rect 14702 22430 14754 22482
rect 14754 22430 14756 22482
rect 14700 22428 14756 22430
rect 15372 23772 15428 23828
rect 14812 22370 14868 22372
rect 14812 22318 14814 22370
rect 14814 22318 14866 22370
rect 14866 22318 14868 22370
rect 14812 22316 14868 22318
rect 14252 21644 14308 21700
rect 15260 22092 15316 22148
rect 16268 24722 16324 24724
rect 16268 24670 16270 24722
rect 16270 24670 16322 24722
rect 16322 24670 16324 24722
rect 16268 24668 16324 24670
rect 15484 23324 15540 23380
rect 16156 23324 16212 23380
rect 14588 21532 14644 21588
rect 15148 21644 15204 21700
rect 15148 20860 15204 20916
rect 13916 19794 13972 19796
rect 13916 19742 13918 19794
rect 13918 19742 13970 19794
rect 13970 19742 13972 19794
rect 13916 19740 13972 19742
rect 13692 19516 13748 19572
rect 12908 19234 12964 19236
rect 12908 19182 12910 19234
rect 12910 19182 12962 19234
rect 12962 19182 12964 19234
rect 12908 19180 12964 19182
rect 13580 19180 13636 19236
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 11228 17388 11284 17444
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 13468 16828 13524 16884
rect 14252 20076 14308 20132
rect 15932 22146 15988 22148
rect 15932 22094 15934 22146
rect 15934 22094 15986 22146
rect 15986 22094 15988 22146
rect 15932 22092 15988 22094
rect 15708 21756 15764 21812
rect 15820 21980 15876 22036
rect 15260 20076 15316 20132
rect 14252 19180 14308 19236
rect 14252 18172 14308 18228
rect 17276 25116 17332 25172
rect 16716 23884 16772 23940
rect 17276 23212 17332 23268
rect 17276 22988 17332 23044
rect 17164 22428 17220 22484
rect 16156 20860 16212 20916
rect 15932 20748 15988 20804
rect 16156 20130 16212 20132
rect 16156 20078 16158 20130
rect 16158 20078 16210 20130
rect 16210 20078 16212 20130
rect 16156 20076 16212 20078
rect 15932 19068 15988 19124
rect 15820 18844 15876 18900
rect 16604 19404 16660 19460
rect 16380 19292 16436 19348
rect 16492 19234 16548 19236
rect 16492 19182 16494 19234
rect 16494 19182 16546 19234
rect 16546 19182 16548 19234
rect 16492 19180 16548 19182
rect 16492 18956 16548 19012
rect 15036 18172 15092 18228
rect 14476 17836 14532 17892
rect 14476 17442 14532 17444
rect 14476 17390 14478 17442
rect 14478 17390 14530 17442
rect 14530 17390 14532 17442
rect 14476 17388 14532 17390
rect 16156 18338 16212 18340
rect 16156 18286 16158 18338
rect 16158 18286 16210 18338
rect 16210 18286 16212 18338
rect 16156 18284 16212 18286
rect 15596 18060 15652 18116
rect 15596 17778 15652 17780
rect 15596 17726 15598 17778
rect 15598 17726 15650 17778
rect 15650 17726 15652 17778
rect 15596 17724 15652 17726
rect 16268 17724 16324 17780
rect 14476 17106 14532 17108
rect 14476 17054 14478 17106
rect 14478 17054 14530 17106
rect 14530 17054 14532 17106
rect 14476 17052 14532 17054
rect 14252 16882 14308 16884
rect 14252 16830 14254 16882
rect 14254 16830 14306 16882
rect 14306 16830 14308 16882
rect 14252 16828 14308 16830
rect 12572 16044 12628 16100
rect 10556 15148 10612 15204
rect 11676 15148 11732 15204
rect 16940 21868 16996 21924
rect 17500 25228 17556 25284
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 21308 28418 21364 28420
rect 21308 28366 21310 28418
rect 21310 28366 21362 28418
rect 21362 28366 21364 28418
rect 21308 28364 21364 28366
rect 21756 27916 21812 27972
rect 18172 25228 18228 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 17612 24108 17668 24164
rect 17500 22988 17556 23044
rect 18284 23660 18340 23716
rect 18732 23212 18788 23268
rect 17388 21980 17444 22036
rect 17164 21868 17220 21924
rect 17388 21810 17444 21812
rect 17388 21758 17390 21810
rect 17390 21758 17442 21810
rect 17442 21758 17444 21810
rect 17388 21756 17444 21758
rect 16828 19292 16884 19348
rect 16716 18844 16772 18900
rect 16604 18620 16660 18676
rect 16492 18450 16548 18452
rect 16492 18398 16494 18450
rect 16494 18398 16546 18450
rect 16546 18398 16548 18450
rect 16492 18396 16548 18398
rect 16604 17836 16660 17892
rect 16380 17442 16436 17444
rect 16380 17390 16382 17442
rect 16382 17390 16434 17442
rect 16434 17390 16436 17442
rect 16380 17388 16436 17390
rect 15372 17106 15428 17108
rect 15372 17054 15374 17106
rect 15374 17054 15426 17106
rect 15426 17054 15428 17106
rect 15372 17052 15428 17054
rect 15596 16940 15652 16996
rect 16380 16940 16436 16996
rect 16044 16882 16100 16884
rect 16044 16830 16046 16882
rect 16046 16830 16098 16882
rect 16098 16830 16100 16882
rect 16044 16828 16100 16830
rect 16268 16770 16324 16772
rect 16268 16718 16270 16770
rect 16270 16718 16322 16770
rect 16322 16718 16324 16770
rect 16268 16716 16324 16718
rect 15708 16604 15764 16660
rect 17164 20802 17220 20804
rect 17164 20750 17166 20802
rect 17166 20750 17218 20802
rect 17218 20750 17220 20802
rect 17164 20748 17220 20750
rect 17164 17836 17220 17892
rect 16940 16604 16996 16660
rect 17724 21532 17780 21588
rect 17500 20076 17556 20132
rect 18844 21868 18900 21924
rect 18172 21420 18228 21476
rect 18284 20914 18340 20916
rect 18284 20862 18286 20914
rect 18286 20862 18338 20914
rect 18338 20862 18340 20914
rect 18284 20860 18340 20862
rect 18396 20076 18452 20132
rect 17836 19964 17892 20020
rect 18732 19852 18788 19908
rect 17612 19516 17668 19572
rect 17388 18620 17444 18676
rect 18508 19404 18564 19460
rect 17836 19122 17892 19124
rect 17836 19070 17838 19122
rect 17838 19070 17890 19122
rect 17890 19070 17892 19122
rect 17836 19068 17892 19070
rect 18172 18844 18228 18900
rect 17836 18396 17892 18452
rect 17612 18284 17668 18340
rect 17164 16098 17220 16100
rect 17164 16046 17166 16098
rect 17166 16046 17218 16098
rect 17218 16046 17220 16098
rect 17164 16044 17220 16046
rect 17388 16828 17444 16884
rect 13804 15148 13860 15204
rect 14476 15484 14532 15540
rect 15036 15484 15092 15540
rect 14924 15202 14980 15204
rect 14924 15150 14926 15202
rect 14926 15150 14978 15202
rect 14978 15150 14980 15202
rect 14924 15148 14980 15150
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 14476 12962 14532 12964
rect 14476 12910 14478 12962
rect 14478 12910 14530 12962
rect 14530 12910 14532 12962
rect 14476 12908 14532 12910
rect 17948 18284 18004 18340
rect 18060 17836 18116 17892
rect 17836 16940 17892 16996
rect 18956 21532 19012 21588
rect 18956 19180 19012 19236
rect 20636 26908 20692 26964
rect 20636 25228 20692 25284
rect 21308 25004 21364 25060
rect 21308 23884 21364 23940
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19740 23212 19796 23268
rect 19404 23042 19460 23044
rect 19404 22990 19406 23042
rect 19406 22990 19458 23042
rect 19458 22990 19460 23042
rect 19404 22988 19460 22990
rect 19740 22316 19796 22372
rect 20188 22540 20244 22596
rect 21308 23548 21364 23604
rect 24780 38274 24836 38276
rect 24780 38222 24782 38274
rect 24782 38222 24834 38274
rect 24834 38222 24836 38274
rect 24780 38220 24836 38222
rect 24220 37436 24276 37492
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 26236 37490 26292 37492
rect 26236 37438 26238 37490
rect 26238 37438 26290 37490
rect 26290 37438 26292 37490
rect 26236 37436 26292 37438
rect 25564 36652 25620 36708
rect 22428 27916 22484 27972
rect 21980 27804 22036 27860
rect 21532 26962 21588 26964
rect 21532 26910 21534 26962
rect 21534 26910 21586 26962
rect 21586 26910 21588 26962
rect 21532 26908 21588 26910
rect 24444 28082 24500 28084
rect 24444 28030 24446 28082
rect 24446 28030 24498 28082
rect 24498 28030 24500 28082
rect 24444 28028 24500 28030
rect 26796 36706 26852 36708
rect 26796 36654 26798 36706
rect 26798 36654 26850 36706
rect 26850 36654 26852 36706
rect 26796 36652 26852 36654
rect 25788 28028 25844 28084
rect 22764 27970 22820 27972
rect 22764 27918 22766 27970
rect 22766 27918 22818 27970
rect 22818 27918 22820 27970
rect 22764 27916 22820 27918
rect 22988 26908 23044 26964
rect 22092 26290 22148 26292
rect 22092 26238 22094 26290
rect 22094 26238 22146 26290
rect 22146 26238 22148 26290
rect 22092 26236 22148 26238
rect 21532 25282 21588 25284
rect 21532 25230 21534 25282
rect 21534 25230 21586 25282
rect 21586 25230 21588 25282
rect 21532 25228 21588 25230
rect 21756 25004 21812 25060
rect 21420 23714 21476 23716
rect 21420 23662 21422 23714
rect 21422 23662 21474 23714
rect 21474 23662 21476 23714
rect 21420 23660 21476 23662
rect 21084 23324 21140 23380
rect 20300 22204 20356 22260
rect 19404 22146 19460 22148
rect 19404 22094 19406 22146
rect 19406 22094 19458 22146
rect 19458 22094 19460 22146
rect 19404 22092 19460 22094
rect 20188 22146 20244 22148
rect 20188 22094 20190 22146
rect 20190 22094 20242 22146
rect 20242 22094 20244 22146
rect 20188 22092 20244 22094
rect 21532 24556 21588 24612
rect 21532 23772 21588 23828
rect 21644 23714 21700 23716
rect 21644 23662 21646 23714
rect 21646 23662 21698 23714
rect 21698 23662 21700 23714
rect 21644 23660 21700 23662
rect 22652 26402 22708 26404
rect 22652 26350 22654 26402
rect 22654 26350 22706 26402
rect 22706 26350 22708 26402
rect 22652 26348 22708 26350
rect 22540 25228 22596 25284
rect 22428 24892 22484 24948
rect 22204 24668 22260 24724
rect 21980 23212 22036 23268
rect 21756 22482 21812 22484
rect 21756 22430 21758 22482
rect 21758 22430 21810 22482
rect 21810 22430 21812 22482
rect 21756 22428 21812 22430
rect 19404 21868 19460 21924
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 21868 22316 21924 22372
rect 23324 25900 23380 25956
rect 23100 25228 23156 25284
rect 23212 23548 23268 23604
rect 23100 22876 23156 22932
rect 22540 22092 22596 22148
rect 19180 21420 19236 21476
rect 18508 17388 18564 17444
rect 18508 17052 18564 17108
rect 18060 16882 18116 16884
rect 18060 16830 18062 16882
rect 18062 16830 18114 16882
rect 18114 16830 18116 16882
rect 18060 16828 18116 16830
rect 19068 18844 19124 18900
rect 18732 16994 18788 16996
rect 18732 16942 18734 16994
rect 18734 16942 18786 16994
rect 18786 16942 18788 16994
rect 18732 16940 18788 16942
rect 18844 18172 18900 18228
rect 17724 16716 17780 16772
rect 18396 16716 18452 16772
rect 18284 16658 18340 16660
rect 18284 16606 18286 16658
rect 18286 16606 18338 16658
rect 18338 16606 18340 16658
rect 18284 16604 18340 16606
rect 17948 15372 18004 15428
rect 18732 16604 18788 16660
rect 17724 15260 17780 15316
rect 17500 14642 17556 14644
rect 17500 14590 17502 14642
rect 17502 14590 17554 14642
rect 17554 14590 17556 14642
rect 17500 14588 17556 14590
rect 20524 21474 20580 21476
rect 20524 21422 20526 21474
rect 20526 21422 20578 21474
rect 20578 21422 20580 21474
rect 20524 21420 20580 21422
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19292 20130 19348 20132
rect 19292 20078 19294 20130
rect 19294 20078 19346 20130
rect 19346 20078 19348 20130
rect 19292 20076 19348 20078
rect 19404 19010 19460 19012
rect 19404 18958 19406 19010
rect 19406 18958 19458 19010
rect 19458 18958 19460 19010
rect 19404 18956 19460 18958
rect 19628 20130 19684 20132
rect 19628 20078 19630 20130
rect 19630 20078 19682 20130
rect 19682 20078 19684 20130
rect 19628 20076 19684 20078
rect 20300 20130 20356 20132
rect 20300 20078 20302 20130
rect 20302 20078 20354 20130
rect 20354 20078 20356 20130
rect 20300 20076 20356 20078
rect 21084 20130 21140 20132
rect 21084 20078 21086 20130
rect 21086 20078 21138 20130
rect 21138 20078 21140 20130
rect 21084 20076 21140 20078
rect 20636 20018 20692 20020
rect 20636 19966 20638 20018
rect 20638 19966 20690 20018
rect 20690 19966 20692 20018
rect 20636 19964 20692 19966
rect 19964 19852 20020 19908
rect 19964 19628 20020 19684
rect 19740 19404 19796 19460
rect 20076 19234 20132 19236
rect 20076 19182 20078 19234
rect 20078 19182 20130 19234
rect 20130 19182 20132 19234
rect 20076 19180 20132 19182
rect 19628 18844 19684 18900
rect 19292 18284 19348 18340
rect 19516 16940 19572 16996
rect 19404 16604 19460 16660
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19964 18450 20020 18452
rect 19964 18398 19966 18450
rect 19966 18398 20018 18450
rect 20018 18398 20020 18450
rect 19964 18396 20020 18398
rect 19740 18284 19796 18340
rect 19740 18060 19796 18116
rect 20972 18620 21028 18676
rect 20748 17666 20804 17668
rect 20748 17614 20750 17666
rect 20750 17614 20802 17666
rect 20802 17614 20804 17666
rect 20748 17612 20804 17614
rect 21196 18172 21252 18228
rect 21308 19516 21364 19572
rect 22204 20972 22260 21028
rect 22988 22146 23044 22148
rect 22988 22094 22990 22146
rect 22990 22094 23042 22146
rect 23042 22094 23044 22146
rect 22988 22092 23044 22094
rect 21532 19516 21588 19572
rect 21532 19122 21588 19124
rect 21532 19070 21534 19122
rect 21534 19070 21586 19122
rect 21586 19070 21588 19122
rect 21532 19068 21588 19070
rect 22428 20076 22484 20132
rect 22092 19068 22148 19124
rect 21420 18396 21476 18452
rect 21644 18450 21700 18452
rect 21644 18398 21646 18450
rect 21646 18398 21698 18450
rect 21698 18398 21700 18450
rect 21644 18396 21700 18398
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19852 17052 19908 17108
rect 20412 16828 20468 16884
rect 21868 16156 21924 16212
rect 20076 15874 20132 15876
rect 20076 15822 20078 15874
rect 20078 15822 20130 15874
rect 20130 15822 20132 15874
rect 20076 15820 20132 15822
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 18956 15426 19012 15428
rect 18956 15374 18958 15426
rect 18958 15374 19010 15426
rect 19010 15374 19012 15426
rect 18956 15372 19012 15374
rect 18732 15314 18788 15316
rect 18732 15262 18734 15314
rect 18734 15262 18786 15314
rect 18786 15262 18788 15314
rect 18732 15260 18788 15262
rect 20300 15372 20356 15428
rect 19852 14588 19908 14644
rect 19180 14140 19236 14196
rect 17948 13916 18004 13972
rect 14924 12908 14980 12964
rect 17724 12962 17780 12964
rect 17724 12910 17726 12962
rect 17726 12910 17778 12962
rect 17778 12910 17780 12962
rect 17724 12908 17780 12910
rect 19740 14252 19796 14308
rect 20748 15820 20804 15876
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19964 12290 20020 12292
rect 19964 12238 19966 12290
rect 19966 12238 20018 12290
rect 20018 12238 20020 12290
rect 19964 12236 20020 12238
rect 20412 12236 20468 12292
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 17500 3612 17556 3668
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 21644 14588 21700 14644
rect 20972 13970 21028 13972
rect 20972 13918 20974 13970
rect 20974 13918 21026 13970
rect 21026 13918 21028 13970
rect 20972 13916 21028 13918
rect 21756 13916 21812 13972
rect 22204 18396 22260 18452
rect 22204 18060 22260 18116
rect 22652 19906 22708 19908
rect 22652 19854 22654 19906
rect 22654 19854 22706 19906
rect 22706 19854 22708 19906
rect 22652 19852 22708 19854
rect 22764 19516 22820 19572
rect 22652 19180 22708 19236
rect 22988 20690 23044 20692
rect 22988 20638 22990 20690
rect 22990 20638 23042 20690
rect 23042 20638 23044 20690
rect 22988 20636 23044 20638
rect 22876 19292 22932 19348
rect 22540 19068 22596 19124
rect 22428 18508 22484 18564
rect 22652 18284 22708 18340
rect 23100 18674 23156 18676
rect 23100 18622 23102 18674
rect 23102 18622 23154 18674
rect 23154 18622 23156 18674
rect 23100 18620 23156 18622
rect 24332 27858 24388 27860
rect 24332 27806 24334 27858
rect 24334 27806 24386 27858
rect 24386 27806 24388 27858
rect 24332 27804 24388 27806
rect 26012 26348 26068 26404
rect 23660 24668 23716 24724
rect 25228 26236 25284 26292
rect 24780 24780 24836 24836
rect 25340 24946 25396 24948
rect 25340 24894 25342 24946
rect 25342 24894 25394 24946
rect 25394 24894 25396 24946
rect 25340 24892 25396 24894
rect 25564 24892 25620 24948
rect 26236 24892 26292 24948
rect 25676 24722 25732 24724
rect 25676 24670 25678 24722
rect 25678 24670 25730 24722
rect 25730 24670 25732 24722
rect 25676 24668 25732 24670
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 27020 24892 27076 24948
rect 26460 24834 26516 24836
rect 26460 24782 26462 24834
rect 26462 24782 26514 24834
rect 26514 24782 26516 24834
rect 26460 24780 26516 24782
rect 37660 24722 37716 24724
rect 37660 24670 37662 24722
rect 37662 24670 37714 24722
rect 37714 24670 37716 24722
rect 37660 24668 37716 24670
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 40012 24220 40068 24276
rect 24108 23660 24164 23716
rect 23884 22876 23940 22932
rect 23660 22316 23716 22372
rect 23324 20972 23380 21028
rect 23324 18562 23380 18564
rect 23324 18510 23326 18562
rect 23326 18510 23378 18562
rect 23378 18510 23380 18562
rect 23324 18508 23380 18510
rect 23660 18450 23716 18452
rect 23660 18398 23662 18450
rect 23662 18398 23714 18450
rect 23714 18398 23716 18450
rect 23660 18396 23716 18398
rect 23436 18338 23492 18340
rect 23436 18286 23438 18338
rect 23438 18286 23490 18338
rect 23490 18286 23492 18338
rect 23436 18284 23492 18286
rect 22652 17666 22708 17668
rect 22652 17614 22654 17666
rect 22654 17614 22706 17666
rect 22706 17614 22708 17666
rect 22652 17612 22708 17614
rect 24332 23378 24388 23380
rect 24332 23326 24334 23378
rect 24334 23326 24386 23378
rect 24386 23326 24388 23378
rect 24332 23324 24388 23326
rect 40012 23548 40068 23604
rect 37660 23436 37716 23492
rect 25228 23324 25284 23380
rect 27356 23212 27412 23268
rect 26572 22258 26628 22260
rect 26572 22206 26574 22258
rect 26574 22206 26626 22258
rect 26626 22206 26628 22258
rect 26572 22204 26628 22206
rect 28700 23212 28756 23268
rect 37660 23154 37716 23156
rect 37660 23102 37662 23154
rect 37662 23102 37714 23154
rect 37714 23102 37716 23154
rect 37660 23100 37716 23102
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 27244 21756 27300 21812
rect 25340 20972 25396 21028
rect 26348 20690 26404 20692
rect 26348 20638 26350 20690
rect 26350 20638 26402 20690
rect 26402 20638 26404 20690
rect 26348 20636 26404 20638
rect 28588 21756 28644 21812
rect 37660 21756 37716 21812
rect 40012 21532 40068 21588
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 25676 20578 25732 20580
rect 25676 20526 25678 20578
rect 25678 20526 25730 20578
rect 25730 20526 25732 20578
rect 25676 20524 25732 20526
rect 26908 20412 26964 20468
rect 24668 19852 24724 19908
rect 26236 19122 26292 19124
rect 26236 19070 26238 19122
rect 26238 19070 26290 19122
rect 26290 19070 26292 19122
rect 26236 19068 26292 19070
rect 26460 19010 26516 19012
rect 26460 18958 26462 19010
rect 26462 18958 26514 19010
rect 26514 18958 26516 19010
rect 26460 18956 26516 18958
rect 26236 18620 26292 18676
rect 22316 16492 22372 16548
rect 21980 15036 22036 15092
rect 21980 14530 22036 14532
rect 21980 14478 21982 14530
rect 21982 14478 22034 14530
rect 22034 14478 22036 14530
rect 21980 14476 22036 14478
rect 22204 14476 22260 14532
rect 22540 14642 22596 14644
rect 22540 14590 22542 14642
rect 22542 14590 22594 14642
rect 22594 14590 22596 14642
rect 22540 14588 22596 14590
rect 23324 16210 23380 16212
rect 23324 16158 23326 16210
rect 23326 16158 23378 16210
rect 23378 16158 23380 16210
rect 23324 16156 23380 16158
rect 23772 16156 23828 16212
rect 24108 15538 24164 15540
rect 24108 15486 24110 15538
rect 24110 15486 24162 15538
rect 24162 15486 24164 15538
rect 24108 15484 24164 15486
rect 27468 19628 27524 19684
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 28364 19234 28420 19236
rect 28364 19182 28366 19234
rect 28366 19182 28418 19234
rect 28418 19182 28420 19234
rect 28364 19180 28420 19182
rect 28924 19180 28980 19236
rect 27244 19122 27300 19124
rect 27244 19070 27246 19122
rect 27246 19070 27298 19122
rect 27298 19070 27300 19122
rect 27244 19068 27300 19070
rect 27132 18956 27188 19012
rect 26796 18508 26852 18564
rect 27804 19010 27860 19012
rect 27804 18958 27806 19010
rect 27806 18958 27858 19010
rect 27858 18958 27860 19010
rect 27804 18956 27860 18958
rect 27580 18508 27636 18564
rect 28588 18396 28644 18452
rect 37660 19234 37716 19236
rect 37660 19182 37662 19234
rect 37662 19182 37714 19234
rect 37714 19182 37716 19234
rect 37660 19180 37716 19182
rect 40012 18844 40068 18900
rect 37660 18450 37716 18452
rect 37660 18398 37662 18450
rect 37662 18398 37714 18450
rect 37714 18398 37716 18450
rect 37660 18396 37716 18398
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 26684 17052 26740 17108
rect 27916 17106 27972 17108
rect 27916 17054 27918 17106
rect 27918 17054 27970 17106
rect 27970 17054 27972 17106
rect 27916 17052 27972 17054
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 25340 16156 25396 16212
rect 25564 16156 25620 16212
rect 26572 16210 26628 16212
rect 26572 16158 26574 16210
rect 26574 16158 26626 16210
rect 26626 16158 26628 16210
rect 26572 16156 26628 16158
rect 25564 15484 25620 15540
rect 23996 15426 24052 15428
rect 23996 15374 23998 15426
rect 23998 15374 24050 15426
rect 24050 15374 24052 15426
rect 23996 15372 24052 15374
rect 23212 15036 23268 15092
rect 23996 15036 24052 15092
rect 22988 14588 23044 14644
rect 23660 14642 23716 14644
rect 23660 14590 23662 14642
rect 23662 14590 23714 14642
rect 23714 14590 23716 14642
rect 23660 14588 23716 14590
rect 22876 14530 22932 14532
rect 22876 14478 22878 14530
rect 22878 14478 22930 14530
rect 22930 14478 22932 14530
rect 22876 14476 22932 14478
rect 23436 14530 23492 14532
rect 23436 14478 23438 14530
rect 23438 14478 23490 14530
rect 23490 14478 23492 14530
rect 23436 14476 23492 14478
rect 23324 13804 23380 13860
rect 25228 13858 25284 13860
rect 25228 13806 25230 13858
rect 25230 13806 25282 13858
rect 25282 13806 25284 13858
rect 25228 13804 25284 13806
rect 24668 13634 24724 13636
rect 24668 13582 24670 13634
rect 24670 13582 24722 13634
rect 24722 13582 24724 13634
rect 24668 13580 24724 13582
rect 25340 13634 25396 13636
rect 25340 13582 25342 13634
rect 25342 13582 25394 13634
rect 25394 13582 25396 13634
rect 25340 13580 25396 13582
rect 21868 12962 21924 12964
rect 21868 12910 21870 12962
rect 21870 12910 21922 12962
rect 21922 12910 21924 12962
rect 21868 12908 21924 12910
rect 25228 12962 25284 12964
rect 25228 12910 25230 12962
rect 25230 12910 25282 12962
rect 25282 12910 25284 12962
rect 25228 12908 25284 12910
rect 20188 4060 20244 4116
rect 18620 3666 18676 3668
rect 18620 3614 18622 3666
rect 18622 3614 18674 3666
rect 18674 3614 18676 3666
rect 18620 3612 18676 3614
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 20860 3612 20916 3668
rect 21420 4114 21476 4116
rect 21420 4062 21422 4114
rect 21422 4062 21474 4114
rect 21474 4062 21476 4114
rect 21420 4060 21476 4062
rect 24220 4060 24276 4116
rect 22092 3666 22148 3668
rect 22092 3614 22094 3666
rect 22094 3614 22146 3666
rect 22146 3614 22148 3666
rect 22092 3612 22148 3614
rect 23548 3612 23604 3668
rect 24892 5180 24948 5236
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 25564 13580 25620 13636
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 25676 12908 25732 12964
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 26124 5234 26180 5236
rect 26124 5182 26126 5234
rect 26126 5182 26178 5234
rect 26178 5182 26180 5234
rect 26124 5180 26180 5182
rect 26236 4114 26292 4116
rect 26236 4062 26238 4114
rect 26238 4062 26290 4114
rect 26290 4062 26292 4114
rect 26236 4060 26292 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 17490 38220 17500 38276
rect 17556 38220 18620 38276
rect 18676 38220 18686 38276
rect 23538 38220 23548 38276
rect 23604 38220 24780 38276
rect 24836 38220 24846 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 18834 37436 18844 37492
rect 18900 37436 19852 37492
rect 19908 37436 19918 37492
rect 21522 37436 21532 37492
rect 21588 37436 22764 37492
rect 22820 37436 22830 37492
rect 24210 37436 24220 37492
rect 24276 37436 26236 37492
rect 26292 37436 26302 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 20178 36652 20188 36708
rect 20244 36652 22316 36708
rect 22372 36652 22382 36708
rect 25554 36652 25564 36708
rect 25620 36652 26796 36708
rect 26852 36652 26862 36708
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 0 35700 800 35728
rect 0 35644 1708 35700
rect 1764 35644 1774 35700
rect 0 35616 800 35644
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 20290 28364 20300 28420
rect 20356 28364 21308 28420
rect 21364 28364 21374 28420
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 24434 28028 24444 28084
rect 24500 28028 25788 28084
rect 25844 28028 25854 28084
rect 16706 27916 16716 27972
rect 16772 27916 17500 27972
rect 17556 27916 17566 27972
rect 21746 27916 21756 27972
rect 21812 27916 22428 27972
rect 22484 27916 22764 27972
rect 22820 27916 22830 27972
rect 16818 27804 16828 27860
rect 16884 27804 18620 27860
rect 18676 27804 21980 27860
rect 22036 27804 24332 27860
rect 24388 27804 24398 27860
rect 17490 27692 17500 27748
rect 17556 27692 17836 27748
rect 17892 27692 17902 27748
rect 0 27636 800 27664
rect 0 27580 4172 27636
rect 4228 27580 4238 27636
rect 17042 27580 17052 27636
rect 17108 27580 17724 27636
rect 17780 27580 17790 27636
rect 0 27552 800 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 14914 27132 14924 27188
rect 14980 27132 16268 27188
rect 16324 27132 16334 27188
rect 18274 26908 18284 26964
rect 18340 26908 19516 26964
rect 19572 26908 20636 26964
rect 20692 26908 20702 26964
rect 21522 26908 21532 26964
rect 21588 26908 22988 26964
rect 23044 26908 23054 26964
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 22642 26348 22652 26404
rect 22708 26348 26012 26404
rect 26068 26348 26078 26404
rect 4274 26236 4284 26292
rect 4340 26236 8428 26292
rect 22082 26236 22092 26292
rect 22148 26236 25228 26292
rect 25284 26236 25294 26292
rect 8372 26180 8428 26236
rect 8372 26124 11116 26180
rect 11172 26124 11182 26180
rect 13234 26124 13244 26180
rect 13300 26124 15932 26180
rect 15988 26124 15998 26180
rect 23324 25956 23380 26236
rect 23314 25900 23324 25956
rect 23380 25900 23390 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 0 25620 800 25648
rect 0 25564 1932 25620
rect 1988 25564 1998 25620
rect 11106 25564 11116 25620
rect 11172 25564 14364 25620
rect 14420 25564 14430 25620
rect 0 25536 800 25564
rect 4274 25452 4284 25508
rect 4340 25452 12796 25508
rect 12852 25452 12862 25508
rect 14914 25228 14924 25284
rect 14980 25228 15484 25284
rect 15540 25228 17500 25284
rect 17556 25228 18172 25284
rect 18228 25228 18238 25284
rect 20626 25228 20636 25284
rect 20692 25228 21532 25284
rect 21588 25228 22540 25284
rect 22596 25228 23100 25284
rect 23156 25228 23166 25284
rect 16146 25116 16156 25172
rect 16212 25116 17276 25172
rect 17332 25116 17342 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 21298 25004 21308 25060
rect 21364 25004 21756 25060
rect 21812 25004 21822 25060
rect 0 24948 800 24976
rect 0 24892 2044 24948
rect 2100 24892 2110 24948
rect 22418 24892 22428 24948
rect 22484 24892 25340 24948
rect 25396 24892 25406 24948
rect 25554 24892 25564 24948
rect 25620 24892 26236 24948
rect 26292 24892 27020 24948
rect 27076 24892 27086 24948
rect 0 24864 800 24892
rect 25564 24836 25620 24892
rect 24770 24780 24780 24836
rect 24836 24780 25620 24836
rect 26450 24780 26460 24836
rect 26516 24780 31948 24836
rect 31892 24724 31948 24780
rect 12786 24668 12796 24724
rect 12852 24668 16268 24724
rect 16324 24668 16334 24724
rect 21532 24668 22204 24724
rect 22260 24668 22270 24724
rect 23650 24668 23660 24724
rect 23716 24668 25676 24724
rect 25732 24668 25742 24724
rect 31892 24668 37660 24724
rect 37716 24668 37726 24724
rect 21532 24612 21588 24668
rect 21522 24556 21532 24612
rect 21588 24556 21598 24612
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 41200 24276 42000 24304
rect 40002 24220 40012 24276
rect 40068 24220 42000 24276
rect 41200 24192 42000 24220
rect 15362 24108 15372 24164
rect 15428 24108 17612 24164
rect 17668 24108 17678 24164
rect 16706 23884 16716 23940
rect 16772 23884 21308 23940
rect 21364 23884 21374 23940
rect 15362 23772 15372 23828
rect 15428 23772 21532 23828
rect 21588 23772 21598 23828
rect 18274 23660 18284 23716
rect 18340 23660 21420 23716
rect 21476 23660 21486 23716
rect 21634 23660 21644 23716
rect 21700 23660 24108 23716
rect 24164 23660 24174 23716
rect 41200 23604 42000 23632
rect 21298 23548 21308 23604
rect 21364 23548 23212 23604
rect 23268 23548 23278 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 41200 23520 42000 23548
rect 31892 23436 37660 23492
rect 37716 23436 37726 23492
rect 15092 23324 15484 23380
rect 15540 23324 16156 23380
rect 16212 23324 21084 23380
rect 21140 23324 24332 23380
rect 24388 23324 25228 23380
rect 25284 23324 25294 23380
rect 15092 23044 15148 23324
rect 31892 23268 31948 23436
rect 17266 23212 17276 23268
rect 17332 23212 18732 23268
rect 18788 23212 18798 23268
rect 19730 23212 19740 23268
rect 19796 23212 21980 23268
rect 22036 23212 22046 23268
rect 27346 23212 27356 23268
rect 27412 23212 28700 23268
rect 28756 23212 31948 23268
rect 31892 23100 37660 23156
rect 37716 23100 37726 23156
rect 11442 22988 11452 23044
rect 11508 22988 13132 23044
rect 13188 22988 14700 23044
rect 14756 22988 15148 23044
rect 17266 22988 17276 23044
rect 17332 22988 17500 23044
rect 17556 22988 19404 23044
rect 19460 22988 19470 23044
rect 31892 22932 31948 23100
rect 41200 22932 42000 22960
rect 23090 22876 23100 22932
rect 23156 22876 23884 22932
rect 23940 22876 31948 22932
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 41200 22848 42000 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 20150 22540 20188 22596
rect 20244 22540 20254 22596
rect 12114 22428 12124 22484
rect 12180 22428 14700 22484
rect 14756 22428 14766 22484
rect 17154 22428 17164 22484
rect 17220 22428 21756 22484
rect 21812 22428 21822 22484
rect 14130 22316 14140 22372
rect 14196 22316 14812 22372
rect 14868 22316 14878 22372
rect 19730 22316 19740 22372
rect 19796 22316 21868 22372
rect 21924 22316 23660 22372
rect 23716 22316 23726 22372
rect 19180 22204 20300 22260
rect 20356 22204 26572 22260
rect 26628 22204 26638 22260
rect 19180 22148 19236 22204
rect 15250 22092 15260 22148
rect 15316 22092 15932 22148
rect 15988 22092 19236 22148
rect 19394 22092 19404 22148
rect 19460 22092 20188 22148
rect 20244 22092 20254 22148
rect 22530 22092 22540 22148
rect 22596 22092 22988 22148
rect 23044 22092 23054 22148
rect 15810 21980 15820 22036
rect 15876 21980 17388 22036
rect 17444 21980 17454 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 16930 21868 16940 21924
rect 16996 21868 17164 21924
rect 17220 21868 17230 21924
rect 18834 21868 18844 21924
rect 18900 21868 19404 21924
rect 19460 21868 19470 21924
rect 15698 21756 15708 21812
rect 15764 21756 17388 21812
rect 17444 21756 17454 21812
rect 27234 21756 27244 21812
rect 27300 21756 28588 21812
rect 28644 21756 37660 21812
rect 37716 21756 37726 21812
rect 14242 21644 14252 21700
rect 14308 21644 15148 21700
rect 15204 21644 15214 21700
rect 41200 21588 42000 21616
rect 4274 21532 4284 21588
rect 4340 21532 9996 21588
rect 10052 21532 10062 21588
rect 14578 21532 14588 21588
rect 14644 21532 17724 21588
rect 17780 21532 18956 21588
rect 19012 21532 19022 21588
rect 40002 21532 40012 21588
rect 40068 21532 42000 21588
rect 41200 21504 42000 21532
rect 4162 21420 4172 21476
rect 4228 21420 18172 21476
rect 18228 21420 18238 21476
rect 19170 21420 19180 21476
rect 19236 21420 20524 21476
rect 20580 21420 20590 21476
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 22194 20972 22204 21028
rect 22260 20972 23324 21028
rect 23380 20972 25340 21028
rect 25396 20972 25406 21028
rect 0 20916 800 20944
rect 0 20860 1932 20916
rect 1988 20860 1998 20916
rect 9986 20860 9996 20916
rect 10052 20860 13244 20916
rect 13300 20860 13310 20916
rect 15138 20860 15148 20916
rect 15204 20860 16156 20916
rect 16212 20860 18284 20916
rect 18340 20860 18350 20916
rect 0 20832 800 20860
rect 15922 20748 15932 20804
rect 15988 20748 17164 20804
rect 17220 20748 17230 20804
rect 22978 20636 22988 20692
rect 23044 20636 26348 20692
rect 26404 20636 26414 20692
rect 12114 20524 12124 20580
rect 12180 20524 13468 20580
rect 13524 20524 13534 20580
rect 25666 20524 25676 20580
rect 25732 20524 26908 20580
rect 26852 20412 26908 20524
rect 26964 20412 26974 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 14242 20076 14252 20132
rect 14308 20076 15148 20132
rect 15250 20076 15260 20132
rect 15316 20076 16156 20132
rect 16212 20076 17500 20132
rect 17556 20076 17566 20132
rect 18386 20076 18396 20132
rect 18452 20076 19292 20132
rect 19348 20076 19358 20132
rect 19618 20076 19628 20132
rect 19684 20076 20300 20132
rect 20356 20076 21084 20132
rect 21140 20076 22428 20132
rect 22484 20076 22494 20132
rect 15092 20020 15148 20076
rect 4274 19964 4284 20020
rect 4340 19964 9996 20020
rect 10052 19964 10062 20020
rect 15092 19964 17836 20020
rect 17892 19964 20636 20020
rect 20692 19964 20702 20020
rect 13570 19852 13580 19908
rect 13636 19852 18732 19908
rect 18788 19852 19964 19908
rect 20020 19852 20188 19908
rect 20244 19852 20254 19908
rect 22642 19852 22652 19908
rect 22708 19852 24668 19908
rect 24724 19852 24734 19908
rect 1922 19740 1932 19796
rect 1988 19740 1998 19796
rect 12114 19740 12124 19796
rect 12180 19740 13916 19796
rect 13972 19740 13982 19796
rect 0 19572 800 19600
rect 1932 19572 1988 19740
rect 19954 19628 19964 19684
rect 20020 19628 27468 19684
rect 27524 19628 27534 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 0 19516 1988 19572
rect 13682 19516 13692 19572
rect 13748 19516 17612 19572
rect 17668 19516 21308 19572
rect 21364 19516 21532 19572
rect 21588 19516 22764 19572
rect 22820 19516 22830 19572
rect 0 19488 800 19516
rect 16594 19404 16604 19460
rect 16660 19404 16698 19460
rect 18498 19404 18508 19460
rect 18564 19404 19740 19460
rect 19796 19404 19806 19460
rect 9986 19292 9996 19348
rect 10052 19292 16380 19348
rect 16436 19292 16446 19348
rect 16818 19292 16828 19348
rect 16884 19292 22876 19348
rect 22932 19292 22942 19348
rect 12898 19180 12908 19236
rect 12964 19180 13580 19236
rect 13636 19180 13646 19236
rect 14242 19180 14252 19236
rect 14308 19180 16492 19236
rect 16548 19180 16558 19236
rect 18946 19180 18956 19236
rect 19012 19180 20076 19236
rect 20132 19180 22652 19236
rect 22708 19180 22718 19236
rect 28354 19180 28364 19236
rect 28420 19180 28924 19236
rect 28980 19180 37660 19236
rect 37716 19180 37726 19236
rect 15922 19068 15932 19124
rect 15988 19068 17836 19124
rect 17892 19068 17902 19124
rect 21522 19068 21532 19124
rect 21588 19068 22092 19124
rect 22148 19068 22540 19124
rect 22596 19068 22606 19124
rect 26226 19068 26236 19124
rect 26292 19068 27244 19124
rect 27300 19068 27310 19124
rect 16482 18956 16492 19012
rect 16548 18956 18228 19012
rect 19394 18956 19404 19012
rect 19460 18956 26460 19012
rect 26516 18956 26526 19012
rect 27122 18956 27132 19012
rect 27188 18956 27804 19012
rect 27860 18956 27870 19012
rect 18172 18900 18228 18956
rect 41200 18900 42000 18928
rect 15810 18844 15820 18900
rect 15876 18844 16716 18900
rect 16772 18844 16782 18900
rect 18162 18844 18172 18900
rect 18228 18844 19068 18900
rect 19124 18844 19628 18900
rect 19684 18844 19694 18900
rect 40002 18844 40012 18900
rect 40068 18844 42000 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 41200 18816 42000 18844
rect 16594 18620 16604 18676
rect 16660 18620 17388 18676
rect 17444 18620 20972 18676
rect 21028 18620 21038 18676
rect 23090 18620 23100 18676
rect 23156 18620 26236 18676
rect 26292 18620 26302 18676
rect 22418 18508 22428 18564
rect 22484 18508 23324 18564
rect 23380 18508 23390 18564
rect 26786 18508 26796 18564
rect 26852 18508 27580 18564
rect 27636 18508 27646 18564
rect 16482 18396 16492 18452
rect 16548 18396 16604 18452
rect 16660 18396 17836 18452
rect 17892 18396 17902 18452
rect 19954 18396 19964 18452
rect 20020 18396 21420 18452
rect 21476 18396 21486 18452
rect 21634 18396 21644 18452
rect 21700 18396 21710 18452
rect 22194 18396 22204 18452
rect 22260 18396 23660 18452
rect 23716 18396 23726 18452
rect 28578 18396 28588 18452
rect 28644 18396 37660 18452
rect 37716 18396 37726 18452
rect 21644 18340 21700 18396
rect 16146 18284 16156 18340
rect 16212 18284 17612 18340
rect 17668 18284 17678 18340
rect 17938 18284 17948 18340
rect 18004 18284 19292 18340
rect 19348 18284 19740 18340
rect 19796 18284 19806 18340
rect 21532 18284 21700 18340
rect 22642 18284 22652 18340
rect 22708 18284 23436 18340
rect 23492 18284 23502 18340
rect 21532 18228 21588 18284
rect 41200 18228 42000 18256
rect 14242 18172 14252 18228
rect 14308 18172 15036 18228
rect 15092 18172 15102 18228
rect 18834 18172 18844 18228
rect 18900 18172 21196 18228
rect 21252 18172 21588 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 41200 18144 42000 18172
rect 15586 18060 15596 18116
rect 15652 18060 19740 18116
rect 19796 18060 22204 18116
rect 22260 18060 22270 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 14466 17836 14476 17892
rect 14532 17836 16604 17892
rect 16660 17836 17164 17892
rect 17220 17836 18060 17892
rect 18116 17836 18126 17892
rect 15586 17724 15596 17780
rect 15652 17724 16268 17780
rect 16324 17724 16334 17780
rect 20738 17612 20748 17668
rect 20804 17612 22652 17668
rect 22708 17612 22718 17668
rect 11218 17388 11228 17444
rect 11284 17388 14476 17444
rect 14532 17388 14542 17444
rect 16370 17388 16380 17444
rect 16436 17388 18508 17444
rect 18564 17388 18574 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 14466 17052 14476 17108
rect 14532 17052 15372 17108
rect 15428 17052 15438 17108
rect 18498 17052 18508 17108
rect 18564 17052 19852 17108
rect 19908 17052 19918 17108
rect 26674 17052 26684 17108
rect 26740 17052 27916 17108
rect 27972 17052 27982 17108
rect 15586 16940 15596 16996
rect 15652 16940 16380 16996
rect 16436 16940 17836 16996
rect 17892 16940 17902 16996
rect 18722 16940 18732 16996
rect 18788 16940 19516 16996
rect 19572 16940 19582 16996
rect 13458 16828 13468 16884
rect 13524 16828 14252 16884
rect 14308 16828 16044 16884
rect 16100 16828 16110 16884
rect 17378 16828 17388 16884
rect 17444 16828 18060 16884
rect 18116 16828 20412 16884
rect 20468 16828 20478 16884
rect 16258 16716 16268 16772
rect 16324 16716 17724 16772
rect 17780 16716 18396 16772
rect 18452 16716 18462 16772
rect 15698 16604 15708 16660
rect 15764 16604 16940 16660
rect 16996 16604 17006 16660
rect 18274 16604 18284 16660
rect 18340 16604 18732 16660
rect 18788 16604 19404 16660
rect 19460 16604 19470 16660
rect 16940 16548 16996 16604
rect 16940 16492 22316 16548
rect 22372 16492 22382 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 21858 16156 21868 16212
rect 21924 16156 23324 16212
rect 23380 16156 23772 16212
rect 23828 16156 25340 16212
rect 25396 16156 25406 16212
rect 25554 16156 25564 16212
rect 25620 16156 26572 16212
rect 26628 16156 26638 16212
rect 12562 16044 12572 16100
rect 12628 16044 17164 16100
rect 17220 16044 17230 16100
rect 20066 15820 20076 15876
rect 20132 15820 20748 15876
rect 20804 15820 20814 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 14466 15484 14476 15540
rect 14532 15484 15036 15540
rect 15092 15484 15102 15540
rect 24098 15484 24108 15540
rect 24164 15484 25564 15540
rect 25620 15484 25630 15540
rect 17938 15372 17948 15428
rect 18004 15372 18956 15428
rect 19012 15372 20300 15428
rect 20356 15372 23996 15428
rect 24052 15372 24062 15428
rect 17714 15260 17724 15316
rect 17780 15260 18732 15316
rect 18788 15260 18798 15316
rect 10546 15148 10556 15204
rect 10612 15148 11676 15204
rect 11732 15148 13804 15204
rect 13860 15148 14924 15204
rect 14980 15148 14990 15204
rect 21970 15036 21980 15092
rect 22036 15036 23212 15092
rect 23268 15036 23996 15092
rect 24052 15036 24062 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 17490 14588 17500 14644
rect 17556 14588 17566 14644
rect 19842 14588 19852 14644
rect 19908 14588 21644 14644
rect 21700 14588 22540 14644
rect 22596 14588 22606 14644
rect 22978 14588 22988 14644
rect 23044 14588 23660 14644
rect 23716 14588 23726 14644
rect 17500 14532 17556 14588
rect 17500 14476 21980 14532
rect 22036 14476 22046 14532
rect 22194 14476 22204 14532
rect 22260 14476 22876 14532
rect 22932 14476 23436 14532
rect 23492 14476 23502 14532
rect 19180 14252 19740 14308
rect 19796 14252 19806 14308
rect 19180 14196 19236 14252
rect 19170 14140 19180 14196
rect 19236 14140 19246 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 17938 13916 17948 13972
rect 18004 13916 20972 13972
rect 21028 13916 21756 13972
rect 21812 13916 21822 13972
rect 23314 13804 23324 13860
rect 23380 13804 25228 13860
rect 25284 13804 25294 13860
rect 24658 13580 24668 13636
rect 24724 13580 25340 13636
rect 25396 13580 25564 13636
rect 25620 13580 25630 13636
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 14466 12908 14476 12964
rect 14532 12908 14924 12964
rect 14980 12908 17724 12964
rect 17780 12908 17790 12964
rect 21858 12908 21868 12964
rect 21924 12908 25228 12964
rect 25284 12908 25676 12964
rect 25732 12908 25742 12964
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 19954 12236 19964 12292
rect 20020 12236 20412 12292
rect 20468 12236 20478 12292
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 24882 5180 24892 5236
rect 24948 5180 26124 5236
rect 26180 5180 26190 5236
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 20178 4060 20188 4116
rect 20244 4060 21420 4116
rect 21476 4060 21486 4116
rect 24210 4060 24220 4116
rect 24276 4060 26236 4116
rect 26292 4060 26302 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 17490 3612 17500 3668
rect 17556 3612 18620 3668
rect 18676 3612 18686 3668
rect 20850 3612 20860 3668
rect 20916 3612 22092 3668
rect 22148 3612 22158 3668
rect 23538 3612 23548 3668
rect 23604 3612 25564 3668
rect 25620 3612 25630 3668
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 20188 22540 20244 22596
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 20188 19852 20244 19908
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 16604 19404 16660 19460
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 16604 18396 16660 18452
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 16604 19460 16660 19470
rect 16604 18452 16660 19404
rect 16604 18386 16660 18396
rect 19808 18844 20128 20356
rect 20188 22596 20244 22606
rect 20188 19908 20244 22540
rect 20188 19842 20244 19852
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14000 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _107_
timestamp 1698175906
transform 1 0 15232 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_
timestamp 1698175906
transform -1 0 15344 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14896 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1698175906
transform 1 0 15680 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22400 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1698175906
transform -1 0 20048 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18144 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1698175906
transform 1 0 19152 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform -1 0 20496 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19936 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform -1 0 18032 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _118_
timestamp 1698175906
transform 1 0 19152 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _119_
timestamp 1698175906
transform -1 0 23296 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15344 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _122_
timestamp 1698175906
transform -1 0 21728 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _123_
timestamp 1698175906
transform -1 0 22176 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _124_
timestamp 1698175906
transform 1 0 15904 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform -1 0 22176 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698175906
transform 1 0 18480 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14224 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16128 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform 1 0 15344 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform 1 0 17696 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19488 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _134_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20272 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _136_
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _137_
timestamp 1698175906
transform 1 0 23184 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _138_
timestamp 1698175906
transform -1 0 22848 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _139_
timestamp 1698175906
transform 1 0 22512 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _140_
timestamp 1698175906
transform -1 0 22512 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _141_
timestamp 1698175906
transform 1 0 25200 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform -1 0 27552 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _143_
timestamp 1698175906
transform -1 0 26656 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _144_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14672 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _145_
timestamp 1698175906
transform -1 0 13104 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _146_
timestamp 1698175906
transform 1 0 13328 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _147_
timestamp 1698175906
transform 1 0 15008 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_
timestamp 1698175906
transform 1 0 15456 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _149_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14448 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _150_
timestamp 1698175906
transform 1 0 22400 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _151_
timestamp 1698175906
transform -1 0 17696 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _152_
timestamp 1698175906
transform -1 0 17024 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _153_
timestamp 1698175906
transform -1 0 14448 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _154_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14784 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _155_
timestamp 1698175906
transform 1 0 14224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _156_
timestamp 1698175906
transform -1 0 17024 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _157_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14672 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _158_
timestamp 1698175906
transform 1 0 16016 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _159_
timestamp 1698175906
transform 1 0 15680 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform -1 0 27664 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _161_
timestamp 1698175906
transform -1 0 26880 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _162_
timestamp 1698175906
transform -1 0 16576 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _163_
timestamp 1698175906
transform 1 0 18144 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _164_
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _165_
timestamp 1698175906
transform -1 0 22288 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _166_
timestamp 1698175906
transform 1 0 24192 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _167_
timestamp 1698175906
transform -1 0 24192 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _168_
timestamp 1698175906
transform -1 0 17696 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _169_
timestamp 1698175906
transform 1 0 15904 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _170_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14784 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _171_
timestamp 1698175906
transform -1 0 17024 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _172_
timestamp 1698175906
transform -1 0 16912 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _173_
timestamp 1698175906
transform -1 0 20160 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _174_
timestamp 1698175906
transform -1 0 20944 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _175_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17696 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _176_
timestamp 1698175906
transform -1 0 20048 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _177_
timestamp 1698175906
transform 1 0 15904 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _178_
timestamp 1698175906
transform 1 0 17024 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _179_
timestamp 1698175906
transform -1 0 18144 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _180_
timestamp 1698175906
transform -1 0 17696 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _181_
timestamp 1698175906
transform -1 0 16464 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _182_
timestamp 1698175906
transform 1 0 23856 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _183_
timestamp 1698175906
transform 1 0 22848 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _184_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23520 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _185_
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _186_
timestamp 1698175906
transform -1 0 21616 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _187_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18704 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _188_
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _189_
timestamp 1698175906
transform 1 0 21728 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _190_
timestamp 1698175906
transform 1 0 22288 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _191_
timestamp 1698175906
transform 1 0 23296 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _192_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14784 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _193_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21952 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _194_
timestamp 1698175906
transform 1 0 23408 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _195_
timestamp 1698175906
transform 1 0 22288 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _196_
timestamp 1698175906
transform -1 0 13776 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _197_
timestamp 1698175906
transform -1 0 14448 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _198_
timestamp 1698175906
transform -1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _199_
timestamp 1698175906
transform -1 0 20496 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _200_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23184 0 -1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _201_
timestamp 1698175906
transform 1 0 27104 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _202_
timestamp 1698175906
transform -1 0 28224 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _203_
timestamp 1698175906
transform 1 0 18704 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _204_
timestamp 1698175906
transform 1 0 26096 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _205_
timestamp 1698175906
transform -1 0 25536 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _206_
timestamp 1698175906
transform -1 0 23408 0 1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _207_
timestamp 1698175906
transform -1 0 18816 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _208_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16912 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _209_
timestamp 1698175906
transform 1 0 17472 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _210_
timestamp 1698175906
transform 1 0 19600 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _211_
timestamp 1698175906
transform 1 0 17808 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20832 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 17696 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 25536 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 10304 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 11424 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 11200 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform -1 0 25648 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform -1 0 13104 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform -1 0 14224 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 25648 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 22736 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform -1 0 15904 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 14784 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 17472 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 14224 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform 1 0 23520 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 19376 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 21728 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 22960 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 21728 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform -1 0 13104 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform 1 0 25872 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 25536 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform 1 0 21616 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform 1 0 16128 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 17360 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _240_
timestamp 1698175906
transform 1 0 25984 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _241_
timestamp 1698175906
transform 1 0 22624 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 20944 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 13776 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 14896 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 14672 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 25872 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 13552 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 14448 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 25424 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 22512 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 16128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 18256 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 21392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform -1 0 17696 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 23296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 22624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 25200 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 21504 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 25200 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 13104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 25648 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 25312 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 25760 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform 1 0 19600 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 20608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 18144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18368 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform 1 0 18928 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 18704 0 -1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698175906
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698175906
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_158 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19040 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_166
timestamp 1698175906
transform 1 0 19936 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_168
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_195
timestamp 1698175906
transform 1 0 23184 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_203
timestamp 1698175906
transform 1 0 24080 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 28000 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 31584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_209
timestamp 1698175906
transform 1 0 24752 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_237
timestamp 1698175906
transform 1 0 27888 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_146
timestamp 1698175906
transform 1 0 17696 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_162
timestamp 1698175906
transform 1 0 19488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_168
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_200
timestamp 1698175906
transform 1 0 23744 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698175906
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698175906
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_181
timestamp 1698175906
transform 1 0 21616 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_211
timestamp 1698175906
transform 1 0 24976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_215
timestamp 1698175906
transform 1 0 25424 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_231
timestamp 1698175906
transform 1 0 27216 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_239
timestamp 1698175906
transform 1 0 28112 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_243
timestamp 1698175906
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_104
timestamp 1698175906
transform 1 0 12992 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_120
timestamp 1698175906
transform 1 0 14784 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_128
timestamp 1698175906
transform 1 0 15680 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_135
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698175906
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_150
timestamp 1698175906
transform 1 0 18144 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_154
timestamp 1698175906
transform 1 0 18592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_156
timestamp 1698175906
transform 1 0 18816 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_167
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_177
timestamp 1698175906
transform 1 0 21168 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_216
timestamp 1698175906
transform 1 0 25536 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_220
timestamp 1698175906
transform 1 0 25984 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_252
timestamp 1698175906
transform 1 0 29568 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_268
timestamp 1698175906
transform 1 0 31360 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_131
timestamp 1698175906
transform 1 0 16016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_135
timestamp 1698175906
transform 1 0 16464 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_179
timestamp 1698175906
transform 1 0 21392 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_205
timestamp 1698175906
transform 1 0 24304 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_237
timestamp 1698175906
transform 1 0 27888 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_88
timestamp 1698175906
transform 1 0 11200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_119
timestamp 1698175906
transform 1 0 14672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_123
timestamp 1698175906
transform 1 0 15120 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698175906
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_150
timestamp 1698175906
transform 1 0 18144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_152
timestamp 1698175906
transform 1 0 18368 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_159
timestamp 1698175906
transform 1 0 19152 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_169
timestamp 1698175906
transform 1 0 20272 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_185
timestamp 1698175906
transform 1 0 22064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_195
timestamp 1698175906
transform 1 0 23184 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_199
timestamp 1698175906
transform 1 0 23632 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698175906
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_69
timestamp 1698175906
transform 1 0 9072 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_85
timestamp 1698175906
transform 1 0 10864 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_93
timestamp 1698175906
transform 1 0 11760 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_97
timestamp 1698175906
transform 1 0 12208 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_129
timestamp 1698175906
transform 1 0 15792 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_137
timestamp 1698175906
transform 1 0 16688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_139
timestamp 1698175906
transform 1 0 16912 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_158
timestamp 1698175906
transform 1 0 19040 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698175906
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_193
timestamp 1698175906
transform 1 0 22960 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_195
timestamp 1698175906
transform 1 0 23184 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_227
timestamp 1698175906
transform 1 0 26768 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_109
timestamp 1698175906
transform 1 0 13552 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_119
timestamp 1698175906
transform 1 0 14672 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_123
timestamp 1698175906
transform 1 0 15120 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698175906
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698175906
transform 1 0 24528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_228
timestamp 1698175906
transform 1 0 26880 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_240
timestamp 1698175906
transform 1 0 28224 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_272
timestamp 1698175906
transform 1 0 31808 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_129
timestamp 1698175906
transform 1 0 15792 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_131
timestamp 1698175906
transform 1 0 16016 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_158
timestamp 1698175906
transform 1 0 19040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_160
timestamp 1698175906
transform 1 0 19264 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_167
timestamp 1698175906
transform 1 0 20048 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_205
timestamp 1698175906
transform 1 0 24304 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_213
timestamp 1698175906
transform 1 0 25200 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_104
timestamp 1698175906
transform 1 0 12992 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_108
timestamp 1698175906
transform 1 0 13440 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_110
timestamp 1698175906
transform 1 0 13664 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_156
timestamp 1698175906
transform 1 0 18816 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_168
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_201
timestamp 1698175906
transform 1 0 23856 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_216
timestamp 1698175906
transform 1 0 25536 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_248
timestamp 1698175906
transform 1 0 29120 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 9072 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698175906
transform 1 0 9520 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_75
timestamp 1698175906
transform 1 0 9744 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_111
timestamp 1698175906
transform 1 0 13776 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_119
timestamp 1698175906
transform 1 0 14672 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_123
timestamp 1698175906
transform 1 0 15120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_152
timestamp 1698175906
transform 1 0 18368 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_154
timestamp 1698175906
transform 1 0 18592 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698175906
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_217
timestamp 1698175906
transform 1 0 25648 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698175906
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 4480 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 8064 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_104
timestamp 1698175906
transform 1 0 12992 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_117
timestamp 1698175906
transform 1 0 14448 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_125
timestamp 1698175906
transform 1 0 15344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_127
timestamp 1698175906
transform 1 0 15568 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_134
timestamp 1698175906
transform 1 0 16352 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_138
timestamp 1698175906
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_158
timestamp 1698175906
transform 1 0 19040 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_184
timestamp 1698175906
transform 1 0 21952 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_196
timestamp 1698175906
transform 1 0 23296 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_204
timestamp 1698175906
transform 1 0 24192 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_208
timestamp 1698175906
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698175906
transform 1 0 32256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 40320 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 9072 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 9520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 9744 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_117
timestamp 1698175906
transform 1 0 14448 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_125
timestamp 1698175906
transform 1 0 15344 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_129
timestamp 1698175906
transform 1 0 15792 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_146
timestamp 1698175906
transform 1 0 17696 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_154
timestamp 1698175906
transform 1 0 18592 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_170
timestamp 1698175906
transform 1 0 20384 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698175906
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_181
timestamp 1698175906
transform 1 0 21616 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_194
timestamp 1698175906
transform 1 0 23072 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_210
timestamp 1698175906
transform 1 0 24864 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_212
timestamp 1698175906
transform 1 0 25088 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_219
timestamp 1698175906
transform 1 0 25872 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_226
timestamp 1698175906
transform 1 0 26656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_228
timestamp 1698175906
transform 1 0 26880 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_234
timestamp 1698175906
transform 1 0 27552 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1698175906
transform 1 0 28448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 4480 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 8064 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_104
timestamp 1698175906
transform 1 0 12992 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_113
timestamp 1698175906
transform 1 0 14000 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_121
timestamp 1698175906
transform 1 0 14896 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_148
timestamp 1698175906
transform 1 0 17920 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_202
timestamp 1698175906
transform 1 0 23968 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_245
timestamp 1698175906
transform 1 0 28784 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698175906
transform 1 0 32368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 40096 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 40320 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_115
timestamp 1698175906
transform 1 0 14224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_125
timestamp 1698175906
transform 1 0 15344 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_149
timestamp 1698175906
transform 1 0 18032 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_157
timestamp 1698175906
transform 1 0 18928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_164
timestamp 1698175906
transform 1 0 19712 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698175906
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_189
timestamp 1698175906
transform 1 0 22512 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_191
timestamp 1698175906
transform 1 0 22736 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_196
timestamp 1698175906
transform 1 0 23296 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_212
timestamp 1698175906
transform 1 0 25088 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_220
timestamp 1698175906
transform 1 0 25984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_222
timestamp 1698175906
transform 1 0 26208 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_228
timestamp 1698175906
transform 1 0 26880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_235
timestamp 1698175906
transform 1 0 27664 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698175906
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_117
timestamp 1698175906
transform 1 0 14448 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_121
timestamp 1698175906
transform 1 0 14896 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698175906
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_149
timestamp 1698175906
transform 1 0 18032 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_153
timestamp 1698175906
transform 1 0 18480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_170
timestamp 1698175906
transform 1 0 20384 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_203
timestamp 1698175906
transform 1 0 24080 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698175906
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_214
timestamp 1698175906
transform 1 0 25312 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_246
timestamp 1698175906
transform 1 0 28896 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698175906
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_115
timestamp 1698175906
transform 1 0 14224 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_119
timestamp 1698175906
transform 1 0 14672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_130
timestamp 1698175906
transform 1 0 15904 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_134
timestamp 1698175906
transform 1 0 16352 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_146
timestamp 1698175906
transform 1 0 17696 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_162
timestamp 1698175906
transform 1 0 19488 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698175906
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_211
timestamp 1698175906
transform 1 0 24976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_215
timestamp 1698175906
transform 1 0 25424 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_231
timestamp 1698175906
transform 1 0 27216 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_239
timestamp 1698175906
transform 1 0 28112 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_88
timestamp 1698175906
transform 1 0 11200 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_96
timestamp 1698175906
transform 1 0 12096 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_100
timestamp 1698175906
transform 1 0 12544 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_146
timestamp 1698175906
transform 1 0 17696 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_205
timestamp 1698175906
transform 1 0 24304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698175906
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_226
timestamp 1698175906
transform 1 0 26656 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_258
timestamp 1698175906
transform 1 0 30240 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_274
timestamp 1698175906
transform 1 0 32032 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698175906
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 36512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 37408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_127
timestamp 1698175906
transform 1 0 15568 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_136
timestamp 1698175906
transform 1 0 16576 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_140
timestamp 1698175906
transform 1 0 17024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_142
timestamp 1698175906
transform 1 0 17248 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698175906
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_179
timestamp 1698175906
transform 1 0 21392 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_190
timestamp 1698175906
transform 1 0 22624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_192
timestamp 1698175906
transform 1 0 22848 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_222
timestamp 1698175906
transform 1 0 26208 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_238
timestamp 1698175906
transform 1 0 28000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698175906
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 4480 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_80
timestamp 1698175906
transform 1 0 10304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_84
timestamp 1698175906
transform 1 0 10752 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_115
timestamp 1698175906
transform 1 0 14224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_119
timestamp 1698175906
transform 1 0 14672 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_127
timestamp 1698175906
transform 1 0 15568 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_131
timestamp 1698175906
transform 1 0 16016 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_133
timestamp 1698175906
transform 1 0 16240 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_158
timestamp 1698175906
transform 1 0 19040 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_166
timestamp 1698175906
transform 1 0 19936 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_170
timestamp 1698175906
transform 1 0 20384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_174
timestamp 1698175906
transform 1 0 20832 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_178
timestamp 1698175906
transform 1 0 21280 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_180
timestamp 1698175906
transform 1 0 21504 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_193
timestamp 1698175906
transform 1 0 22960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_195
timestamp 1698175906
transform 1 0 23184 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_204
timestamp 1698175906
transform 1 0 24192 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698175906
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_115
timestamp 1698175906
transform 1 0 14224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_119
timestamp 1698175906
transform 1 0 14672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_149
timestamp 1698175906
transform 1 0 18032 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_153
timestamp 1698175906
transform 1 0 18480 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_169
timestamp 1698175906
transform 1 0 20272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698175906
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_186
timestamp 1698175906
transform 1 0 22176 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_188
timestamp 1698175906
transform 1 0 22400 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_220
timestamp 1698175906
transform 1 0 25984 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_236
timestamp 1698175906
transform 1 0 27776 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_104
timestamp 1698175906
transform 1 0 12992 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_120
timestamp 1698175906
transform 1 0 14784 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_128
timestamp 1698175906
transform 1 0 15680 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_132
timestamp 1698175906
transform 1 0 16128 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_134
timestamp 1698175906
transform 1 0 16352 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_149
timestamp 1698175906
transform 1 0 18032 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_156
timestamp 1698175906
transform 1 0 18816 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_160
timestamp 1698175906
transform 1 0 19264 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_196
timestamp 1698175906
transform 1 0 23296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_198
timestamp 1698175906
transform 1 0 23520 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_123
timestamp 1698175906
transform 1 0 15120 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_131
timestamp 1698175906
transform 1 0 16016 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_161
timestamp 1698175906
transform 1 0 19376 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_165
timestamp 1698175906
transform 1 0 19824 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_173
timestamp 1698175906
transform 1 0 20720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_181
timestamp 1698175906
transform 1 0 21616 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_189
timestamp 1698175906
transform 1 0 22512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_192
timestamp 1698175906
transform 1 0 22848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_224
timestamp 1698175906
transform 1 0 26432 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_240
timestamp 1698175906
transform 1 0 28224 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698175906
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_6
timestamp 1698175906
transform 1 0 2016 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_22
timestamp 1698175906
transform 1 0 3808 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_30
timestamp 1698175906
transform 1 0 4704 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_203
timestamp 1698175906
transform 1 0 24080 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_215
timestamp 1698175906
transform 1 0 25424 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_243
timestamp 1698175906
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_150
timestamp 1698175906
transform 1 0 18144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_154
timestamp 1698175906
transform 1 0 18592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 28000 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 31584 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita39_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 25424 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita39_26
timestamp 1698175906
transform -1 0 2016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17472 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 18704 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 37520 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 20272 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 27328 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 21616 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 37520 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 25648 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 24976 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform -1 0 4480 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 4480 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform -1 0 4480 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 24192 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 20944 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 24864 41200 24976 42000 0 FreeSans 448 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 18816 41200 18928 42000 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 20160 41200 20272 42000 0 FreeSans 448 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 41200 24192 42000 24304 0 FreeSans 448 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 0 35616 800 35728 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 23520 41200 23632 42000 0 FreeSans 448 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 21504 41200 21616 42000 0 FreeSans 448 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 41200 18816 42000 18928 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 25536 41200 25648 42000 0 FreeSans 448 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 17472 41200 17584 42000 0 FreeSans 448 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 24192 41200 24304 42000 0 FreeSans 448 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 41200 21504 42000 21616 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal3 13440 22456 13440 22456 0 _000_
rlabel metal2 24696 19600 24696 19600 0 _001_
rlabel metal2 12152 19544 12152 19544 0 _002_
rlabel metal2 15960 25872 15960 25872 0 _003_
rlabel metal2 26600 22792 26600 22792 0 _004_
rlabel metal2 23688 27496 23688 27496 0 _005_
rlabel metal2 14952 24304 14952 24304 0 _006_
rlabel metal2 16072 26936 16072 26936 0 _007_
rlabel metal2 18424 13496 18424 13496 0 _008_
rlabel metal2 15176 13440 15176 13440 0 _009_
rlabel metal2 24472 16800 24472 16800 0 _010_
rlabel metal2 20328 28168 20328 28168 0 _011_
rlabel metal2 22680 24248 22680 24248 0 _012_
rlabel metal2 23856 25592 23856 25592 0 _013_
rlabel metal2 22624 15288 22624 15288 0 _014_
rlabel metal2 12152 20608 12152 20608 0 _015_
rlabel metal2 27608 18760 27608 18760 0 _016_
rlabel metal2 26544 17752 26544 17752 0 _017_
rlabel metal2 22568 14056 22568 14056 0 _018_
rlabel metal3 17416 27608 17416 27608 0 _019_
rlabel metal2 18256 24920 18256 24920 0 _020_
rlabel metal2 22008 22736 22008 22736 0 _021_
rlabel metal2 18648 14840 18648 14840 0 _022_
rlabel metal2 26376 21224 26376 21224 0 _023_
rlabel metal3 12880 17416 12880 17416 0 _024_
rlabel metal2 12600 16016 12600 16016 0 _025_
rlabel metal2 17304 23576 17304 23576 0 _026_
rlabel metal2 14672 25480 14672 25480 0 _027_
rlabel metal2 15064 24864 15064 24864 0 _028_
rlabel metal2 15736 25536 15736 25536 0 _029_
rlabel metal2 21336 23688 21336 23688 0 _030_
rlabel metal2 26936 22232 26936 22232 0 _031_
rlabel metal2 17752 16800 17752 16800 0 _032_
rlabel metal3 21672 18368 21672 18368 0 _033_
rlabel metal3 22904 23688 22904 23688 0 _034_
rlabel metal2 22008 27440 22008 27440 0 _035_
rlabel metal2 24024 27720 24024 27720 0 _036_
rlabel metal2 16072 25200 16072 25200 0 _037_
rlabel metal2 15624 24080 15624 24080 0 _038_
rlabel metal2 16744 26992 16744 26992 0 _039_
rlabel metal2 19768 12376 19768 12376 0 _040_
rlabel metal3 17752 16856 17752 16856 0 _041_
rlabel metal2 19320 13944 19320 13944 0 _042_
rlabel metal2 17640 17304 17640 17304 0 _043_
rlabel metal2 17304 15288 17304 15288 0 _044_
rlabel metal2 17416 14224 17416 14224 0 _045_
rlabel metal2 16296 14056 16296 14056 0 _046_
rlabel metal2 24360 15904 24360 15904 0 _047_
rlabel metal2 23576 17696 23576 17696 0 _048_
rlabel metal2 21672 27832 21672 27832 0 _049_
rlabel metal2 22848 14728 22848 14728 0 _050_
rlabel metal3 23912 24920 23912 24920 0 _051_
rlabel metal2 23352 26376 23352 26376 0 _052_
rlabel metal2 14280 20412 14280 20412 0 _053_
rlabel metal3 22568 14504 22568 14504 0 _054_
rlabel metal3 23352 14616 23352 14616 0 _055_
rlabel metal2 13552 20216 13552 20216 0 _056_
rlabel metal2 28000 19208 28000 19208 0 _057_
rlabel metal2 27496 19432 27496 19432 0 _058_
rlabel metal2 26264 18872 26264 18872 0 _059_
rlabel metal2 26712 18032 26712 18032 0 _060_
rlabel metal3 22960 18984 22960 18984 0 _061_
rlabel metal3 24304 13832 24304 13832 0 _062_
rlabel metal2 18032 28056 18032 28056 0 _063_
rlabel metal2 17640 27356 17640 27356 0 _064_
rlabel metal2 19880 24472 19880 24472 0 _065_
rlabel metal2 14392 17304 14392 17304 0 _066_
rlabel metal2 16912 20888 16912 20888 0 _067_
rlabel metal2 14840 16016 14840 16016 0 _068_
rlabel metal2 15960 20384 15960 20384 0 _069_
rlabel metal2 21560 23576 21560 23576 0 _070_
rlabel metal2 21896 18872 21896 18872 0 _071_
rlabel metal2 19544 17192 19544 17192 0 _072_
rlabel metal3 18872 20104 18872 20104 0 _073_
rlabel metal2 22400 20664 22400 20664 0 _074_
rlabel metal2 13496 19992 13496 19992 0 _075_
rlabel metal2 20888 22344 20888 22344 0 _076_
rlabel metal2 19376 22344 19376 22344 0 _077_
rlabel metal2 22064 22232 22064 22232 0 _078_
rlabel metal2 22400 22120 22400 22120 0 _079_
rlabel metal2 16408 16856 16408 16856 0 _080_
rlabel metal2 21448 20104 21448 20104 0 _081_
rlabel metal2 13720 20160 13720 20160 0 _082_
rlabel metal2 16632 21168 16632 21168 0 _083_
rlabel metal2 24024 14784 24024 14784 0 _084_
rlabel metal2 21672 14504 21672 14504 0 _085_
rlabel metal3 18872 16632 18872 16632 0 _086_
rlabel metal2 20216 14112 20216 14112 0 _087_
rlabel metal2 16408 18144 16408 18144 0 _088_
rlabel metal2 16296 21392 16296 21392 0 _089_
rlabel metal2 19768 18984 19768 18984 0 _090_
rlabel metal2 20104 15456 20104 15456 0 _091_
rlabel metal3 16576 21784 16576 21784 0 _092_
rlabel metal2 14616 21840 14616 21840 0 _093_
rlabel metal2 22680 17976 22680 17976 0 _094_
rlabel metal3 22288 26936 22288 26936 0 _095_
rlabel metal3 24696 20664 24696 20664 0 _096_
rlabel metal2 25256 25536 25256 25536 0 _097_
rlabel metal2 27440 20776 27440 20776 0 _098_
rlabel metal2 26768 20664 26768 20664 0 _099_
rlabel metal2 13216 15960 13216 15960 0 _100_
rlabel metal2 14896 22344 14896 22344 0 _101_
rlabel metal2 15904 22344 15904 22344 0 _102_
rlabel metal2 20272 23688 20272 23688 0 _103_
rlabel metal2 17416 18816 17416 18816 0 _104_
rlabel metal3 15400 19208 15400 19208 0 _105_
rlabel metal3 2478 27608 2478 27608 0 clk
rlabel metal3 19880 21448 19880 21448 0 clknet_0_clk
rlabel metal2 21784 13832 21784 13832 0 clknet_1_0__leaf_clk
rlabel metal2 13160 21112 13160 21112 0 clknet_1_1__leaf_clk
rlabel metal2 14168 16464 14168 16464 0 dut39.count\[0\]
rlabel metal3 14784 15512 14784 15512 0 dut39.count\[1\]
rlabel metal2 14280 22344 14280 22344 0 dut39.count\[2\]
rlabel metal2 22120 19152 22120 19152 0 dut39.count\[3\]
rlabel metal2 17752 5964 17752 5964 0 net1
rlabel metal2 28616 18088 28616 18088 0 net10
rlabel metal2 26040 25984 26040 25984 0 net11
rlabel metal3 25480 13608 25480 13608 0 net12
rlabel metal2 17864 27440 17864 27440 0 net13
rlabel metal2 24584 5964 24584 5964 0 net14
rlabel metal3 11648 20888 11648 20888 0 net15
rlabel metal2 12824 25032 12824 25032 0 net16
rlabel metal3 25144 28056 25144 28056 0 net17
rlabel metal2 28728 23128 28728 23128 0 net18
rlabel metal3 6356 26264 6356 26264 0 net19
rlabel metal2 25480 9716 25480 9716 0 net2
rlabel metal2 10024 19656 10024 19656 0 net20
rlabel metal2 23128 28280 23128 28280 0 net21
rlabel metal2 28616 21616 28616 21616 0 net22
rlabel metal3 31920 23016 31920 23016 0 net23
rlabel metal2 21112 5964 21112 5964 0 net24
rlabel metal2 25144 37520 25144 37520 0 net25
rlabel metal3 1246 35672 1246 35672 0 net26
rlabel metal2 18536 28392 18536 28392 0 net3
rlabel metal2 20888 31920 20888 31920 0 net4
rlabel metal3 31920 24752 31920 24752 0 net5
rlabel metal2 20496 13048 20496 13048 0 net6
rlabel metal2 27048 31472 27048 31472 0 net7
rlabel metal3 22624 27944 22624 27944 0 net8
rlabel metal2 28952 18760 28952 18760 0 net9
rlabel metal2 17528 2198 17528 2198 0 segm[10]
rlabel metal2 24248 2422 24248 2422 0 segm[11]
rlabel metal3 19376 37464 19376 37464 0 segm[12]
rlabel metal2 20216 38962 20216 38962 0 segm[13]
rlabel metal2 40040 24360 40040 24360 0 segm[1]
rlabel metal2 20216 2422 20216 2422 0 segm[2]
rlabel metal3 24192 38248 24192 38248 0 segm[4]
rlabel metal2 21560 39354 21560 39354 0 segm[5]
rlabel metal2 40040 19096 40040 19096 0 segm[6]
rlabel metal3 40642 18200 40642 18200 0 segm[7]
rlabel metal2 25592 38962 25592 38962 0 segm[8]
rlabel metal2 24920 2982 24920 2982 0 segm[9]
rlabel metal2 17528 39746 17528 39746 0 sel[0]
rlabel metal2 23576 2198 23576 2198 0 sel[10]
rlabel metal3 1358 20888 1358 20888 0 sel[11]
rlabel metal3 1414 24920 1414 24920 0 sel[1]
rlabel metal2 24248 39354 24248 39354 0 sel[2]
rlabel metal2 40040 23800 40040 23800 0 sel[3]
rlabel metal3 1358 25592 1358 25592 0 sel[4]
rlabel metal3 1358 19544 1358 19544 0 sel[5]
rlabel metal2 22232 39690 22232 39690 0 sel[6]
rlabel metal2 40040 22008 40040 22008 0 sel[7]
rlabel metal3 40642 22904 40642 22904 0 sel[8]
rlabel metal2 20888 2198 20888 2198 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
