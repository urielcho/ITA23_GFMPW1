magic
tech gf180mcuD
magscale 1 10
timestamp 1699641927
<< metal1 >>
rect 17266 38558 17278 38610
rect 17330 38607 17342 38610
rect 18162 38607 18174 38610
rect 17330 38561 18174 38607
rect 17330 38558 17342 38561
rect 18162 38558 18174 38561
rect 18226 38558 18238 38610
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 18622 38274 18674 38286
rect 18622 38210 18674 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 17826 37998 17838 38050
rect 17890 37998 17902 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 17278 37938 17330 37950
rect 17278 37874 17330 37886
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 18398 37490 18450 37502
rect 18398 37426 18450 37438
rect 17378 37214 17390 37266
rect 17442 37214 17454 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 17378 27806 17390 27858
rect 17442 27806 17454 27858
rect 20626 27806 20638 27858
rect 20690 27806 20702 27858
rect 18286 27746 18338 27758
rect 18286 27682 18338 27694
rect 20414 27746 20466 27758
rect 21410 27694 21422 27746
rect 21474 27694 21486 27746
rect 23538 27694 23550 27746
rect 23602 27694 23614 27746
rect 20414 27682 20466 27694
rect 17390 27634 17442 27646
rect 17390 27570 17442 27582
rect 17726 27634 17778 27646
rect 17726 27570 17778 27582
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 21858 27246 21870 27298
rect 21922 27246 21934 27298
rect 1934 27186 1986 27198
rect 21422 27186 21474 27198
rect 15138 27134 15150 27186
rect 15202 27134 15214 27186
rect 17266 27134 17278 27186
rect 17330 27134 17342 27186
rect 20514 27134 20526 27186
rect 20578 27134 20590 27186
rect 1934 27122 1986 27134
rect 21422 27122 21474 27134
rect 22542 27186 22594 27198
rect 40014 27186 40066 27198
rect 27458 27134 27470 27186
rect 27522 27134 27534 27186
rect 22542 27122 22594 27134
rect 40014 27122 40066 27134
rect 4274 27022 4286 27074
rect 4338 27022 4350 27074
rect 14354 27022 14366 27074
rect 14418 27022 14430 27074
rect 17602 27022 17614 27074
rect 17666 27022 17678 27074
rect 21522 27022 21534 27074
rect 21586 27022 21598 27074
rect 22082 27022 22094 27074
rect 22146 27022 22158 27074
rect 24658 27022 24670 27074
rect 24722 27022 24734 27074
rect 27906 27022 27918 27074
rect 27970 27022 27982 27074
rect 37650 27022 37662 27074
rect 37714 27022 37726 27074
rect 21310 26962 21362 26974
rect 12114 26910 12126 26962
rect 12178 26910 12190 26962
rect 18386 26910 18398 26962
rect 18450 26910 18462 26962
rect 21310 26898 21362 26910
rect 22430 26962 22482 26974
rect 22430 26898 22482 26910
rect 22654 26962 22706 26974
rect 22654 26898 22706 26910
rect 24222 26962 24274 26974
rect 25330 26910 25342 26962
rect 25394 26910 25406 26962
rect 28130 26910 28142 26962
rect 28194 26910 28206 26962
rect 24222 26898 24274 26910
rect 12462 26850 12514 26862
rect 12462 26786 12514 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 17726 26514 17778 26526
rect 17726 26450 17778 26462
rect 17838 26514 17890 26526
rect 17838 26450 17890 26462
rect 18734 26514 18786 26526
rect 18734 26450 18786 26462
rect 18846 26514 18898 26526
rect 20638 26514 20690 26526
rect 19618 26462 19630 26514
rect 19682 26462 19694 26514
rect 18846 26450 18898 26462
rect 20638 26450 20690 26462
rect 25342 26514 25394 26526
rect 25342 26450 25394 26462
rect 26574 26514 26626 26526
rect 26574 26450 26626 26462
rect 17614 26290 17666 26302
rect 18958 26290 19010 26302
rect 4274 26238 4286 26290
rect 4338 26238 4350 26290
rect 13122 26238 13134 26290
rect 13186 26238 13198 26290
rect 13794 26238 13806 26290
rect 13858 26238 13870 26290
rect 17378 26238 17390 26290
rect 17442 26238 17454 26290
rect 18050 26238 18062 26290
rect 18114 26238 18126 26290
rect 18386 26238 18398 26290
rect 18450 26238 18462 26290
rect 17614 26226 17666 26238
rect 18958 26226 19010 26238
rect 19294 26290 19346 26302
rect 19294 26226 19346 26238
rect 21086 26290 21138 26302
rect 25230 26290 25282 26302
rect 21522 26238 21534 26290
rect 21586 26238 21598 26290
rect 21086 26226 21138 26238
rect 25230 26226 25282 26238
rect 25454 26290 25506 26302
rect 25454 26226 25506 26238
rect 25902 26290 25954 26302
rect 25902 26226 25954 26238
rect 26350 26290 26402 26302
rect 26350 26226 26402 26238
rect 26686 26290 26738 26302
rect 37874 26238 37886 26290
rect 37938 26238 37950 26290
rect 26686 26226 26738 26238
rect 10210 26126 10222 26178
rect 10274 26126 10286 26178
rect 12338 26126 12350 26178
rect 12402 26126 12414 26178
rect 14466 26126 14478 26178
rect 14530 26126 14542 26178
rect 16594 26126 16606 26178
rect 16658 26126 16670 26178
rect 22194 26126 22206 26178
rect 22258 26126 22270 26178
rect 24322 26126 24334 26178
rect 24386 26126 24398 26178
rect 39890 26126 39902 26178
rect 39954 26126 39966 26178
rect 1934 26066 1986 26078
rect 1934 26002 1986 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 11678 25730 11730 25742
rect 11678 25666 11730 25678
rect 18398 25730 18450 25742
rect 18398 25666 18450 25678
rect 21758 25730 21810 25742
rect 21758 25666 21810 25678
rect 16046 25618 16098 25630
rect 2034 25566 2046 25618
rect 2098 25566 2110 25618
rect 16930 25566 16942 25618
rect 16994 25566 17006 25618
rect 16046 25554 16098 25566
rect 16158 25506 16210 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 12338 25454 12350 25506
rect 12402 25454 12414 25506
rect 16158 25442 16210 25454
rect 16606 25506 16658 25518
rect 16606 25442 16658 25454
rect 17054 25506 17106 25518
rect 18286 25506 18338 25518
rect 17490 25454 17502 25506
rect 17554 25454 17566 25506
rect 17054 25442 17106 25454
rect 18286 25442 18338 25454
rect 22430 25506 22482 25518
rect 22430 25442 22482 25454
rect 11678 25394 11730 25406
rect 11678 25330 11730 25342
rect 11790 25394 11842 25406
rect 17278 25394 17330 25406
rect 21758 25394 21810 25406
rect 12114 25342 12126 25394
rect 12178 25342 12190 25394
rect 18834 25342 18846 25394
rect 18898 25342 18910 25394
rect 11790 25330 11842 25342
rect 17278 25330 17330 25342
rect 21758 25330 21810 25342
rect 21870 25394 21922 25406
rect 21870 25330 21922 25342
rect 22094 25394 22146 25406
rect 22094 25330 22146 25342
rect 13582 25282 13634 25294
rect 13582 25218 13634 25230
rect 15934 25282 15986 25294
rect 15934 25218 15986 25230
rect 16942 25282 16994 25294
rect 16942 25218 16994 25230
rect 18398 25282 18450 25294
rect 18398 25218 18450 25230
rect 19182 25282 19234 25294
rect 19182 25218 19234 25230
rect 22318 25282 22370 25294
rect 22318 25218 22370 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 12350 24946 12402 24958
rect 12350 24882 12402 24894
rect 12574 24946 12626 24958
rect 12574 24882 12626 24894
rect 16830 24946 16882 24958
rect 22642 24894 22654 24946
rect 22706 24894 22718 24946
rect 16830 24882 16882 24894
rect 20638 24834 20690 24846
rect 19842 24782 19854 24834
rect 19906 24782 19918 24834
rect 20638 24770 20690 24782
rect 21870 24834 21922 24846
rect 22418 24782 22430 24834
rect 22482 24782 22494 24834
rect 26114 24782 26126 24834
rect 26178 24782 26190 24834
rect 21870 24770 21922 24782
rect 12686 24722 12738 24734
rect 25790 24722 25842 24734
rect 20066 24670 20078 24722
rect 20130 24670 20142 24722
rect 22194 24670 22206 24722
rect 22258 24670 22270 24722
rect 12686 24658 12738 24670
rect 25790 24658 25842 24670
rect 21410 24558 21422 24610
rect 21474 24558 21486 24610
rect 20526 24498 20578 24510
rect 20526 24434 20578 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 23886 24162 23938 24174
rect 23886 24098 23938 24110
rect 1934 24050 1986 24062
rect 19070 24050 19122 24062
rect 13458 23998 13470 24050
rect 13522 23998 13534 24050
rect 1934 23986 1986 23998
rect 19070 23986 19122 23998
rect 40014 24050 40066 24062
rect 40014 23986 40066 23998
rect 17502 23938 17554 23950
rect 19854 23938 19906 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 16258 23886 16270 23938
rect 16322 23886 16334 23938
rect 16930 23886 16942 23938
rect 16994 23886 17006 23938
rect 19618 23886 19630 23938
rect 19682 23886 19694 23938
rect 17502 23874 17554 23886
rect 19854 23874 19906 23886
rect 20526 23938 20578 23950
rect 20526 23874 20578 23886
rect 21982 23938 22034 23950
rect 21982 23874 22034 23886
rect 22542 23938 22594 23950
rect 22542 23874 22594 23886
rect 23438 23938 23490 23950
rect 23438 23874 23490 23886
rect 24110 23938 24162 23950
rect 24110 23874 24162 23886
rect 25118 23938 25170 23950
rect 25118 23874 25170 23886
rect 25678 23938 25730 23950
rect 25678 23874 25730 23886
rect 26462 23938 26514 23950
rect 26462 23874 26514 23886
rect 26798 23938 26850 23950
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 26798 23874 26850 23886
rect 24334 23826 24386 23838
rect 15586 23774 15598 23826
rect 15650 23774 15662 23826
rect 20178 23774 20190 23826
rect 20242 23774 20254 23826
rect 24334 23762 24386 23774
rect 24446 23826 24498 23838
rect 24446 23762 24498 23774
rect 24670 23826 24722 23838
rect 24670 23762 24722 23774
rect 25902 23826 25954 23838
rect 25902 23762 25954 23774
rect 25006 23714 25058 23726
rect 16706 23662 16718 23714
rect 16770 23662 16782 23714
rect 23090 23662 23102 23714
rect 23154 23662 23166 23714
rect 25006 23650 25058 23662
rect 25230 23714 25282 23726
rect 25230 23650 25282 23662
rect 26014 23714 26066 23726
rect 26014 23650 26066 23662
rect 26238 23714 26290 23726
rect 26238 23650 26290 23662
rect 26686 23714 26738 23726
rect 26686 23650 26738 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 14926 23378 14978 23390
rect 14926 23314 14978 23326
rect 15374 23378 15426 23390
rect 15374 23314 15426 23326
rect 15486 23378 15538 23390
rect 15486 23314 15538 23326
rect 24670 23378 24722 23390
rect 24670 23314 24722 23326
rect 14254 23266 14306 23278
rect 14254 23202 14306 23214
rect 14366 23266 14418 23278
rect 18722 23214 18734 23266
rect 18786 23214 18798 23266
rect 26002 23214 26014 23266
rect 26066 23214 26078 23266
rect 14366 23202 14418 23214
rect 15710 23154 15762 23166
rect 4274 23102 4286 23154
rect 4338 23102 4350 23154
rect 13794 23102 13806 23154
rect 13858 23102 13870 23154
rect 15922 23102 15934 23154
rect 15986 23102 15998 23154
rect 23090 23102 23102 23154
rect 23154 23102 23166 23154
rect 25218 23102 25230 23154
rect 25282 23102 25294 23154
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 15710 23090 15762 23102
rect 14814 23042 14866 23054
rect 10994 22990 11006 23042
rect 11058 22990 11070 23042
rect 13122 22990 13134 23042
rect 13186 22990 13198 23042
rect 14814 22978 14866 22990
rect 15598 23042 15650 23054
rect 28130 22990 28142 23042
rect 28194 22990 28206 23042
rect 15598 22978 15650 22990
rect 1934 22930 1986 22942
rect 1934 22866 1986 22878
rect 14366 22930 14418 22942
rect 14366 22866 14418 22878
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 15486 22594 15538 22606
rect 15486 22530 15538 22542
rect 1934 22482 1986 22494
rect 1934 22418 1986 22430
rect 14142 22482 14194 22494
rect 14142 22418 14194 22430
rect 17950 22482 18002 22494
rect 17950 22418 18002 22430
rect 19742 22482 19794 22494
rect 23438 22482 23490 22494
rect 20178 22430 20190 22482
rect 20242 22430 20254 22482
rect 19742 22418 19794 22430
rect 23438 22418 23490 22430
rect 24334 22482 24386 22494
rect 25442 22430 25454 22482
rect 25506 22430 25518 22482
rect 27570 22430 27582 22482
rect 27634 22430 27646 22482
rect 24334 22418 24386 22430
rect 15262 22370 15314 22382
rect 4274 22318 4286 22370
rect 4338 22318 4350 22370
rect 15262 22306 15314 22318
rect 17726 22370 17778 22382
rect 18498 22318 18510 22370
rect 18562 22318 18574 22370
rect 19170 22318 19182 22370
rect 19234 22318 19246 22370
rect 20290 22318 20302 22370
rect 20354 22318 20366 22370
rect 21746 22318 21758 22370
rect 21810 22318 21822 22370
rect 24658 22318 24670 22370
rect 24722 22318 24734 22370
rect 17726 22306 17778 22318
rect 15822 22258 15874 22270
rect 18610 22206 18622 22258
rect 18674 22206 18686 22258
rect 22754 22206 22766 22258
rect 22818 22206 22830 22258
rect 15822 22194 15874 22206
rect 15598 22146 15650 22158
rect 23326 22146 23378 22158
rect 17378 22094 17390 22146
rect 17442 22094 17454 22146
rect 19282 22094 19294 22146
rect 19346 22094 19358 22146
rect 21858 22094 21870 22146
rect 21922 22094 21934 22146
rect 15598 22082 15650 22094
rect 23326 22082 23378 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 13918 21810 13970 21822
rect 13918 21746 13970 21758
rect 18062 21810 18114 21822
rect 18062 21746 18114 21758
rect 18174 21810 18226 21822
rect 22094 21810 22146 21822
rect 19618 21758 19630 21810
rect 19682 21758 19694 21810
rect 18174 21746 18226 21758
rect 22094 21746 22146 21758
rect 13358 21698 13410 21710
rect 13358 21634 13410 21646
rect 13470 21698 13522 21710
rect 13470 21634 13522 21646
rect 17838 21698 17890 21710
rect 17838 21634 17890 21646
rect 17950 21698 18002 21710
rect 21758 21698 21810 21710
rect 18946 21646 18958 21698
rect 19010 21646 19022 21698
rect 19170 21646 19182 21698
rect 19234 21646 19246 21698
rect 21634 21646 21646 21698
rect 21698 21646 21710 21698
rect 17950 21634 18002 21646
rect 21758 21634 21810 21646
rect 21870 21698 21922 21710
rect 21870 21634 21922 21646
rect 22318 21698 22370 21710
rect 22978 21646 22990 21698
rect 23042 21646 23054 21698
rect 23202 21646 23214 21698
rect 23266 21646 23278 21698
rect 22318 21634 22370 21646
rect 13134 21586 13186 21598
rect 22542 21586 22594 21598
rect 12898 21534 12910 21586
rect 12962 21534 12974 21586
rect 17490 21534 17502 21586
rect 17554 21534 17566 21586
rect 18610 21534 18622 21586
rect 18674 21534 18686 21586
rect 20514 21534 20526 21586
rect 20578 21534 20590 21586
rect 13134 21522 13186 21534
rect 22542 21522 22594 21534
rect 23998 21586 24050 21598
rect 23998 21522 24050 21534
rect 37326 21586 37378 21598
rect 37762 21534 37774 21586
rect 37826 21534 37838 21586
rect 37326 21522 37378 21534
rect 20974 21474 21026 21486
rect 9986 21422 9998 21474
rect 10050 21422 10062 21474
rect 12114 21422 12126 21474
rect 12178 21422 12190 21474
rect 21746 21422 21758 21474
rect 21810 21422 21822 21474
rect 39890 21422 39902 21474
rect 39954 21422 39966 21474
rect 20974 21410 21026 21422
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 18062 21026 18114 21038
rect 18062 20962 18114 20974
rect 18398 21026 18450 21038
rect 18398 20962 18450 20974
rect 20078 20914 20130 20926
rect 40014 20914 40066 20926
rect 16146 20862 16158 20914
rect 16210 20862 16222 20914
rect 22530 20862 22542 20914
rect 22594 20862 22606 20914
rect 20078 20850 20130 20862
rect 40014 20850 40066 20862
rect 12238 20802 12290 20814
rect 12238 20738 12290 20750
rect 12574 20802 12626 20814
rect 22430 20802 22482 20814
rect 26350 20802 26402 20814
rect 15586 20750 15598 20802
rect 15650 20750 15662 20802
rect 16818 20750 16830 20802
rect 16882 20750 16894 20802
rect 17266 20750 17278 20802
rect 17330 20750 17342 20802
rect 18722 20750 18734 20802
rect 18786 20750 18798 20802
rect 20514 20750 20526 20802
rect 20578 20750 20590 20802
rect 22866 20750 22878 20802
rect 22930 20750 22942 20802
rect 12574 20738 12626 20750
rect 22430 20738 22482 20750
rect 26350 20738 26402 20750
rect 27246 20802 27298 20814
rect 27246 20738 27298 20750
rect 27358 20802 27410 20814
rect 37650 20750 37662 20802
rect 37714 20750 37726 20802
rect 27358 20738 27410 20750
rect 12462 20690 12514 20702
rect 17390 20690 17442 20702
rect 25902 20690 25954 20702
rect 15922 20638 15934 20690
rect 15986 20638 15998 20690
rect 18946 20638 18958 20690
rect 19010 20638 19022 20690
rect 21858 20638 21870 20690
rect 21922 20638 21934 20690
rect 12462 20626 12514 20638
rect 17390 20626 17442 20638
rect 25902 20626 25954 20638
rect 26798 20690 26850 20702
rect 26798 20626 26850 20638
rect 27694 20690 27746 20702
rect 27694 20626 27746 20638
rect 18174 20578 18226 20590
rect 21534 20578 21586 20590
rect 25230 20578 25282 20590
rect 19282 20526 19294 20578
rect 19346 20526 19358 20578
rect 22978 20526 22990 20578
rect 23042 20526 23054 20578
rect 18174 20514 18226 20526
rect 21534 20514 21586 20526
rect 25230 20514 25282 20526
rect 25678 20578 25730 20590
rect 25678 20514 25730 20526
rect 25790 20578 25842 20590
rect 25790 20514 25842 20526
rect 26574 20578 26626 20590
rect 26574 20514 26626 20526
rect 26686 20578 26738 20590
rect 26686 20514 26738 20526
rect 27582 20578 27634 20590
rect 27582 20514 27634 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 16270 20242 16322 20254
rect 16270 20178 16322 20190
rect 15710 20130 15762 20142
rect 13010 20078 13022 20130
rect 13074 20078 13086 20130
rect 15710 20066 15762 20078
rect 15822 20130 15874 20142
rect 28702 20130 28754 20142
rect 16594 20078 16606 20130
rect 16658 20078 16670 20130
rect 26226 20078 26238 20130
rect 26290 20078 26302 20130
rect 15822 20066 15874 20078
rect 28702 20066 28754 20078
rect 28814 20130 28866 20142
rect 28814 20066 28866 20078
rect 17726 20018 17778 20030
rect 12226 19966 12238 20018
rect 12290 19966 12302 20018
rect 17726 19954 17778 19966
rect 18286 20018 18338 20030
rect 18286 19954 18338 19966
rect 18734 20018 18786 20030
rect 19058 19966 19070 20018
rect 19122 19966 19134 20018
rect 25442 19966 25454 20018
rect 25506 19966 25518 20018
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 18734 19954 18786 19966
rect 15138 19854 15150 19906
rect 15202 19854 15214 19906
rect 23090 19854 23102 19906
rect 23154 19854 23166 19906
rect 28354 19854 28366 19906
rect 28418 19854 28430 19906
rect 15822 19794 15874 19806
rect 15822 19730 15874 19742
rect 28814 19794 28866 19806
rect 28814 19730 28866 19742
rect 40014 19794 40066 19806
rect 40014 19730 40066 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 15822 19458 15874 19470
rect 15822 19394 15874 19406
rect 19842 19294 19854 19346
rect 19906 19294 19918 19346
rect 21410 19294 21422 19346
rect 21474 19294 21486 19346
rect 26114 19294 26126 19346
rect 26178 19294 26190 19346
rect 28242 19294 28254 19346
rect 28306 19294 28318 19346
rect 15934 19234 15986 19246
rect 17726 19234 17778 19246
rect 16594 19182 16606 19234
rect 16658 19182 16670 19234
rect 19730 19182 19742 19234
rect 19794 19182 19806 19234
rect 20066 19182 20078 19234
rect 20130 19182 20142 19234
rect 24210 19182 24222 19234
rect 24274 19182 24286 19234
rect 25442 19182 25454 19234
rect 25506 19182 25518 19234
rect 15934 19170 15986 19182
rect 17726 19170 17778 19182
rect 18062 19122 18114 19134
rect 18062 19058 18114 19070
rect 18846 19122 18898 19134
rect 23538 19070 23550 19122
rect 23602 19070 23614 19122
rect 18846 19058 18898 19070
rect 15374 19010 15426 19022
rect 17166 19010 17218 19022
rect 16818 18958 16830 19010
rect 16882 18958 16894 19010
rect 15374 18946 15426 18958
rect 17166 18946 17218 18958
rect 18174 19010 18226 19022
rect 25006 19010 25058 19022
rect 19618 18958 19630 19010
rect 19682 18958 19694 19010
rect 18174 18946 18226 18958
rect 25006 18946 25058 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 15486 18674 15538 18686
rect 15486 18610 15538 18622
rect 23662 18674 23714 18686
rect 23662 18610 23714 18622
rect 18386 18510 18398 18562
rect 18450 18510 18462 18562
rect 19730 18510 19742 18562
rect 19794 18510 19806 18562
rect 20962 18510 20974 18562
rect 21026 18510 21038 18562
rect 16718 18450 16770 18462
rect 22654 18450 22706 18462
rect 12226 18398 12238 18450
rect 12290 18398 12302 18450
rect 16482 18398 16494 18450
rect 16546 18398 16558 18450
rect 17938 18398 17950 18450
rect 18002 18398 18014 18450
rect 19394 18398 19406 18450
rect 19458 18398 19470 18450
rect 21858 18398 21870 18450
rect 21922 18398 21934 18450
rect 22418 18398 22430 18450
rect 22482 18398 22494 18450
rect 16718 18386 16770 18398
rect 22654 18386 22706 18398
rect 22766 18450 22818 18462
rect 23874 18398 23886 18450
rect 23938 18398 23950 18450
rect 22766 18386 22818 18398
rect 15822 18338 15874 18350
rect 12898 18286 12910 18338
rect 12962 18286 12974 18338
rect 15026 18286 15038 18338
rect 15090 18286 15102 18338
rect 15822 18274 15874 18286
rect 23550 18226 23602 18238
rect 23202 18174 23214 18226
rect 23266 18174 23278 18226
rect 23550 18162 23602 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 22094 17890 22146 17902
rect 22094 17826 22146 17838
rect 18174 17778 18226 17790
rect 18174 17714 18226 17726
rect 20638 17778 20690 17790
rect 21870 17778 21922 17790
rect 21522 17726 21534 17778
rect 21586 17726 21598 17778
rect 20638 17714 20690 17726
rect 21870 17714 21922 17726
rect 26014 17778 26066 17790
rect 26014 17714 26066 17726
rect 40014 17778 40066 17790
rect 40014 17714 40066 17726
rect 13806 17666 13858 17678
rect 13806 17602 13858 17614
rect 17726 17666 17778 17678
rect 17726 17602 17778 17614
rect 18622 17666 18674 17678
rect 18622 17602 18674 17614
rect 18958 17666 19010 17678
rect 18958 17602 19010 17614
rect 19742 17666 19794 17678
rect 19742 17602 19794 17614
rect 21646 17666 21698 17678
rect 21646 17602 21698 17614
rect 22318 17666 22370 17678
rect 22318 17602 22370 17614
rect 22542 17666 22594 17678
rect 22542 17602 22594 17614
rect 26126 17666 26178 17678
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 26126 17602 26178 17614
rect 13470 17554 13522 17566
rect 13470 17490 13522 17502
rect 17950 17554 18002 17566
rect 17950 17490 18002 17502
rect 18286 17554 18338 17566
rect 18286 17490 18338 17502
rect 19182 17554 19234 17566
rect 19182 17490 19234 17502
rect 22990 17554 23042 17566
rect 22990 17490 23042 17502
rect 23214 17554 23266 17566
rect 23214 17490 23266 17502
rect 18846 17442 18898 17454
rect 18846 17378 18898 17390
rect 19406 17442 19458 17454
rect 19406 17378 19458 17390
rect 19630 17442 19682 17454
rect 19630 17378 19682 17390
rect 20750 17442 20802 17454
rect 20750 17378 20802 17390
rect 21422 17442 21474 17454
rect 21422 17378 21474 17390
rect 22878 17442 22930 17454
rect 22878 17378 22930 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 18510 17106 18562 17118
rect 18510 17042 18562 17054
rect 18734 17106 18786 17118
rect 18734 17042 18786 17054
rect 14690 16942 14702 16994
rect 14754 16942 14766 16994
rect 17502 16882 17554 16894
rect 14018 16830 14030 16882
rect 14082 16830 14094 16882
rect 17502 16818 17554 16830
rect 19070 16882 19122 16894
rect 23090 16830 23102 16882
rect 23154 16830 23166 16882
rect 19070 16818 19122 16830
rect 16818 16718 16830 16770
rect 16882 16718 16894 16770
rect 19506 16718 19518 16770
rect 19570 16718 19582 16770
rect 18846 16658 18898 16670
rect 18846 16594 18898 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 17826 16158 17838 16210
rect 17890 16158 17902 16210
rect 24770 16158 24782 16210
rect 24834 16158 24846 16210
rect 26898 16158 26910 16210
rect 26962 16158 26974 16210
rect 18286 16098 18338 16110
rect 20750 16098 20802 16110
rect 17938 16046 17950 16098
rect 18002 16046 18014 16098
rect 18946 16046 18958 16098
rect 19010 16046 19022 16098
rect 21634 16046 21646 16098
rect 21698 16046 21710 16098
rect 22754 16046 22766 16098
rect 22818 16046 22830 16098
rect 23986 16046 23998 16098
rect 24050 16046 24062 16098
rect 18286 16034 18338 16046
rect 20750 16034 20802 16046
rect 22990 15986 23042 15998
rect 22990 15922 23042 15934
rect 17726 15874 17778 15886
rect 21870 15874 21922 15886
rect 19170 15822 19182 15874
rect 19234 15822 19246 15874
rect 20402 15822 20414 15874
rect 20466 15822 20478 15874
rect 17726 15810 17778 15822
rect 21870 15810 21922 15822
rect 21982 15874 22034 15886
rect 21982 15810 22034 15822
rect 22094 15874 22146 15886
rect 22094 15810 22146 15822
rect 22206 15874 22258 15886
rect 22206 15810 22258 15822
rect 23662 15874 23714 15886
rect 23662 15810 23714 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 19518 15538 19570 15550
rect 19518 15474 19570 15486
rect 21758 15538 21810 15550
rect 21758 15474 21810 15486
rect 18174 15426 18226 15438
rect 18174 15362 18226 15374
rect 18510 15426 18562 15438
rect 18510 15362 18562 15374
rect 18846 15426 18898 15438
rect 22542 15426 22594 15438
rect 21410 15374 21422 15426
rect 21474 15374 21486 15426
rect 18846 15362 18898 15374
rect 22542 15362 22594 15374
rect 22766 15426 22818 15438
rect 22766 15362 22818 15374
rect 25230 15426 25282 15438
rect 25554 15374 25566 15426
rect 25618 15374 25630 15426
rect 25230 15362 25282 15374
rect 17614 15314 17666 15326
rect 17614 15250 17666 15262
rect 17726 15314 17778 15326
rect 17726 15250 17778 15262
rect 17838 15314 17890 15326
rect 17838 15250 17890 15262
rect 19070 15314 19122 15326
rect 19070 15250 19122 15262
rect 22430 15314 22482 15326
rect 22430 15250 22482 15262
rect 18622 15202 18674 15214
rect 18622 15138 18674 15150
rect 19170 15038 19182 15090
rect 19234 15087 19246 15090
rect 19618 15087 19630 15090
rect 19234 15041 19630 15087
rect 19234 15038 19246 15041
rect 19618 15038 19630 15041
rect 19682 15038 19694 15090
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 21534 14642 21586 14654
rect 16706 14590 16718 14642
rect 16770 14590 16782 14642
rect 18834 14590 18846 14642
rect 18898 14590 18910 14642
rect 23538 14590 23550 14642
rect 23602 14590 23614 14642
rect 25666 14590 25678 14642
rect 25730 14590 25742 14642
rect 21534 14578 21586 14590
rect 19518 14530 19570 14542
rect 16034 14478 16046 14530
rect 16098 14478 16110 14530
rect 19282 14478 19294 14530
rect 19346 14478 19358 14530
rect 19518 14466 19570 14478
rect 19854 14530 19906 14542
rect 21870 14530 21922 14542
rect 20402 14478 20414 14530
rect 20466 14478 20478 14530
rect 19854 14466 19906 14478
rect 21870 14466 21922 14478
rect 22318 14530 22370 14542
rect 22754 14478 22766 14530
rect 22818 14478 22830 14530
rect 22318 14466 22370 14478
rect 22206 14418 22258 14430
rect 22206 14354 22258 14366
rect 19630 14306 19682 14318
rect 19630 14242 19682 14254
rect 19742 14306 19794 14318
rect 22094 14306 22146 14318
rect 20626 14254 20638 14306
rect 20690 14254 20702 14306
rect 19742 14242 19794 14254
rect 22094 14242 22146 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 17502 13970 17554 13982
rect 17502 13906 17554 13918
rect 18958 13970 19010 13982
rect 18958 13906 19010 13918
rect 19070 13970 19122 13982
rect 19070 13906 19122 13918
rect 24558 13970 24610 13982
rect 24558 13906 24610 13918
rect 18734 13858 18786 13870
rect 14690 13806 14702 13858
rect 14754 13806 14766 13858
rect 18734 13794 18786 13806
rect 19742 13858 19794 13870
rect 19742 13794 19794 13806
rect 19182 13746 19234 13758
rect 20078 13746 20130 13758
rect 14018 13694 14030 13746
rect 14082 13694 14094 13746
rect 19394 13694 19406 13746
rect 19458 13694 19470 13746
rect 19182 13682 19234 13694
rect 20078 13682 20130 13694
rect 20302 13746 20354 13758
rect 21186 13694 21198 13746
rect 21250 13694 21262 13746
rect 20302 13682 20354 13694
rect 20190 13634 20242 13646
rect 16818 13582 16830 13634
rect 16882 13582 16894 13634
rect 21970 13582 21982 13634
rect 22034 13582 22046 13634
rect 24098 13582 24110 13634
rect 24162 13582 24174 13634
rect 20190 13570 20242 13582
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 21758 13074 21810 13086
rect 18498 13022 18510 13074
rect 18562 13022 18574 13074
rect 20626 13022 20638 13074
rect 20690 13022 20702 13074
rect 21758 13010 21810 13022
rect 21534 12962 21586 12974
rect 17714 12910 17726 12962
rect 17778 12910 17790 12962
rect 21534 12898 21586 12910
rect 21870 12962 21922 12974
rect 21870 12898 21922 12910
rect 22094 12962 22146 12974
rect 22094 12898 22146 12910
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 20974 12402 21026 12414
rect 20974 12338 21026 12350
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 18734 5234 18786 5246
rect 18734 5170 18786 5182
rect 24782 5234 24834 5246
rect 24782 5170 24834 5182
rect 17826 5070 17838 5122
rect 17890 5070 17902 5122
rect 23762 5070 23774 5122
rect 23826 5070 23838 5122
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 17490 4286 17502 4338
rect 17554 4286 17566 4338
rect 20402 4286 20414 4338
rect 20466 4286 20478 4338
rect 25778 4286 25790 4338
rect 25842 4286 25854 4338
rect 18510 4114 18562 4126
rect 18510 4050 18562 4062
rect 21422 4114 21474 4126
rect 21422 4050 21474 4062
rect 26798 4114 26850 4126
rect 26798 4050 26850 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 22094 3666 22146 3678
rect 18834 3614 18846 3666
rect 18898 3614 18910 3666
rect 22094 3602 22146 3614
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 19730 3502 19742 3554
rect 19794 3502 19806 3554
rect 21074 3502 21086 3554
rect 21138 3502 21150 3554
rect 24994 3502 25006 3554
rect 25058 3502 25070 3554
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 17278 38558 17330 38610
rect 18174 38558 18226 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 18622 38222 18674 38274
rect 25566 38222 25618 38274
rect 17838 37998 17890 38050
rect 24558 37998 24610 38050
rect 17278 37886 17330 37938
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 18398 37438 18450 37490
rect 17390 37214 17442 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 17390 27806 17442 27858
rect 20638 27806 20690 27858
rect 18286 27694 18338 27746
rect 20414 27694 20466 27746
rect 21422 27694 21474 27746
rect 23550 27694 23602 27746
rect 17390 27582 17442 27634
rect 17726 27582 17778 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 21870 27246 21922 27298
rect 1934 27134 1986 27186
rect 15150 27134 15202 27186
rect 17278 27134 17330 27186
rect 20526 27134 20578 27186
rect 21422 27134 21474 27186
rect 22542 27134 22594 27186
rect 27470 27134 27522 27186
rect 40014 27134 40066 27186
rect 4286 27022 4338 27074
rect 14366 27022 14418 27074
rect 17614 27022 17666 27074
rect 21534 27022 21586 27074
rect 22094 27022 22146 27074
rect 24670 27022 24722 27074
rect 27918 27022 27970 27074
rect 37662 27022 37714 27074
rect 12126 26910 12178 26962
rect 18398 26910 18450 26962
rect 21310 26910 21362 26962
rect 22430 26910 22482 26962
rect 22654 26910 22706 26962
rect 24222 26910 24274 26962
rect 25342 26910 25394 26962
rect 28142 26910 28194 26962
rect 12462 26798 12514 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 17726 26462 17778 26514
rect 17838 26462 17890 26514
rect 18734 26462 18786 26514
rect 18846 26462 18898 26514
rect 19630 26462 19682 26514
rect 20638 26462 20690 26514
rect 25342 26462 25394 26514
rect 26574 26462 26626 26514
rect 4286 26238 4338 26290
rect 13134 26238 13186 26290
rect 13806 26238 13858 26290
rect 17390 26238 17442 26290
rect 17614 26238 17666 26290
rect 18062 26238 18114 26290
rect 18398 26238 18450 26290
rect 18958 26238 19010 26290
rect 19294 26238 19346 26290
rect 21086 26238 21138 26290
rect 21534 26238 21586 26290
rect 25230 26238 25282 26290
rect 25454 26238 25506 26290
rect 25902 26238 25954 26290
rect 26350 26238 26402 26290
rect 26686 26238 26738 26290
rect 37886 26238 37938 26290
rect 10222 26126 10274 26178
rect 12350 26126 12402 26178
rect 14478 26126 14530 26178
rect 16606 26126 16658 26178
rect 22206 26126 22258 26178
rect 24334 26126 24386 26178
rect 39902 26126 39954 26178
rect 1934 26014 1986 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 11678 25678 11730 25730
rect 18398 25678 18450 25730
rect 21758 25678 21810 25730
rect 2046 25566 2098 25618
rect 16046 25566 16098 25618
rect 16942 25566 16994 25618
rect 4286 25454 4338 25506
rect 12350 25454 12402 25506
rect 16158 25454 16210 25506
rect 16606 25454 16658 25506
rect 17054 25454 17106 25506
rect 17502 25454 17554 25506
rect 18286 25454 18338 25506
rect 22430 25454 22482 25506
rect 11678 25342 11730 25394
rect 11790 25342 11842 25394
rect 12126 25342 12178 25394
rect 17278 25342 17330 25394
rect 18846 25342 18898 25394
rect 21758 25342 21810 25394
rect 21870 25342 21922 25394
rect 22094 25342 22146 25394
rect 13582 25230 13634 25282
rect 15934 25230 15986 25282
rect 16942 25230 16994 25282
rect 18398 25230 18450 25282
rect 19182 25230 19234 25282
rect 22318 25230 22370 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 12350 24894 12402 24946
rect 12574 24894 12626 24946
rect 16830 24894 16882 24946
rect 22654 24894 22706 24946
rect 19854 24782 19906 24834
rect 20638 24782 20690 24834
rect 21870 24782 21922 24834
rect 22430 24782 22482 24834
rect 26126 24782 26178 24834
rect 12686 24670 12738 24722
rect 20078 24670 20130 24722
rect 22206 24670 22258 24722
rect 25790 24670 25842 24722
rect 21422 24558 21474 24610
rect 20526 24446 20578 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 23886 24110 23938 24162
rect 1934 23998 1986 24050
rect 13470 23998 13522 24050
rect 19070 23998 19122 24050
rect 40014 23998 40066 24050
rect 4286 23886 4338 23938
rect 16270 23886 16322 23938
rect 16942 23886 16994 23938
rect 17502 23886 17554 23938
rect 19630 23886 19682 23938
rect 19854 23886 19906 23938
rect 20526 23886 20578 23938
rect 21982 23886 22034 23938
rect 22542 23886 22594 23938
rect 23438 23886 23490 23938
rect 24110 23886 24162 23938
rect 25118 23886 25170 23938
rect 25678 23886 25730 23938
rect 26462 23886 26514 23938
rect 26798 23886 26850 23938
rect 37662 23886 37714 23938
rect 15598 23774 15650 23826
rect 20190 23774 20242 23826
rect 24334 23774 24386 23826
rect 24446 23774 24498 23826
rect 24670 23774 24722 23826
rect 25902 23774 25954 23826
rect 16718 23662 16770 23714
rect 23102 23662 23154 23714
rect 25006 23662 25058 23714
rect 25230 23662 25282 23714
rect 26014 23662 26066 23714
rect 26238 23662 26290 23714
rect 26686 23662 26738 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 14926 23326 14978 23378
rect 15374 23326 15426 23378
rect 15486 23326 15538 23378
rect 24670 23326 24722 23378
rect 14254 23214 14306 23266
rect 14366 23214 14418 23266
rect 18734 23214 18786 23266
rect 26014 23214 26066 23266
rect 4286 23102 4338 23154
rect 13806 23102 13858 23154
rect 15710 23102 15762 23154
rect 15934 23102 15986 23154
rect 23102 23102 23154 23154
rect 25230 23102 25282 23154
rect 37662 23102 37714 23154
rect 11006 22990 11058 23042
rect 13134 22990 13186 23042
rect 14814 22990 14866 23042
rect 15598 22990 15650 23042
rect 28142 22990 28194 23042
rect 1934 22878 1986 22930
rect 14366 22878 14418 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 15486 22542 15538 22594
rect 1934 22430 1986 22482
rect 14142 22430 14194 22482
rect 17950 22430 18002 22482
rect 19742 22430 19794 22482
rect 20190 22430 20242 22482
rect 23438 22430 23490 22482
rect 24334 22430 24386 22482
rect 25454 22430 25506 22482
rect 27582 22430 27634 22482
rect 4286 22318 4338 22370
rect 15262 22318 15314 22370
rect 17726 22318 17778 22370
rect 18510 22318 18562 22370
rect 19182 22318 19234 22370
rect 20302 22318 20354 22370
rect 21758 22318 21810 22370
rect 24670 22318 24722 22370
rect 15822 22206 15874 22258
rect 18622 22206 18674 22258
rect 22766 22206 22818 22258
rect 15598 22094 15650 22146
rect 17390 22094 17442 22146
rect 19294 22094 19346 22146
rect 21870 22094 21922 22146
rect 23326 22094 23378 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 13918 21758 13970 21810
rect 18062 21758 18114 21810
rect 18174 21758 18226 21810
rect 19630 21758 19682 21810
rect 22094 21758 22146 21810
rect 13358 21646 13410 21698
rect 13470 21646 13522 21698
rect 17838 21646 17890 21698
rect 17950 21646 18002 21698
rect 18958 21646 19010 21698
rect 19182 21646 19234 21698
rect 21646 21646 21698 21698
rect 21758 21646 21810 21698
rect 21870 21646 21922 21698
rect 22318 21646 22370 21698
rect 22990 21646 23042 21698
rect 23214 21646 23266 21698
rect 12910 21534 12962 21586
rect 13134 21534 13186 21586
rect 17502 21534 17554 21586
rect 18622 21534 18674 21586
rect 20526 21534 20578 21586
rect 22542 21534 22594 21586
rect 23998 21534 24050 21586
rect 37326 21534 37378 21586
rect 37774 21534 37826 21586
rect 9998 21422 10050 21474
rect 12126 21422 12178 21474
rect 20974 21422 21026 21474
rect 21758 21422 21810 21474
rect 39902 21422 39954 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 18062 20974 18114 21026
rect 18398 20974 18450 21026
rect 16158 20862 16210 20914
rect 20078 20862 20130 20914
rect 22542 20862 22594 20914
rect 40014 20862 40066 20914
rect 12238 20750 12290 20802
rect 12574 20750 12626 20802
rect 15598 20750 15650 20802
rect 16830 20750 16882 20802
rect 17278 20750 17330 20802
rect 18734 20750 18786 20802
rect 20526 20750 20578 20802
rect 22430 20750 22482 20802
rect 22878 20750 22930 20802
rect 26350 20750 26402 20802
rect 27246 20750 27298 20802
rect 27358 20750 27410 20802
rect 37662 20750 37714 20802
rect 12462 20638 12514 20690
rect 15934 20638 15986 20690
rect 17390 20638 17442 20690
rect 18958 20638 19010 20690
rect 21870 20638 21922 20690
rect 25902 20638 25954 20690
rect 26798 20638 26850 20690
rect 27694 20638 27746 20690
rect 18174 20526 18226 20578
rect 19294 20526 19346 20578
rect 21534 20526 21586 20578
rect 22990 20526 23042 20578
rect 25230 20526 25282 20578
rect 25678 20526 25730 20578
rect 25790 20526 25842 20578
rect 26574 20526 26626 20578
rect 26686 20526 26738 20578
rect 27582 20526 27634 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 16270 20190 16322 20242
rect 13022 20078 13074 20130
rect 15710 20078 15762 20130
rect 15822 20078 15874 20130
rect 16606 20078 16658 20130
rect 26238 20078 26290 20130
rect 28702 20078 28754 20130
rect 28814 20078 28866 20130
rect 12238 19966 12290 20018
rect 17726 19966 17778 20018
rect 18286 19966 18338 20018
rect 18734 19966 18786 20018
rect 19070 19966 19122 20018
rect 25454 19966 25506 20018
rect 37662 19966 37714 20018
rect 15150 19854 15202 19906
rect 23102 19854 23154 19906
rect 28366 19854 28418 19906
rect 15822 19742 15874 19794
rect 28814 19742 28866 19794
rect 40014 19742 40066 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 15822 19406 15874 19458
rect 19854 19294 19906 19346
rect 21422 19294 21474 19346
rect 26126 19294 26178 19346
rect 28254 19294 28306 19346
rect 15934 19182 15986 19234
rect 16606 19182 16658 19234
rect 17726 19182 17778 19234
rect 19742 19182 19794 19234
rect 20078 19182 20130 19234
rect 24222 19182 24274 19234
rect 25454 19182 25506 19234
rect 18062 19070 18114 19122
rect 18846 19070 18898 19122
rect 23550 19070 23602 19122
rect 15374 18958 15426 19010
rect 16830 18958 16882 19010
rect 17166 18958 17218 19010
rect 18174 18958 18226 19010
rect 19630 18958 19682 19010
rect 25006 18958 25058 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 15486 18622 15538 18674
rect 23662 18622 23714 18674
rect 18398 18510 18450 18562
rect 19742 18510 19794 18562
rect 20974 18510 21026 18562
rect 12238 18398 12290 18450
rect 16494 18398 16546 18450
rect 16718 18398 16770 18450
rect 17950 18398 18002 18450
rect 19406 18398 19458 18450
rect 21870 18398 21922 18450
rect 22430 18398 22482 18450
rect 22654 18398 22706 18450
rect 22766 18398 22818 18450
rect 23886 18398 23938 18450
rect 12910 18286 12962 18338
rect 15038 18286 15090 18338
rect 15822 18286 15874 18338
rect 23214 18174 23266 18226
rect 23550 18174 23602 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 22094 17838 22146 17890
rect 18174 17726 18226 17778
rect 20638 17726 20690 17778
rect 21534 17726 21586 17778
rect 21870 17726 21922 17778
rect 26014 17726 26066 17778
rect 40014 17726 40066 17778
rect 13806 17614 13858 17666
rect 17726 17614 17778 17666
rect 18622 17614 18674 17666
rect 18958 17614 19010 17666
rect 19742 17614 19794 17666
rect 21646 17614 21698 17666
rect 22318 17614 22370 17666
rect 22542 17614 22594 17666
rect 26126 17614 26178 17666
rect 37662 17614 37714 17666
rect 13470 17502 13522 17554
rect 17950 17502 18002 17554
rect 18286 17502 18338 17554
rect 19182 17502 19234 17554
rect 22990 17502 23042 17554
rect 23214 17502 23266 17554
rect 18846 17390 18898 17442
rect 19406 17390 19458 17442
rect 19630 17390 19682 17442
rect 20750 17390 20802 17442
rect 21422 17390 21474 17442
rect 22878 17390 22930 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 18510 17054 18562 17106
rect 18734 17054 18786 17106
rect 14702 16942 14754 16994
rect 14030 16830 14082 16882
rect 17502 16830 17554 16882
rect 19070 16830 19122 16882
rect 23102 16830 23154 16882
rect 16830 16718 16882 16770
rect 19518 16718 19570 16770
rect 18846 16606 18898 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 17838 16158 17890 16210
rect 24782 16158 24834 16210
rect 26910 16158 26962 16210
rect 17950 16046 18002 16098
rect 18286 16046 18338 16098
rect 18958 16046 19010 16098
rect 20750 16046 20802 16098
rect 21646 16046 21698 16098
rect 22766 16046 22818 16098
rect 23998 16046 24050 16098
rect 22990 15934 23042 15986
rect 17726 15822 17778 15874
rect 19182 15822 19234 15874
rect 20414 15822 20466 15874
rect 21870 15822 21922 15874
rect 21982 15822 22034 15874
rect 22094 15822 22146 15874
rect 22206 15822 22258 15874
rect 23662 15822 23714 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 19518 15486 19570 15538
rect 21758 15486 21810 15538
rect 18174 15374 18226 15426
rect 18510 15374 18562 15426
rect 18846 15374 18898 15426
rect 21422 15374 21474 15426
rect 22542 15374 22594 15426
rect 22766 15374 22818 15426
rect 25230 15374 25282 15426
rect 25566 15374 25618 15426
rect 17614 15262 17666 15314
rect 17726 15262 17778 15314
rect 17838 15262 17890 15314
rect 19070 15262 19122 15314
rect 22430 15262 22482 15314
rect 18622 15150 18674 15202
rect 19182 15038 19234 15090
rect 19630 15038 19682 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 16718 14590 16770 14642
rect 18846 14590 18898 14642
rect 21534 14590 21586 14642
rect 23550 14590 23602 14642
rect 25678 14590 25730 14642
rect 16046 14478 16098 14530
rect 19294 14478 19346 14530
rect 19518 14478 19570 14530
rect 19854 14478 19906 14530
rect 20414 14478 20466 14530
rect 21870 14478 21922 14530
rect 22318 14478 22370 14530
rect 22766 14478 22818 14530
rect 22206 14366 22258 14418
rect 19630 14254 19682 14306
rect 19742 14254 19794 14306
rect 20638 14254 20690 14306
rect 22094 14254 22146 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 17502 13918 17554 13970
rect 18958 13918 19010 13970
rect 19070 13918 19122 13970
rect 24558 13918 24610 13970
rect 14702 13806 14754 13858
rect 18734 13806 18786 13858
rect 19742 13806 19794 13858
rect 14030 13694 14082 13746
rect 19182 13694 19234 13746
rect 19406 13694 19458 13746
rect 20078 13694 20130 13746
rect 20302 13694 20354 13746
rect 21198 13694 21250 13746
rect 16830 13582 16882 13634
rect 20190 13582 20242 13634
rect 21982 13582 22034 13634
rect 24110 13582 24162 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 18510 13022 18562 13074
rect 20638 13022 20690 13074
rect 21758 13022 21810 13074
rect 17726 12910 17778 12962
rect 21534 12910 21586 12962
rect 21870 12910 21922 12962
rect 22094 12910 22146 12962
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 20974 12350 21026 12402
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 18734 5182 18786 5234
rect 24782 5182 24834 5234
rect 17838 5070 17890 5122
rect 23774 5070 23826 5122
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 17502 4286 17554 4338
rect 20414 4286 20466 4338
rect 25790 4286 25842 4338
rect 18510 4062 18562 4114
rect 21422 4062 21474 4114
rect 26798 4062 26850 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18846 3614 18898 3666
rect 22094 3614 22146 3666
rect 25566 3614 25618 3666
rect 19742 3502 19794 3554
rect 21086 3502 21138 3554
rect 25006 3502 25058 3554
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 16800 41200 16912 42000
rect 17472 41200 17584 42000
rect 18144 41200 18256 42000
rect 22848 41200 22960 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 16828 37492 16884 41200
rect 17276 38610 17332 38622
rect 17276 38558 17278 38610
rect 17330 38558 17332 38610
rect 17276 37938 17332 38558
rect 17500 38276 17556 41200
rect 18172 38610 18228 41200
rect 18172 38558 18174 38610
rect 18226 38558 18228 38610
rect 18172 38546 18228 38558
rect 17500 38210 17556 38220
rect 18620 38276 18676 38286
rect 18620 38182 18676 38220
rect 22876 38276 22932 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 22876 38210 22932 38220
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 17276 37886 17278 37938
rect 17330 37886 17332 37938
rect 17276 37874 17332 37886
rect 17836 38050 17892 38062
rect 17836 37998 17838 38050
rect 17890 37998 17892 38050
rect 16828 37426 16884 37436
rect 17388 37268 17444 37278
rect 17052 37266 17444 37268
rect 17052 37214 17390 37266
rect 17442 37214 17444 37266
rect 17052 37212 17444 37214
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4172 27636 4228 27646
rect 1932 27186 1988 27198
rect 1932 27134 1934 27186
rect 1986 27134 1988 27186
rect 1932 26292 1988 27134
rect 1932 26226 1988 26236
rect 1932 26066 1988 26078
rect 1932 26014 1934 26066
rect 1986 26014 1988 26066
rect 1932 25620 1988 26014
rect 1932 25554 1988 25564
rect 2044 25618 2100 25630
rect 2044 25566 2046 25618
rect 2098 25566 2100 25618
rect 2044 24948 2100 25566
rect 2044 24882 2100 24892
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 1932 23538 1988 23548
rect 1932 22932 1988 22942
rect 1932 22838 1988 22876
rect 1932 22482 1988 22494
rect 1932 22430 1934 22482
rect 1986 22430 1988 22482
rect 1932 21588 1988 22430
rect 1932 21522 1988 21532
rect 4172 20020 4228 27580
rect 15148 27636 15204 27646
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 15148 27186 15204 27580
rect 15148 27134 15150 27186
rect 15202 27134 15204 27186
rect 15148 27122 15204 27134
rect 4284 27076 4340 27086
rect 4284 26982 4340 27020
rect 12124 27076 12180 27086
rect 12124 26962 12180 27020
rect 12124 26910 12126 26962
rect 12178 26910 12180 26962
rect 12124 26898 12180 26910
rect 14364 27074 14420 27086
rect 14364 27022 14366 27074
rect 14418 27022 14420 27074
rect 12460 26850 12516 26862
rect 12460 26798 12462 26850
rect 12514 26798 12516 26850
rect 4284 26292 4340 26302
rect 4284 26198 4340 26236
rect 12124 26292 12180 26302
rect 10220 26178 10276 26190
rect 10220 26126 10222 26178
rect 10274 26126 10276 26178
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4284 25508 4340 25518
rect 4284 25414 4340 25452
rect 10220 25508 10276 26126
rect 11676 25732 11732 25742
rect 11676 25638 11732 25676
rect 10220 25442 10276 25452
rect 11676 25396 11732 25406
rect 11676 25302 11732 25340
rect 11788 25396 11844 25406
rect 11788 25394 12068 25396
rect 11788 25342 11790 25394
rect 11842 25342 12068 25394
rect 11788 25340 12068 25342
rect 11788 25330 11844 25340
rect 12012 25060 12068 25340
rect 12124 25394 12180 26236
rect 12348 26178 12404 26190
rect 12348 26126 12350 26178
rect 12402 26126 12404 26178
rect 12348 25732 12404 26126
rect 12348 25666 12404 25676
rect 12348 25508 12404 25518
rect 12460 25508 12516 26798
rect 13132 26292 13188 26302
rect 13132 26198 13188 26236
rect 13804 26292 13860 26302
rect 12404 25452 12628 25508
rect 12348 25414 12404 25452
rect 12124 25342 12126 25394
rect 12178 25342 12180 25394
rect 12124 25330 12180 25342
rect 12012 25004 12404 25060
rect 12348 24946 12404 25004
rect 12348 24894 12350 24946
rect 12402 24894 12404 24946
rect 12348 24882 12404 24894
rect 12572 24946 12628 25452
rect 13580 25284 13636 25294
rect 13804 25284 13860 26236
rect 13580 25282 13860 25284
rect 13580 25230 13582 25282
rect 13634 25230 13860 25282
rect 13580 25228 13860 25230
rect 13580 25218 13636 25228
rect 12572 24894 12574 24946
rect 12626 24894 12628 24946
rect 12572 24882 12628 24894
rect 13804 25172 13860 25228
rect 14364 25172 14420 27022
rect 16828 26964 16884 26974
rect 16156 26292 16212 26302
rect 14476 26180 14532 26190
rect 14476 26086 14532 26124
rect 16044 26180 16100 26190
rect 16044 25618 16100 26124
rect 16044 25566 16046 25618
rect 16098 25566 16100 25618
rect 16044 25554 16100 25566
rect 16156 25506 16212 26236
rect 16604 26180 16660 26190
rect 16604 26086 16660 26124
rect 16156 25454 16158 25506
rect 16210 25454 16212 25506
rect 16156 25442 16212 25454
rect 16604 25620 16660 25630
rect 16604 25506 16660 25564
rect 16604 25454 16606 25506
rect 16658 25454 16660 25506
rect 16604 25442 16660 25454
rect 15932 25284 15988 25294
rect 14476 25172 14532 25182
rect 14364 25116 14476 25172
rect 12684 24722 12740 24734
rect 12684 24670 12686 24722
rect 12738 24670 12740 24722
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4284 23938 4340 23950
rect 4284 23886 4286 23938
rect 4338 23886 4340 23938
rect 4284 23828 4340 23886
rect 4284 23762 4340 23772
rect 12684 23604 12740 24670
rect 13468 24050 13524 24062
rect 13468 23998 13470 24050
rect 13522 23998 13524 24050
rect 13468 23828 13524 23998
rect 13468 23762 13524 23772
rect 12684 23538 12740 23548
rect 13468 23492 13524 23502
rect 11004 23268 11060 23278
rect 4284 23156 4340 23166
rect 4284 23062 4340 23100
rect 11004 23042 11060 23212
rect 11004 22990 11006 23042
rect 11058 22990 11060 23042
rect 11004 22978 11060 22990
rect 13132 23042 13188 23054
rect 13132 22990 13134 23042
rect 13186 22990 13188 23042
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 13132 22596 13188 22990
rect 13132 22530 13188 22540
rect 4284 22370 4340 22382
rect 4284 22318 4286 22370
rect 4338 22318 4340 22370
rect 4284 21476 4340 22318
rect 12908 21812 12964 21822
rect 4284 21410 4340 21420
rect 9996 21700 10052 21710
rect 9996 21474 10052 21644
rect 12908 21586 12964 21756
rect 13356 21700 13412 21710
rect 13356 21606 13412 21644
rect 13468 21698 13524 23436
rect 13804 23156 13860 25116
rect 14476 25106 14532 25116
rect 15596 23828 15652 23838
rect 14924 23826 15652 23828
rect 14924 23774 15598 23826
rect 15650 23774 15652 23826
rect 14924 23772 15652 23774
rect 14252 23492 14308 23502
rect 14252 23266 14308 23436
rect 14924 23378 14980 23772
rect 15596 23762 15652 23772
rect 15484 23604 15540 23614
rect 14924 23326 14926 23378
rect 14978 23326 14980 23378
rect 14924 23314 14980 23326
rect 15372 23380 15428 23390
rect 15372 23286 15428 23324
rect 15484 23378 15540 23548
rect 15484 23326 15486 23378
rect 15538 23326 15540 23378
rect 15484 23314 15540 23326
rect 14252 23214 14254 23266
rect 14306 23214 14308 23266
rect 14252 23202 14308 23214
rect 14364 23268 14420 23278
rect 14364 23174 14420 23212
rect 13804 23154 14196 23156
rect 13804 23102 13806 23154
rect 13858 23102 14196 23154
rect 13804 23100 14196 23102
rect 13804 23090 13860 23100
rect 13916 21812 13972 23100
rect 14140 22482 14196 23100
rect 15708 23154 15764 23166
rect 15708 23102 15710 23154
rect 15762 23102 15764 23154
rect 14812 23044 14868 23054
rect 14812 22950 14868 22988
rect 15596 23044 15652 23054
rect 15596 22950 15652 22988
rect 14364 22932 14420 22942
rect 14364 22838 14420 22876
rect 15260 22932 15316 22942
rect 14140 22430 14142 22482
rect 14194 22430 14196 22482
rect 14140 22418 14196 22430
rect 15260 22370 15316 22876
rect 15484 22596 15540 22606
rect 15484 22502 15540 22540
rect 15260 22318 15262 22370
rect 15314 22318 15316 22370
rect 15260 22306 15316 22318
rect 13916 21718 13972 21756
rect 15596 22146 15652 22158
rect 15596 22094 15598 22146
rect 15650 22094 15652 22146
rect 15596 21812 15652 22094
rect 15596 21746 15652 21756
rect 15708 22148 15764 23102
rect 15932 23156 15988 25228
rect 16268 25172 16324 25182
rect 16268 23940 16324 25116
rect 16828 25172 16884 26908
rect 17052 26180 17108 37212
rect 17388 37202 17444 37212
rect 17388 27860 17444 27870
rect 17836 27860 17892 37998
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 18396 37492 18452 37502
rect 18396 37398 18452 37436
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 17164 27858 17444 27860
rect 17164 27806 17390 27858
rect 17442 27806 17444 27858
rect 17164 27804 17444 27806
rect 17164 26852 17220 27804
rect 17388 27794 17444 27804
rect 17500 27804 17892 27860
rect 17388 27636 17444 27646
rect 17388 27542 17444 27580
rect 17500 27412 17556 27804
rect 17276 27356 17556 27412
rect 17724 27634 17780 27646
rect 17724 27582 17726 27634
rect 17778 27582 17780 27634
rect 17276 27186 17332 27356
rect 17276 27134 17278 27186
rect 17330 27134 17332 27186
rect 17276 27122 17332 27134
rect 17612 27074 17668 27086
rect 17612 27022 17614 27074
rect 17666 27022 17668 27074
rect 17612 26964 17668 27022
rect 17612 26898 17668 26908
rect 17164 26786 17220 26796
rect 17500 26852 17556 26862
rect 16940 25620 16996 25630
rect 16940 25526 16996 25564
rect 17052 25506 17108 26124
rect 17052 25454 17054 25506
rect 17106 25454 17108 25506
rect 17052 25442 17108 25454
rect 17388 26290 17444 26302
rect 17388 26238 17390 26290
rect 17442 26238 17444 26290
rect 17276 25396 17332 25406
rect 17276 25302 17332 25340
rect 16828 24946 16884 25116
rect 16828 24894 16830 24946
rect 16882 24894 16884 24946
rect 16828 24882 16884 24894
rect 16940 25282 16996 25294
rect 16940 25230 16942 25282
rect 16994 25230 16996 25282
rect 16268 23846 16324 23884
rect 16940 23938 16996 25230
rect 17388 25284 17444 26238
rect 17500 25508 17556 26796
rect 17724 26514 17780 27582
rect 17724 26462 17726 26514
rect 17778 26462 17780 26514
rect 17724 26450 17780 26462
rect 17836 26514 17892 27804
rect 20636 27858 20692 27870
rect 20636 27806 20638 27858
rect 20690 27806 20692 27858
rect 18284 27748 18340 27758
rect 18284 26964 18340 27692
rect 20412 27748 20468 27758
rect 20636 27748 20692 27806
rect 20468 27692 20804 27748
rect 20412 27654 20468 27692
rect 20524 27188 20580 27198
rect 20524 27186 20692 27188
rect 20524 27134 20526 27186
rect 20578 27134 20692 27186
rect 20524 27132 20692 27134
rect 20524 27122 20580 27132
rect 20412 27076 20468 27086
rect 18284 26898 18340 26908
rect 18396 26962 18452 26974
rect 18396 26910 18398 26962
rect 18450 26910 18452 26962
rect 18396 26908 18452 26910
rect 20412 26908 20468 27020
rect 18396 26852 18900 26908
rect 20412 26852 20580 26908
rect 17836 26462 17838 26514
rect 17890 26462 17892 26514
rect 17836 26450 17892 26462
rect 18732 26516 18788 26526
rect 18732 26422 18788 26460
rect 18844 26514 18900 26852
rect 20524 26786 20580 26796
rect 20636 26740 20692 27132
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20636 26674 20692 26684
rect 20748 26908 20804 27692
rect 21420 27746 21476 27758
rect 22764 27748 22820 27758
rect 21420 27694 21422 27746
rect 21474 27694 21476 27746
rect 21420 27186 21476 27694
rect 22652 27692 22764 27748
rect 21868 27300 21924 27310
rect 21868 27298 22596 27300
rect 21868 27246 21870 27298
rect 21922 27246 22596 27298
rect 21868 27244 22596 27246
rect 21868 27234 21924 27244
rect 21420 27134 21422 27186
rect 21474 27134 21476 27186
rect 21420 27122 21476 27134
rect 21532 27132 21812 27188
rect 21532 27076 21588 27132
rect 21532 26982 21588 27020
rect 21308 26962 21364 26974
rect 21308 26910 21310 26962
rect 21362 26910 21364 26962
rect 20748 26852 21140 26908
rect 19836 26618 20100 26628
rect 18844 26462 18846 26514
rect 18898 26462 18900 26514
rect 18844 26450 18900 26462
rect 19628 26516 19684 26526
rect 19628 26422 19684 26460
rect 20636 26516 20692 26526
rect 20748 26516 20804 26852
rect 20636 26514 20804 26516
rect 20636 26462 20638 26514
rect 20690 26462 20804 26514
rect 20636 26460 20804 26462
rect 20636 26450 20692 26460
rect 17500 25414 17556 25452
rect 17612 26290 17668 26302
rect 17612 26238 17614 26290
rect 17666 26238 17668 26290
rect 17388 25218 17444 25228
rect 17612 24164 17668 26238
rect 18060 26290 18116 26302
rect 18060 26238 18062 26290
rect 18114 26238 18116 26290
rect 18060 25172 18116 26238
rect 18396 26290 18452 26302
rect 18396 26238 18398 26290
rect 18450 26238 18452 26290
rect 18396 25730 18452 26238
rect 18396 25678 18398 25730
rect 18450 25678 18452 25730
rect 18396 25666 18452 25678
rect 18956 26292 19012 26302
rect 18284 25508 18340 25518
rect 18844 25508 18900 25518
rect 18284 25506 18564 25508
rect 18284 25454 18286 25506
rect 18338 25454 18564 25506
rect 18284 25452 18564 25454
rect 18284 25396 18340 25452
rect 18284 25330 18340 25340
rect 18396 25282 18452 25294
rect 18396 25230 18398 25282
rect 18450 25230 18452 25282
rect 18396 25172 18452 25230
rect 18060 25116 18452 25172
rect 18396 24836 18452 25116
rect 17612 24098 17668 24108
rect 18172 24164 18228 24174
rect 16940 23886 16942 23938
rect 16994 23886 16996 23938
rect 16716 23714 16772 23726
rect 16716 23662 16718 23714
rect 16770 23662 16772 23714
rect 16716 23380 16772 23662
rect 16940 23604 16996 23886
rect 17500 23940 17556 23950
rect 17500 23846 17556 23884
rect 16940 23538 16996 23548
rect 17612 23716 17668 23726
rect 16716 23314 16772 23324
rect 15932 23154 16100 23156
rect 15932 23102 15934 23154
rect 15986 23102 16100 23154
rect 15932 23100 16100 23102
rect 15932 23090 15988 23100
rect 15820 22260 15876 22270
rect 15820 22166 15876 22204
rect 13468 21646 13470 21698
rect 13522 21646 13524 21698
rect 13468 21634 13524 21646
rect 13132 21588 13188 21598
rect 12908 21534 12910 21586
rect 12962 21534 12964 21586
rect 12908 21522 12964 21534
rect 13020 21586 13188 21588
rect 13020 21534 13134 21586
rect 13186 21534 13188 21586
rect 13020 21532 13188 21534
rect 9996 21422 9998 21474
rect 10050 21422 10052 21474
rect 9996 21410 10052 21422
rect 12124 21476 12180 21486
rect 12124 21474 12292 21476
rect 12124 21422 12126 21474
rect 12178 21422 12292 21474
rect 12124 21420 12292 21422
rect 12124 21410 12180 21420
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 12236 20802 12292 21420
rect 12236 20750 12238 20802
rect 12290 20750 12292 20802
rect 12236 20738 12292 20750
rect 12460 21252 12516 21262
rect 12460 20690 12516 21196
rect 13020 21028 13076 21532
rect 13132 21522 13188 21532
rect 12572 20972 13076 21028
rect 12572 20802 12628 20972
rect 12572 20750 12574 20802
rect 12626 20750 12628 20802
rect 12572 20738 12628 20750
rect 15148 20804 15204 20814
rect 12460 20638 12462 20690
rect 12514 20638 12516 20690
rect 12460 20626 12516 20638
rect 13020 20132 13076 20142
rect 13020 20038 13076 20076
rect 4172 19954 4228 19964
rect 12236 20018 12292 20030
rect 12236 19966 12238 20018
rect 12290 19966 12292 20018
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 12236 19012 12292 19966
rect 15148 19906 15204 20748
rect 15596 20802 15652 20814
rect 15596 20750 15598 20802
rect 15650 20750 15652 20802
rect 15148 19854 15150 19906
rect 15202 19854 15204 19906
rect 15148 19842 15204 19854
rect 15484 20132 15540 20142
rect 15484 19460 15540 20076
rect 15484 19394 15540 19404
rect 12236 18450 12292 18956
rect 12236 18398 12238 18450
rect 12290 18398 12292 18450
rect 12236 18386 12292 18398
rect 14028 19012 14084 19022
rect 12908 18340 12964 18350
rect 13804 18340 13860 18350
rect 12908 18338 13524 18340
rect 12908 18286 12910 18338
rect 12962 18286 13524 18338
rect 12908 18284 13524 18286
rect 12908 18274 12964 18284
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 13468 17554 13524 18284
rect 13804 17666 13860 18284
rect 13804 17614 13806 17666
rect 13858 17614 13860 17666
rect 13804 17602 13860 17614
rect 13468 17502 13470 17554
rect 13522 17502 13524 17554
rect 13468 17490 13524 17502
rect 14028 16884 14084 18956
rect 15372 19012 15428 19022
rect 15428 18956 15540 19012
rect 15372 18918 15428 18956
rect 15036 18900 15092 18910
rect 15036 18338 15092 18844
rect 15484 18674 15540 18956
rect 15596 18900 15652 20750
rect 15708 20130 15764 22092
rect 15932 20804 15988 20814
rect 15932 20690 15988 20748
rect 15932 20638 15934 20690
rect 15986 20638 15988 20690
rect 15932 20626 15988 20638
rect 16044 20356 16100 23100
rect 16156 22372 16212 22382
rect 16156 20914 16212 22316
rect 17388 22146 17444 22158
rect 17388 22094 17390 22146
rect 17442 22094 17444 22146
rect 17388 21252 17444 22094
rect 17388 21186 17444 21196
rect 17500 21700 17556 21710
rect 17500 21586 17556 21644
rect 17500 21534 17502 21586
rect 17554 21534 17556 21586
rect 16156 20862 16158 20914
rect 16210 20862 16212 20914
rect 16156 20850 16212 20862
rect 16268 20804 16324 20814
rect 16156 20356 16212 20366
rect 16044 20300 16156 20356
rect 16156 20290 16212 20300
rect 16268 20242 16324 20748
rect 16828 20804 16884 20814
rect 16828 20710 16884 20748
rect 17276 20802 17332 20814
rect 17276 20750 17278 20802
rect 17330 20750 17332 20802
rect 16268 20190 16270 20242
rect 16322 20190 16324 20242
rect 16268 20178 16324 20190
rect 16940 20244 16996 20254
rect 15708 20078 15710 20130
rect 15762 20078 15764 20130
rect 15708 20066 15764 20078
rect 15820 20132 15876 20142
rect 15820 20038 15876 20076
rect 16604 20130 16660 20142
rect 16604 20078 16606 20130
rect 16658 20078 16660 20130
rect 16604 19908 16660 20078
rect 15820 19796 15876 19806
rect 15708 19794 15876 19796
rect 15708 19742 15822 19794
rect 15874 19742 15876 19794
rect 15708 19740 15876 19742
rect 15708 19124 15764 19740
rect 15820 19730 15876 19740
rect 15820 19460 15876 19470
rect 15820 19366 15876 19404
rect 15932 19236 15988 19246
rect 15932 19142 15988 19180
rect 16604 19236 16660 19852
rect 16604 19142 16660 19180
rect 15708 19068 15876 19124
rect 15708 18900 15764 18910
rect 15596 18844 15708 18900
rect 15708 18834 15764 18844
rect 15484 18622 15486 18674
rect 15538 18622 15540 18674
rect 15484 18610 15540 18622
rect 15820 18564 15876 19068
rect 16828 19012 16884 19022
rect 16492 18956 16828 19012
rect 15820 18508 15988 18564
rect 15932 18452 15988 18508
rect 15932 18386 15988 18396
rect 16492 18450 16548 18956
rect 16828 18918 16884 18956
rect 16940 18788 16996 20188
rect 17276 20132 17332 20750
rect 17388 20690 17444 20702
rect 17388 20638 17390 20690
rect 17442 20638 17444 20690
rect 17388 20356 17444 20638
rect 17388 20290 17444 20300
rect 17500 20244 17556 21534
rect 17500 20178 17556 20188
rect 17276 20066 17332 20076
rect 17164 19010 17220 19022
rect 17164 18958 17166 19010
rect 17218 18958 17220 19010
rect 17164 18900 17220 18958
rect 17164 18834 17220 18844
rect 16492 18398 16494 18450
rect 16546 18398 16548 18450
rect 16492 18386 16548 18398
rect 16716 18732 16996 18788
rect 16716 18450 16772 18732
rect 16716 18398 16718 18450
rect 16770 18398 16772 18450
rect 16716 18386 16772 18398
rect 15036 18286 15038 18338
rect 15090 18286 15092 18338
rect 15036 18274 15092 18286
rect 15820 18340 15876 18350
rect 15820 18246 15876 18284
rect 17612 18228 17668 23660
rect 17948 22484 18004 22494
rect 17948 22390 18004 22428
rect 17724 22370 17780 22382
rect 17724 22318 17726 22370
rect 17778 22318 17780 22370
rect 17724 22260 17780 22318
rect 17724 22194 17780 22204
rect 18060 21812 18116 21822
rect 18060 21718 18116 21756
rect 18172 21810 18228 24108
rect 18396 23716 18452 24780
rect 18396 23650 18452 23660
rect 18508 22372 18564 25452
rect 18844 25394 18900 25452
rect 18844 25342 18846 25394
rect 18898 25342 18900 25394
rect 18844 25330 18900 25342
rect 18956 24948 19012 26236
rect 19292 26290 19348 26302
rect 19292 26238 19294 26290
rect 19346 26238 19348 26290
rect 19292 25396 19348 26238
rect 21084 26292 21140 26852
rect 21308 26516 21364 26910
rect 21308 26450 21364 26460
rect 21644 26964 21700 26974
rect 21532 26292 21588 26302
rect 21644 26292 21700 26908
rect 21756 26908 21812 27132
rect 22540 27186 22596 27244
rect 22540 27134 22542 27186
rect 22594 27134 22596 27186
rect 22540 27122 22596 27134
rect 22092 27076 22148 27086
rect 22092 26982 22148 27020
rect 22428 26962 22484 26974
rect 22428 26910 22430 26962
rect 22482 26910 22484 26962
rect 22428 26908 22484 26910
rect 21756 26852 22484 26908
rect 22652 26962 22708 27692
rect 22764 27682 22820 27692
rect 23548 27748 23604 27758
rect 23548 27654 23604 27692
rect 24556 27748 24612 37998
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 24556 27682 24612 27692
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 26908 27188 26964 27198
rect 22652 26910 22654 26962
rect 22706 26910 22708 26962
rect 22652 26898 22708 26910
rect 22764 27076 22820 27086
rect 21084 26290 21700 26292
rect 21084 26238 21086 26290
rect 21138 26238 21534 26290
rect 21586 26238 21700 26290
rect 21084 26236 21700 26238
rect 22540 26516 22596 26526
rect 21084 26226 21140 26236
rect 21532 26226 21588 26236
rect 22204 26180 22260 26190
rect 21756 26178 22260 26180
rect 21756 26126 22206 26178
rect 22258 26126 22260 26178
rect 21756 26124 22260 26126
rect 21756 25730 21812 26124
rect 22204 26114 22260 26124
rect 21756 25678 21758 25730
rect 21810 25678 21812 25730
rect 21756 25666 21812 25678
rect 21532 25620 21588 25630
rect 21588 25564 21700 25620
rect 21532 25554 21588 25564
rect 21644 25396 21700 25564
rect 22428 25508 22484 25546
rect 22540 25508 22596 26460
rect 22484 25452 22596 25508
rect 22428 25442 22484 25452
rect 21756 25396 21812 25406
rect 21644 25394 21812 25396
rect 21644 25342 21758 25394
rect 21810 25342 21812 25394
rect 21644 25340 21812 25342
rect 19292 25330 19348 25340
rect 18956 24882 19012 24892
rect 19180 25282 19236 25294
rect 19180 25230 19182 25282
rect 19234 25230 19236 25282
rect 19068 24164 19124 24174
rect 19068 24050 19124 24108
rect 19068 23998 19070 24050
rect 19122 23998 19124 24050
rect 19068 23986 19124 23998
rect 18732 23940 18788 23950
rect 18508 22278 18564 22316
rect 18620 23828 18676 23838
rect 18620 22484 18676 23772
rect 18732 23716 18788 23884
rect 19180 23828 19236 25230
rect 21756 25284 21812 25340
rect 21868 25396 21924 25406
rect 22092 25396 22148 25406
rect 21868 25394 22148 25396
rect 21868 25342 21870 25394
rect 21922 25342 22094 25394
rect 22146 25342 22148 25394
rect 21868 25340 22148 25342
rect 21868 25330 21924 25340
rect 22092 25330 22148 25340
rect 22316 25284 22372 25294
rect 21756 25218 21812 25228
rect 22204 25282 22372 25284
rect 22204 25230 22318 25282
rect 22370 25230 22372 25282
rect 22204 25228 22372 25230
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19852 24836 19908 24846
rect 19852 24742 19908 24780
rect 20636 24836 20692 24846
rect 20636 24742 20692 24780
rect 21868 24836 21924 24846
rect 21868 24742 21924 24780
rect 19740 24724 19796 24734
rect 19628 23940 19684 23950
rect 19628 23846 19684 23884
rect 19180 23762 19236 23772
rect 19740 23716 19796 24668
rect 20076 24722 20132 24734
rect 20076 24670 20078 24722
rect 20130 24670 20132 24722
rect 19852 24052 19908 24062
rect 19852 23938 19908 23996
rect 19852 23886 19854 23938
rect 19906 23886 19908 23938
rect 19852 23874 19908 23886
rect 20076 23940 20132 24670
rect 22204 24722 22260 25228
rect 22316 25218 22372 25228
rect 22764 25172 22820 27020
rect 24668 27074 24724 27086
rect 24668 27022 24670 27074
rect 24722 27022 24724 27074
rect 24220 26964 24276 27002
rect 24220 26898 24276 26908
rect 24668 26964 24724 27022
rect 24668 26898 24724 26908
rect 25340 26962 25396 26974
rect 25340 26910 25342 26962
rect 25394 26910 25396 26962
rect 22428 25116 22820 25172
rect 22876 26740 22932 26750
rect 22204 24670 22206 24722
rect 22258 24670 22260 24722
rect 21420 24610 21476 24622
rect 21420 24558 21422 24610
rect 21474 24558 21476 24610
rect 20076 23874 20132 23884
rect 20524 24498 20580 24510
rect 20524 24446 20526 24498
rect 20578 24446 20580 24498
rect 20524 24052 20580 24446
rect 20524 23938 20580 23996
rect 20524 23886 20526 23938
rect 20578 23886 20580 23938
rect 20524 23874 20580 23886
rect 18732 23266 18788 23660
rect 18732 23214 18734 23266
rect 18786 23214 18788 23266
rect 18732 23202 18788 23214
rect 19628 23660 19796 23716
rect 20188 23828 20244 23838
rect 19628 23604 19684 23660
rect 19628 22596 19684 23548
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19628 22540 19796 22596
rect 18620 22258 18676 22428
rect 19740 22482 19796 22540
rect 19740 22430 19742 22482
rect 19794 22430 19796 22482
rect 19740 22418 19796 22430
rect 20188 22482 20244 23772
rect 20188 22430 20190 22482
rect 20242 22430 20244 22482
rect 20188 22418 20244 22430
rect 18620 22206 18622 22258
rect 18674 22206 18676 22258
rect 18620 22194 18676 22206
rect 19180 22370 19236 22382
rect 19180 22318 19182 22370
rect 19234 22318 19236 22370
rect 19180 21924 19236 22318
rect 19628 22372 19684 22382
rect 19292 22148 19348 22158
rect 19292 22146 19460 22148
rect 19292 22094 19294 22146
rect 19346 22094 19460 22146
rect 19292 22092 19460 22094
rect 19292 22082 19348 22092
rect 18172 21758 18174 21810
rect 18226 21758 18228 21810
rect 17836 21698 17892 21710
rect 17836 21646 17838 21698
rect 17890 21646 17892 21698
rect 17724 20132 17780 20142
rect 17724 20018 17780 20076
rect 17724 19966 17726 20018
rect 17778 19966 17780 20018
rect 17724 19234 17780 19966
rect 17836 19460 17892 21646
rect 17948 21698 18004 21710
rect 17948 21646 17950 21698
rect 18002 21646 18004 21698
rect 17948 21140 18004 21646
rect 18060 21140 18116 21150
rect 17948 21084 18060 21140
rect 18060 21026 18116 21084
rect 18060 20974 18062 21026
rect 18114 20974 18116 21026
rect 18060 20962 18116 20974
rect 18172 20804 18228 21758
rect 18844 21868 19236 21924
rect 18620 21588 18676 21598
rect 18844 21588 18900 21868
rect 18620 21586 18900 21588
rect 18620 21534 18622 21586
rect 18674 21534 18900 21586
rect 18620 21532 18900 21534
rect 18956 21698 19012 21710
rect 18956 21646 18958 21698
rect 19010 21646 19012 21698
rect 18396 21028 18452 21038
rect 18396 20934 18452 20972
rect 17836 19394 17892 19404
rect 17948 20748 18228 20804
rect 18620 20916 18676 21532
rect 18844 21364 18900 21374
rect 17724 19182 17726 19234
rect 17778 19182 17780 19234
rect 17724 18564 17780 19182
rect 17724 18498 17780 18508
rect 17948 18450 18004 20748
rect 18060 20580 18116 20590
rect 18060 19348 18116 20524
rect 18172 20580 18228 20590
rect 18620 20580 18676 20860
rect 18732 21140 18788 21150
rect 18732 20802 18788 21084
rect 18732 20750 18734 20802
rect 18786 20750 18788 20802
rect 18732 20738 18788 20750
rect 18172 20578 18676 20580
rect 18172 20526 18174 20578
rect 18226 20526 18676 20578
rect 18172 20524 18676 20526
rect 18172 20514 18228 20524
rect 18396 20356 18452 20366
rect 18284 20132 18340 20142
rect 18284 20018 18340 20076
rect 18284 19966 18286 20018
rect 18338 19966 18340 20018
rect 18284 19954 18340 19966
rect 18060 19292 18228 19348
rect 18060 19122 18116 19134
rect 18060 19070 18062 19122
rect 18114 19070 18116 19122
rect 18060 18900 18116 19070
rect 18172 19010 18228 19292
rect 18172 18958 18174 19010
rect 18226 18958 18228 19010
rect 18172 18946 18228 18958
rect 18060 18834 18116 18844
rect 18396 18562 18452 20300
rect 18844 20244 18900 21308
rect 18956 21252 19012 21646
rect 18956 20690 19012 21196
rect 18956 20638 18958 20690
rect 19010 20638 19012 20690
rect 18956 20580 19012 20638
rect 18956 20514 19012 20524
rect 19180 21698 19236 21710
rect 19180 21646 19182 21698
rect 19234 21646 19236 21698
rect 18620 20188 18900 20244
rect 18620 19460 18676 20188
rect 18732 20020 18788 20030
rect 19068 20020 19124 20030
rect 18788 20018 19124 20020
rect 18788 19966 19070 20018
rect 19122 19966 19124 20018
rect 18788 19964 19124 19966
rect 18732 19926 18788 19964
rect 19068 19954 19124 19964
rect 19180 19908 19236 21646
rect 18620 19404 19012 19460
rect 18844 19124 18900 19134
rect 18844 19030 18900 19068
rect 18396 18510 18398 18562
rect 18450 18510 18452 18562
rect 18396 18498 18452 18510
rect 17948 18398 17950 18450
rect 18002 18398 18004 18450
rect 17948 18386 18004 18398
rect 17612 18172 18116 18228
rect 17724 17668 17780 17678
rect 17724 17574 17780 17612
rect 17948 17556 18004 17566
rect 17836 17554 18004 17556
rect 17836 17502 17950 17554
rect 18002 17502 18004 17554
rect 17836 17500 18004 17502
rect 18060 17556 18116 18172
rect 18172 17780 18228 17790
rect 18172 17778 18676 17780
rect 18172 17726 18174 17778
rect 18226 17726 18676 17778
rect 18172 17724 18676 17726
rect 18172 17714 18228 17724
rect 18620 17666 18676 17724
rect 18620 17614 18622 17666
rect 18674 17614 18676 17666
rect 18620 17602 18676 17614
rect 18956 17666 19012 19404
rect 19180 18676 19236 19852
rect 19180 18610 19236 18620
rect 19292 20580 19348 20590
rect 19292 18228 19348 20524
rect 18956 17614 18958 17666
rect 19010 17614 19012 17666
rect 18284 17556 18340 17566
rect 18060 17554 18340 17556
rect 18060 17502 18286 17554
rect 18338 17502 18340 17554
rect 18060 17500 18340 17502
rect 14700 17332 14756 17342
rect 14700 16994 14756 17276
rect 17836 17108 17892 17500
rect 17948 17490 18004 17500
rect 14700 16942 14702 16994
rect 14754 16942 14756 16994
rect 14700 16930 14756 16942
rect 16828 17052 17892 17108
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 14028 13746 14084 16828
rect 16044 16884 16100 16894
rect 14700 15316 14756 15326
rect 14700 13858 14756 15260
rect 16044 14530 16100 16828
rect 16828 16770 16884 17052
rect 16828 16718 16830 16770
rect 16882 16718 16884 16770
rect 16828 16706 16884 16718
rect 16828 15876 16884 15886
rect 16716 15204 16772 15214
rect 16716 14642 16772 15148
rect 16716 14590 16718 14642
rect 16770 14590 16772 14642
rect 16716 14578 16772 14590
rect 16044 14478 16046 14530
rect 16098 14478 16100 14530
rect 16044 14466 16100 14478
rect 14700 13806 14702 13858
rect 14754 13806 14756 13858
rect 14700 13794 14756 13806
rect 14028 13694 14030 13746
rect 14082 13694 14084 13746
rect 14028 13682 14084 13694
rect 16828 13634 16884 15820
rect 17164 15148 17220 17052
rect 16940 15092 17220 15148
rect 17500 16884 17556 16894
rect 16940 13748 16996 15092
rect 17500 13972 17556 16828
rect 17836 16210 17892 16222
rect 17836 16158 17838 16210
rect 17890 16158 17892 16210
rect 17724 15876 17780 15886
rect 17724 15782 17780 15820
rect 17612 15540 17668 15550
rect 17612 15314 17668 15484
rect 17612 15262 17614 15314
rect 17666 15262 17668 15314
rect 17612 15250 17668 15262
rect 17724 15316 17780 15326
rect 17724 15222 17780 15260
rect 17836 15314 17892 16158
rect 17948 16100 18004 16110
rect 18172 16100 18228 17500
rect 18284 17490 18340 17500
rect 18508 17444 18564 17454
rect 18508 17106 18564 17388
rect 18844 17442 18900 17454
rect 18844 17390 18846 17442
rect 18898 17390 18900 17442
rect 18732 17332 18788 17342
rect 18844 17332 18900 17390
rect 18788 17276 18900 17332
rect 18732 17266 18788 17276
rect 18956 17220 19012 17614
rect 19068 18172 19348 18228
rect 19404 18450 19460 22092
rect 19628 21810 19684 22316
rect 20300 22370 20356 22382
rect 20300 22318 20302 22370
rect 20354 22318 20356 22370
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19628 21758 19630 21810
rect 19682 21758 19684 21810
rect 19628 21746 19684 21758
rect 19628 21028 19684 21038
rect 19628 20244 19684 20972
rect 20076 20916 20132 20926
rect 20300 20916 20356 22318
rect 21420 22260 21476 24558
rect 21980 23940 22036 23950
rect 21420 22194 21476 22204
rect 21756 22372 21812 22382
rect 21980 22372 22036 23884
rect 21756 22370 22036 22372
rect 21756 22318 21758 22370
rect 21810 22318 22036 22370
rect 21756 22316 22036 22318
rect 22092 23716 22148 23726
rect 22204 23716 22260 24670
rect 22148 23660 22260 23716
rect 22316 25060 22372 25070
rect 20132 20860 20356 20916
rect 20524 21812 20580 21822
rect 20524 21586 20580 21756
rect 21644 21698 21700 21710
rect 21644 21646 21646 21698
rect 21698 21646 21700 21698
rect 21644 21588 21700 21646
rect 21756 21698 21812 22316
rect 21868 22148 21924 22158
rect 21924 22092 22036 22148
rect 21868 22054 21924 22092
rect 21756 21646 21758 21698
rect 21810 21646 21812 21698
rect 21756 21634 21812 21646
rect 21868 21700 21924 21710
rect 21868 21606 21924 21644
rect 20524 21534 20526 21586
rect 20578 21534 20580 21586
rect 20076 20822 20132 20860
rect 20524 20804 20580 21534
rect 21420 21532 21644 21588
rect 20972 21476 21028 21486
rect 20972 21382 21028 21420
rect 20188 20802 20580 20804
rect 20188 20750 20526 20802
rect 20578 20750 20580 20802
rect 20188 20748 20580 20750
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20244 20244 20748
rect 20524 20738 20580 20748
rect 19628 20188 19908 20244
rect 19852 19346 19908 20188
rect 19852 19294 19854 19346
rect 19906 19294 19908 19346
rect 19852 19282 19908 19294
rect 20076 20188 20244 20244
rect 19740 19236 19796 19246
rect 19516 19234 19796 19236
rect 19516 19182 19742 19234
rect 19794 19182 19796 19234
rect 19516 19180 19796 19182
rect 19516 18900 19572 19180
rect 19740 19170 19796 19180
rect 20076 19234 20132 20188
rect 21420 19346 21476 21532
rect 21644 21522 21700 21532
rect 21756 21474 21812 21486
rect 21756 21422 21758 21474
rect 21810 21422 21812 21474
rect 21420 19294 21422 19346
rect 21474 19294 21476 19346
rect 21420 19282 21476 19294
rect 21532 20578 21588 20590
rect 21532 20526 21534 20578
rect 21586 20526 21588 20578
rect 20076 19182 20078 19234
rect 20130 19182 20132 19234
rect 20076 19170 20132 19182
rect 19516 18834 19572 18844
rect 19628 19010 19684 19022
rect 19628 18958 19630 19010
rect 19682 18958 19684 19010
rect 19404 18398 19406 18450
rect 19458 18398 19460 18450
rect 19068 17444 19124 18172
rect 19292 18004 19348 18014
rect 19180 17556 19236 17566
rect 19180 17462 19236 17500
rect 19068 17378 19124 17388
rect 18844 17164 19012 17220
rect 18508 17054 18510 17106
rect 18562 17054 18564 17106
rect 18508 16772 18564 17054
rect 18732 17108 18788 17118
rect 18844 17108 18900 17164
rect 18732 17106 18900 17108
rect 18732 17054 18734 17106
rect 18786 17054 18900 17106
rect 18732 17052 18900 17054
rect 18732 17042 18788 17052
rect 19068 16884 19124 16894
rect 19292 16884 19348 17948
rect 19404 17892 19460 18398
rect 19404 17826 19460 17836
rect 19516 18676 19572 18686
rect 19404 17442 19460 17454
rect 19404 17390 19406 17442
rect 19458 17390 19460 17442
rect 19404 17108 19460 17390
rect 19516 17444 19572 18620
rect 19628 17668 19684 18958
rect 21532 19012 21588 20526
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19740 18562 19796 18574
rect 19740 18510 19742 18562
rect 19794 18510 19796 18562
rect 19740 18004 19796 18510
rect 20972 18564 21028 18574
rect 20972 18470 21028 18508
rect 21532 18228 21588 18956
rect 21756 18564 21812 21422
rect 21868 20692 21924 20702
rect 21868 20598 21924 20636
rect 21980 20468 22036 22092
rect 22092 21810 22148 23660
rect 22092 21758 22094 21810
rect 22146 21758 22148 21810
rect 22092 21746 22148 21758
rect 22316 21698 22372 25004
rect 22316 21646 22318 21698
rect 22370 21646 22372 21698
rect 22316 21634 22372 21646
rect 22428 24834 22484 25116
rect 22652 24948 22708 24958
rect 22652 24854 22708 24892
rect 22428 24782 22430 24834
rect 22482 24782 22484 24834
rect 22428 21476 22484 24782
rect 22876 24276 22932 26684
rect 25340 26514 25396 26910
rect 26908 26852 26964 27132
rect 27468 27188 27524 27198
rect 27468 27094 27524 27132
rect 27916 27188 27972 27198
rect 27916 27074 27972 27132
rect 40012 27186 40068 27198
rect 40012 27134 40014 27186
rect 40066 27134 40068 27186
rect 27916 27022 27918 27074
rect 27970 27022 27972 27074
rect 27916 27010 27972 27022
rect 37660 27076 37716 27086
rect 37660 26982 37716 27020
rect 28140 26964 28196 26974
rect 28140 26870 28196 26908
rect 37884 26964 37940 26974
rect 25340 26462 25342 26514
rect 25394 26462 25396 26514
rect 25340 26450 25396 26462
rect 26572 26796 26964 26852
rect 26572 26514 26628 26796
rect 26572 26462 26574 26514
rect 26626 26462 26628 26514
rect 26572 26450 26628 26462
rect 25228 26290 25284 26302
rect 25228 26238 25230 26290
rect 25282 26238 25284 26290
rect 24332 26178 24388 26190
rect 24332 26126 24334 26178
rect 24386 26126 24388 26178
rect 23884 24948 23940 24958
rect 23436 24836 23492 24846
rect 22540 24220 23380 24276
rect 22540 23938 22596 24220
rect 22540 23886 22542 23938
rect 22594 23886 22596 23938
rect 22540 23874 22596 23886
rect 23100 23716 23156 23726
rect 23100 23622 23156 23660
rect 23100 23154 23156 23166
rect 23100 23102 23102 23154
rect 23154 23102 23156 23154
rect 22764 22260 22820 22270
rect 22540 22148 22596 22158
rect 22540 21586 22596 22092
rect 22540 21534 22542 21586
rect 22594 21534 22596 21586
rect 22540 21522 22596 21534
rect 22428 20804 22484 21420
rect 22540 21028 22596 21038
rect 22764 21028 22820 22204
rect 22988 21698 23044 21710
rect 22988 21646 22990 21698
rect 23042 21646 23044 21698
rect 22596 20972 22820 21028
rect 22876 21252 22932 21262
rect 22540 20914 22596 20972
rect 22540 20862 22542 20914
rect 22594 20862 22596 20914
rect 22540 20850 22596 20862
rect 21756 18498 21812 18508
rect 21868 20412 22036 20468
rect 22092 20802 22484 20804
rect 22092 20750 22430 20802
rect 22482 20750 22484 20802
rect 22092 20748 22484 20750
rect 19740 17938 19796 17948
rect 21420 18172 21588 18228
rect 21644 18452 21700 18462
rect 20636 17780 20692 17790
rect 20636 17686 20692 17724
rect 19740 17668 19796 17678
rect 19628 17612 19740 17668
rect 19740 17574 19796 17612
rect 19628 17444 19684 17454
rect 19516 17442 19684 17444
rect 19516 17390 19630 17442
rect 19682 17390 19684 17442
rect 19516 17388 19684 17390
rect 19628 17378 19684 17388
rect 20748 17444 20804 17454
rect 21420 17444 21476 18172
rect 21532 17780 21588 17790
rect 21532 17686 21588 17724
rect 21644 17666 21700 18396
rect 21868 18450 21924 20412
rect 21868 18398 21870 18450
rect 21922 18398 21924 18450
rect 21868 18386 21924 18398
rect 22092 17890 22148 20748
rect 22428 20738 22484 20748
rect 22876 20802 22932 21196
rect 22876 20750 22878 20802
rect 22930 20750 22932 20802
rect 22876 20738 22932 20750
rect 22988 20804 23044 21646
rect 22988 20738 23044 20748
rect 22988 20580 23044 20590
rect 22876 20578 23044 20580
rect 22876 20526 22990 20578
rect 23042 20526 23044 20578
rect 22876 20524 23044 20526
rect 22764 18564 22820 18574
rect 22092 17838 22094 17890
rect 22146 17838 22148 17890
rect 22092 17826 22148 17838
rect 22428 18450 22484 18462
rect 22428 18398 22430 18450
rect 22482 18398 22484 18450
rect 21868 17780 21924 17790
rect 21868 17686 21924 17724
rect 21644 17614 21646 17666
rect 21698 17614 21700 17666
rect 21644 17602 21700 17614
rect 22316 17668 22372 17678
rect 22316 17574 22372 17612
rect 20748 17350 20804 17388
rect 20860 17442 21476 17444
rect 20860 17390 21422 17442
rect 21474 17390 21476 17442
rect 20860 17388 21476 17390
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 17108 19684 17118
rect 19404 17052 19628 17108
rect 19516 16884 19572 16894
rect 19068 16882 19460 16884
rect 19068 16830 19070 16882
rect 19122 16830 19460 16882
rect 19068 16828 19460 16830
rect 19068 16818 19124 16828
rect 17948 16098 18228 16100
rect 17948 16046 17950 16098
rect 18002 16046 18228 16098
rect 17948 16044 18228 16046
rect 18284 16716 18788 16772
rect 18284 16098 18340 16716
rect 18284 16046 18286 16098
rect 18338 16046 18340 16098
rect 17948 16034 18004 16044
rect 18284 16034 18340 16046
rect 18172 15428 18228 15438
rect 18508 15428 18564 15438
rect 18172 15426 18508 15428
rect 18172 15374 18174 15426
rect 18226 15374 18508 15426
rect 18172 15372 18508 15374
rect 18172 15362 18228 15372
rect 18508 15334 18564 15372
rect 17836 15262 17838 15314
rect 17890 15262 17892 15314
rect 17836 15250 17892 15262
rect 18620 15204 18676 15242
rect 18620 15138 18676 15148
rect 17500 13970 17780 13972
rect 17500 13918 17502 13970
rect 17554 13918 17780 13970
rect 17500 13916 17780 13918
rect 17500 13906 17556 13916
rect 16940 13692 17668 13748
rect 16828 13582 16830 13634
rect 16882 13582 16884 13634
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 16828 8428 16884 13582
rect 17612 8428 17668 13692
rect 17724 12962 17780 13916
rect 18732 13858 18788 16716
rect 18844 16660 18900 16670
rect 18844 16566 18900 16604
rect 18956 16100 19012 16110
rect 18956 16006 19012 16044
rect 18844 15876 18900 15886
rect 18844 15426 18900 15820
rect 18844 15374 18846 15426
rect 18898 15374 18900 15426
rect 18844 15362 18900 15374
rect 19180 15874 19236 15886
rect 19180 15822 19182 15874
rect 19234 15822 19236 15874
rect 19068 15314 19124 15326
rect 19068 15262 19070 15314
rect 19122 15262 19124 15314
rect 18732 13806 18734 13858
rect 18786 13806 18788 13858
rect 18732 13794 18788 13806
rect 18844 14642 18900 14654
rect 18844 14590 18846 14642
rect 18898 14590 18900 14642
rect 18508 13636 18564 13646
rect 18508 13074 18564 13580
rect 18844 13524 18900 14590
rect 18956 14532 19012 14542
rect 18956 13970 19012 14476
rect 18956 13918 18958 13970
rect 19010 13918 19012 13970
rect 18956 13906 19012 13918
rect 19068 13970 19124 15262
rect 19180 15090 19236 15822
rect 19180 15038 19182 15090
rect 19234 15038 19236 15090
rect 19180 14308 19236 15038
rect 19292 15540 19348 15550
rect 19292 14530 19348 15484
rect 19292 14478 19294 14530
rect 19346 14478 19348 14530
rect 19292 14466 19348 14478
rect 19404 14532 19460 16828
rect 19516 16770 19572 16828
rect 19516 16718 19518 16770
rect 19570 16718 19572 16770
rect 19516 15538 19572 16718
rect 19516 15486 19518 15538
rect 19570 15486 19572 15538
rect 19516 15204 19572 15486
rect 19628 15540 19684 17052
rect 20748 16100 20804 16110
rect 20860 16100 20916 17388
rect 21420 17378 21476 17388
rect 22204 17556 22260 17566
rect 20748 16098 20916 16100
rect 20748 16046 20750 16098
rect 20802 16046 20916 16098
rect 20748 16044 20916 16046
rect 21644 16660 21700 16670
rect 21644 16098 21700 16604
rect 21644 16046 21646 16098
rect 21698 16046 21700 16098
rect 20748 16034 20804 16044
rect 21644 16034 21700 16046
rect 21756 16100 21812 16110
rect 20412 15876 20468 15886
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19628 15474 19684 15484
rect 19516 15138 19572 15148
rect 19852 15316 19908 15326
rect 19628 15092 19684 15102
rect 19852 15092 19908 15260
rect 20412 15148 20468 15820
rect 21756 15538 21812 16044
rect 21756 15486 21758 15538
rect 21810 15486 21812 15538
rect 21756 15474 21812 15486
rect 21868 15874 21924 15886
rect 21868 15822 21870 15874
rect 21922 15822 21924 15874
rect 21868 15540 21924 15822
rect 21868 15474 21924 15484
rect 21980 15874 22036 15886
rect 21980 15822 21982 15874
rect 22034 15822 22036 15874
rect 21420 15428 21476 15438
rect 21476 15372 21700 15428
rect 21420 15334 21476 15372
rect 19628 15090 19908 15092
rect 19628 15038 19630 15090
rect 19682 15038 19908 15090
rect 19628 15036 19908 15038
rect 19628 15026 19684 15036
rect 19516 14532 19572 14542
rect 19460 14530 19572 14532
rect 19460 14478 19518 14530
rect 19570 14478 19572 14530
rect 19460 14476 19572 14478
rect 19404 14438 19460 14476
rect 19516 14466 19572 14476
rect 19852 14530 19908 15036
rect 19852 14478 19854 14530
rect 19906 14478 19908 14530
rect 19852 14466 19908 14478
rect 20076 15092 20468 15148
rect 21196 15204 21252 15214
rect 19180 14252 19460 14308
rect 19068 13918 19070 13970
rect 19122 13918 19124 13970
rect 19068 13906 19124 13918
rect 19180 13746 19236 13758
rect 19180 13694 19182 13746
rect 19234 13694 19236 13746
rect 19180 13524 19236 13694
rect 19404 13746 19460 14252
rect 19628 14306 19684 14318
rect 19628 14254 19630 14306
rect 19682 14254 19684 14306
rect 19628 13860 19684 14254
rect 19740 14308 19796 14346
rect 20076 14308 20132 15092
rect 21196 14644 21252 15148
rect 21532 14644 21588 14654
rect 21196 14642 21588 14644
rect 21196 14590 21534 14642
rect 21586 14590 21588 14642
rect 21196 14588 21588 14590
rect 20412 14530 20468 14542
rect 20412 14478 20414 14530
rect 20466 14478 20468 14530
rect 20412 14308 20468 14478
rect 20076 14252 20244 14308
rect 19740 14242 19796 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20188 13972 20244 14252
rect 20076 13916 20244 13972
rect 19740 13860 19796 13870
rect 19628 13858 19796 13860
rect 19628 13806 19742 13858
rect 19794 13806 19796 13858
rect 19628 13804 19796 13806
rect 19740 13794 19796 13804
rect 19404 13694 19406 13746
rect 19458 13694 19460 13746
rect 19404 13682 19460 13694
rect 20076 13746 20132 13916
rect 20076 13694 20078 13746
rect 20130 13694 20132 13746
rect 18844 13468 19236 13524
rect 18508 13022 18510 13074
rect 18562 13022 18564 13074
rect 18508 13010 18564 13022
rect 17724 12910 17726 12962
rect 17778 12910 17780 12962
rect 17724 12898 17780 12910
rect 19180 8428 19236 13468
rect 20076 13524 20132 13694
rect 20300 13746 20356 13758
rect 20300 13694 20302 13746
rect 20354 13694 20356 13746
rect 20188 13636 20244 13646
rect 20188 13542 20244 13580
rect 20076 13458 20132 13468
rect 20300 12964 20356 13694
rect 20412 13076 20468 14252
rect 20636 14308 20692 14318
rect 20636 14306 20804 14308
rect 20636 14254 20638 14306
rect 20690 14254 20804 14306
rect 20636 14252 20804 14254
rect 20636 14242 20692 14252
rect 20636 13076 20692 13086
rect 20412 13074 20692 13076
rect 20412 13022 20638 13074
rect 20690 13022 20692 13074
rect 20412 13020 20692 13022
rect 20300 12898 20356 12908
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20636 8428 20692 13020
rect 16828 8372 17556 8428
rect 17612 8372 17892 8428
rect 19180 8372 19684 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 17500 4338 17556 8372
rect 17500 4286 17502 4338
rect 17554 4286 17556 4338
rect 17500 4274 17556 4286
rect 17724 5236 17780 5246
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 17724 980 17780 5180
rect 17836 5122 17892 8372
rect 18732 5236 18788 5246
rect 18732 5142 18788 5180
rect 17836 5070 17838 5122
rect 17890 5070 17892 5122
rect 17836 5058 17892 5070
rect 18508 4116 18564 4126
rect 17500 924 17780 980
rect 18172 4114 18564 4116
rect 18172 4062 18510 4114
rect 18562 4062 18564 4114
rect 18172 4060 18564 4062
rect 17500 800 17556 924
rect 18172 800 18228 4060
rect 18508 4050 18564 4060
rect 18844 3666 18900 3678
rect 18844 3614 18846 3666
rect 18898 3614 18900 3666
rect 18844 800 18900 3614
rect 19628 3556 19684 8372
rect 20412 8372 20692 8428
rect 20748 8428 20804 14252
rect 21196 13748 21252 14588
rect 21532 14532 21588 14588
rect 21532 14466 21588 14476
rect 20972 13746 21252 13748
rect 20972 13694 21198 13746
rect 21250 13694 21252 13746
rect 20972 13692 21252 13694
rect 20972 12402 21028 13692
rect 21196 13682 21252 13692
rect 21532 12964 21588 12974
rect 21644 12964 21700 15372
rect 21868 15316 21924 15326
rect 21868 14530 21924 15260
rect 21980 14644 22036 15822
rect 22092 15876 22148 15886
rect 22092 15782 22148 15820
rect 22204 15874 22260 17500
rect 22428 17108 22484 18398
rect 22652 18452 22708 18462
rect 22652 18358 22708 18396
rect 22764 18450 22820 18508
rect 22764 18398 22766 18450
rect 22818 18398 22820 18450
rect 22764 18386 22820 18398
rect 22540 17666 22596 17678
rect 22876 17668 22932 20524
rect 22988 20514 23044 20524
rect 22540 17614 22542 17666
rect 22594 17614 22596 17666
rect 22540 17444 22596 17614
rect 22540 17378 22596 17388
rect 22764 17612 22932 17668
rect 23100 19906 23156 23102
rect 23324 22484 23380 24220
rect 23436 23938 23492 24780
rect 23884 24162 23940 24892
rect 24332 24836 24388 26126
rect 25228 24948 25284 26238
rect 25452 26290 25508 26302
rect 25452 26238 25454 26290
rect 25506 26238 25508 26290
rect 25452 25508 25508 26238
rect 25900 26292 25956 26302
rect 26348 26292 26404 26302
rect 25900 26290 26404 26292
rect 25900 26238 25902 26290
rect 25954 26238 26350 26290
rect 26402 26238 26404 26290
rect 25900 26236 26404 26238
rect 25900 26226 25956 26236
rect 26348 26226 26404 26236
rect 26684 26290 26740 26302
rect 26684 26238 26686 26290
rect 26738 26238 26740 26290
rect 25452 25442 25508 25452
rect 25228 24882 25284 24892
rect 24332 24770 24388 24780
rect 26124 24834 26180 24846
rect 26124 24782 26126 24834
rect 26178 24782 26180 24834
rect 25788 24724 25844 24734
rect 23884 24110 23886 24162
rect 23938 24110 23940 24162
rect 23884 24098 23940 24110
rect 25564 24668 25788 24724
rect 23436 23886 23438 23938
rect 23490 23886 23492 23938
rect 23436 23874 23492 23886
rect 24108 23938 24164 23950
rect 24108 23886 24110 23938
rect 24162 23886 24164 23938
rect 23436 22484 23492 22494
rect 23324 22482 23492 22484
rect 23324 22430 23438 22482
rect 23490 22430 23492 22482
rect 23324 22428 23492 22430
rect 23436 22418 23492 22428
rect 23324 22146 23380 22158
rect 23324 22094 23326 22146
rect 23378 22094 23380 22146
rect 23324 21812 23380 22094
rect 23324 21746 23380 21756
rect 23212 21700 23268 21710
rect 23212 21606 23268 21644
rect 23996 21588 24052 21598
rect 23996 21494 24052 21532
rect 24108 21252 24164 23886
rect 25116 23940 25172 23950
rect 25116 23938 25508 23940
rect 25116 23886 25118 23938
rect 25170 23886 25508 23938
rect 25116 23884 25508 23886
rect 25116 23874 25172 23884
rect 24332 23826 24388 23838
rect 24332 23774 24334 23826
rect 24386 23774 24388 23826
rect 24332 23268 24388 23774
rect 24332 23202 24388 23212
rect 24444 23826 24500 23838
rect 24444 23774 24446 23826
rect 24498 23774 24500 23826
rect 24444 22708 24500 23774
rect 24668 23828 24724 23838
rect 24668 23826 24836 23828
rect 24668 23774 24670 23826
rect 24722 23774 24836 23826
rect 24668 23772 24836 23774
rect 24668 23762 24724 23772
rect 24780 23604 24836 23772
rect 24780 23538 24836 23548
rect 25004 23714 25060 23726
rect 25004 23662 25006 23714
rect 25058 23662 25060 23714
rect 24108 21186 24164 21196
rect 24220 22652 24500 22708
rect 24668 23492 24724 23502
rect 24668 23378 24724 23436
rect 24668 23326 24670 23378
rect 24722 23326 24724 23378
rect 24220 20692 24276 22652
rect 24332 22484 24388 22494
rect 24668 22484 24724 23326
rect 24332 22482 24724 22484
rect 24332 22430 24334 22482
rect 24386 22430 24724 22482
rect 24332 22428 24724 22430
rect 24332 22418 24388 22428
rect 24668 22370 24724 22428
rect 24668 22318 24670 22370
rect 24722 22318 24724 22370
rect 24668 22306 24724 22318
rect 25004 22372 25060 23662
rect 25228 23716 25284 23754
rect 25228 23650 25284 23660
rect 25228 23492 25284 23502
rect 25228 23154 25284 23436
rect 25228 23102 25230 23154
rect 25282 23102 25284 23154
rect 25228 23090 25284 23102
rect 25452 22482 25508 23884
rect 25564 23716 25620 24668
rect 25788 24630 25844 24668
rect 26124 24164 26180 24782
rect 26124 24108 26628 24164
rect 25676 23996 26068 24052
rect 25676 23938 25732 23996
rect 25676 23886 25678 23938
rect 25730 23886 25732 23938
rect 25676 23874 25732 23886
rect 26012 23940 26068 23996
rect 26460 23940 26516 23950
rect 26012 23938 26516 23940
rect 26012 23886 26462 23938
rect 26514 23886 26516 23938
rect 26012 23884 26516 23886
rect 26460 23874 26516 23884
rect 26572 23940 26628 24108
rect 26684 23940 26740 26238
rect 37884 26290 37940 26908
rect 37884 26238 37886 26290
rect 37938 26238 37940 26290
rect 37884 26226 37940 26238
rect 39900 26852 39956 26862
rect 39900 26178 39956 26796
rect 40012 26292 40068 27134
rect 40012 26226 40068 26236
rect 39900 26126 39902 26178
rect 39954 26126 39956 26178
rect 39900 26114 39956 26126
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 26796 23940 26852 23950
rect 26572 23938 26852 23940
rect 26572 23886 26798 23938
rect 26850 23886 26852 23938
rect 26572 23884 26852 23886
rect 25900 23826 25956 23838
rect 25900 23774 25902 23826
rect 25954 23774 25956 23826
rect 25900 23716 25956 23774
rect 25564 23660 25956 23716
rect 26012 23716 26068 23726
rect 26236 23716 26292 23726
rect 26012 23622 26068 23660
rect 26124 23714 26292 23716
rect 26124 23662 26238 23714
rect 26290 23662 26292 23714
rect 26124 23660 26292 23662
rect 26124 23604 26180 23660
rect 26236 23650 26292 23660
rect 26124 23538 26180 23548
rect 26012 23268 26068 23278
rect 26012 23174 26068 23212
rect 25452 22430 25454 22482
rect 25506 22430 25508 22482
rect 25452 22418 25508 22430
rect 25004 22306 25060 22316
rect 26572 21476 26628 23884
rect 26796 23874 26852 23884
rect 28140 23940 28196 23950
rect 26684 23714 26740 23726
rect 26684 23662 26686 23714
rect 26738 23662 26740 23714
rect 26684 23604 26740 23662
rect 28140 23604 28196 23884
rect 37660 23940 37716 23950
rect 37660 23846 37716 23884
rect 26684 23548 26964 23604
rect 26908 22484 26964 23548
rect 28140 23042 28196 23548
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 28140 22990 28142 23042
rect 28194 22990 28196 23042
rect 28140 22978 28196 22990
rect 37660 23154 37716 23166
rect 37660 23102 37662 23154
rect 37714 23102 37716 23154
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 27020 22484 27076 22494
rect 26908 22428 27020 22484
rect 27020 22418 27076 22428
rect 27580 22484 27636 22494
rect 27580 22390 27636 22428
rect 37660 22484 37716 23102
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 37660 22418 37716 22428
rect 37324 21588 37380 21598
rect 37324 21494 37380 21532
rect 37772 21588 37828 21598
rect 37772 21494 37828 21532
rect 26572 21410 26628 21420
rect 27692 21476 27748 21486
rect 26348 20804 26404 20814
rect 26348 20710 26404 20748
rect 27244 20802 27300 20814
rect 27244 20750 27246 20802
rect 27298 20750 27300 20802
rect 24220 20626 24276 20636
rect 25900 20692 25956 20702
rect 25900 20598 25956 20636
rect 26796 20692 26852 20702
rect 26796 20598 26852 20636
rect 25228 20578 25284 20590
rect 25228 20526 25230 20578
rect 25282 20526 25284 20578
rect 25228 20020 25284 20526
rect 25676 20580 25732 20590
rect 25676 20486 25732 20524
rect 25788 20578 25844 20590
rect 25788 20526 25790 20578
rect 25842 20526 25844 20578
rect 25788 20244 25844 20526
rect 26572 20578 26628 20590
rect 26572 20526 26574 20578
rect 26626 20526 26628 20578
rect 25788 20188 26292 20244
rect 26236 20130 26292 20188
rect 26236 20078 26238 20130
rect 26290 20078 26292 20130
rect 26236 20066 26292 20078
rect 25452 20020 25508 20030
rect 25228 20018 25508 20020
rect 25228 19966 25454 20018
rect 25506 19966 25508 20018
rect 25228 19964 25508 19966
rect 23100 19854 23102 19906
rect 23154 19854 23156 19906
rect 22428 17042 22484 17052
rect 22764 16100 22820 17612
rect 22988 17554 23044 17566
rect 22988 17502 22990 17554
rect 23042 17502 23044 17554
rect 22876 17442 22932 17454
rect 22876 17390 22878 17442
rect 22930 17390 22932 17442
rect 22876 16212 22932 17390
rect 22988 17108 23044 17502
rect 22988 17042 23044 17052
rect 23100 16882 23156 19854
rect 24220 19234 24276 19246
rect 24220 19182 24222 19234
rect 24274 19182 24276 19234
rect 23548 19124 23604 19134
rect 23548 19122 23716 19124
rect 23548 19070 23550 19122
rect 23602 19070 23716 19122
rect 23548 19068 23716 19070
rect 23548 19058 23604 19068
rect 23660 18674 23716 19068
rect 23660 18622 23662 18674
rect 23714 18622 23716 18674
rect 23660 18610 23716 18622
rect 24220 19012 24276 19182
rect 25452 19234 25508 19964
rect 26572 19908 26628 20526
rect 25452 19182 25454 19234
rect 25506 19182 25508 19234
rect 23884 18452 23940 18462
rect 23772 18450 23940 18452
rect 23772 18398 23886 18450
rect 23938 18398 23940 18450
rect 23772 18396 23940 18398
rect 23212 18228 23268 18238
rect 23548 18228 23604 18238
rect 23212 18226 23604 18228
rect 23212 18174 23214 18226
rect 23266 18174 23550 18226
rect 23602 18174 23604 18226
rect 23212 18172 23604 18174
rect 23212 18162 23268 18172
rect 23548 18162 23604 18172
rect 23100 16830 23102 16882
rect 23154 16830 23156 16882
rect 23100 16818 23156 16830
rect 23212 17556 23268 17566
rect 23212 16212 23268 17500
rect 23772 17556 23828 18396
rect 23884 18386 23940 18396
rect 23772 17490 23828 17500
rect 22876 16146 22932 16156
rect 22988 16156 23268 16212
rect 22764 16006 22820 16044
rect 22988 15986 23044 16156
rect 22988 15934 22990 15986
rect 23042 15934 23044 15986
rect 22988 15922 23044 15934
rect 23996 16100 24052 16110
rect 24220 16100 24276 18956
rect 25004 19012 25060 19022
rect 25004 18918 25060 18956
rect 25452 19012 25508 19182
rect 25452 18946 25508 18956
rect 26012 19852 26628 19908
rect 26684 20578 26740 20590
rect 26684 20526 26686 20578
rect 26738 20526 26740 20578
rect 25900 18452 25956 18462
rect 26012 18452 26068 19852
rect 26684 19796 26740 20526
rect 26124 19740 26740 19796
rect 27244 19796 27300 20750
rect 27356 20804 27412 20814
rect 27356 20710 27412 20748
rect 27692 20690 27748 21420
rect 39900 21474 39956 21486
rect 39900 21422 39902 21474
rect 39954 21422 39956 21474
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 39900 20916 39956 21422
rect 39900 20850 39956 20860
rect 40012 20914 40068 20926
rect 40012 20862 40014 20914
rect 40066 20862 40068 20914
rect 37660 20804 37716 20814
rect 37660 20710 37716 20748
rect 27692 20638 27694 20690
rect 27746 20638 27748 20690
rect 27580 20580 27636 20590
rect 27580 20486 27636 20524
rect 27692 20468 27748 20638
rect 27692 20402 27748 20412
rect 28364 20580 28420 20590
rect 26124 19346 26180 19740
rect 27244 19730 27300 19740
rect 28252 20132 28308 20142
rect 26124 19294 26126 19346
rect 26178 19294 26180 19346
rect 26124 19282 26180 19294
rect 28252 19346 28308 20076
rect 28364 19906 28420 20524
rect 28700 20468 28756 20478
rect 28700 20130 28756 20412
rect 40012 20244 40068 20862
rect 40012 20178 40068 20188
rect 28700 20078 28702 20130
rect 28754 20078 28756 20130
rect 28700 20066 28756 20078
rect 28812 20132 28868 20142
rect 28812 20038 28868 20076
rect 37660 20020 37716 20030
rect 37660 19926 37716 19964
rect 28364 19854 28366 19906
rect 28418 19854 28420 19906
rect 28364 19842 28420 19854
rect 28812 19796 28868 19806
rect 28812 19702 28868 19740
rect 40012 19794 40068 19806
rect 40012 19742 40014 19794
rect 40066 19742 40068 19794
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 40012 19572 40068 19742
rect 40012 19506 40068 19516
rect 28252 19294 28254 19346
rect 28306 19294 28308 19346
rect 28252 19282 28308 19294
rect 25956 18396 26068 18452
rect 25900 18386 25956 18396
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 26012 17780 26068 17790
rect 26012 17686 26068 17724
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 26124 17668 26180 17678
rect 26124 17574 26180 17612
rect 26908 17668 26964 17678
rect 24780 16212 24836 16222
rect 24780 16118 24836 16156
rect 26908 16210 26964 17612
rect 37660 17668 37716 17678
rect 37660 17574 37716 17612
rect 40012 17556 40068 17726
rect 40012 17490 40068 17500
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 26908 16158 26910 16210
rect 26962 16158 26964 16210
rect 26908 16146 26964 16158
rect 23996 16098 24276 16100
rect 23996 16046 23998 16098
rect 24050 16046 24276 16098
rect 23996 16044 24276 16046
rect 22204 15822 22206 15874
rect 22258 15822 22260 15874
rect 22204 15810 22260 15822
rect 22316 15876 22372 15886
rect 21980 14578 22036 14588
rect 21868 14478 21870 14530
rect 21922 14478 21924 14530
rect 21868 14466 21924 14478
rect 22316 14530 22372 15820
rect 23660 15876 23716 15886
rect 23996 15876 24052 16044
rect 23660 15874 24052 15876
rect 23660 15822 23662 15874
rect 23714 15822 24052 15874
rect 23660 15820 24052 15822
rect 22652 15540 22708 15550
rect 22708 15484 22820 15540
rect 22652 15474 22708 15484
rect 22540 15428 22596 15438
rect 22540 15334 22596 15372
rect 22764 15426 22820 15484
rect 22764 15374 22766 15426
rect 22818 15374 22820 15426
rect 22764 15362 22820 15374
rect 22428 15316 22484 15326
rect 22428 15222 22484 15260
rect 23548 14644 23604 14654
rect 23548 14550 23604 14588
rect 22316 14478 22318 14530
rect 22370 14478 22372 14530
rect 22316 14466 22372 14478
rect 22764 14532 22820 14542
rect 22764 14438 22820 14476
rect 22204 14418 22260 14430
rect 22204 14366 22206 14418
rect 22258 14366 22260 14418
rect 22092 14306 22148 14318
rect 22092 14254 22094 14306
rect 22146 14254 22148 14306
rect 21980 13636 22036 13646
rect 21756 13634 22036 13636
rect 21756 13582 21982 13634
rect 22034 13582 22036 13634
rect 21756 13580 22036 13582
rect 21756 13074 21812 13580
rect 21980 13570 22036 13580
rect 21756 13022 21758 13074
rect 21810 13022 21812 13074
rect 21756 13010 21812 13022
rect 21868 13412 21924 13422
rect 21588 12908 21700 12964
rect 21868 12962 21924 13356
rect 21868 12910 21870 12962
rect 21922 12910 21924 12962
rect 21532 12870 21588 12908
rect 21868 12898 21924 12910
rect 22092 12962 22148 14254
rect 22204 13636 22260 14366
rect 23660 14308 23716 15820
rect 25228 15428 25284 15438
rect 25284 15372 25396 15428
rect 25228 15334 25284 15372
rect 25340 14644 25396 15372
rect 25564 15426 25620 15438
rect 25564 15374 25566 15426
rect 25618 15374 25620 15426
rect 25564 15148 25620 15374
rect 25564 15092 25844 15148
rect 25676 14644 25732 14654
rect 25340 14642 25732 14644
rect 25340 14590 25678 14642
rect 25730 14590 25732 14642
rect 25340 14588 25732 14590
rect 23660 14242 23716 14252
rect 24556 14308 24612 14318
rect 24556 13970 24612 14252
rect 24556 13918 24558 13970
rect 24610 13918 24612 13970
rect 24556 13906 24612 13918
rect 22204 13570 22260 13580
rect 24108 13636 24164 13646
rect 22092 12910 22094 12962
rect 22146 12910 22148 12962
rect 22092 12898 22148 12910
rect 20972 12350 20974 12402
rect 21026 12350 21028 12402
rect 20972 12338 21028 12350
rect 24108 8428 24164 13580
rect 20748 8372 21140 8428
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 20412 4338 20468 8372
rect 20412 4286 20414 4338
rect 20466 4286 20468 4338
rect 20412 4274 20468 4286
rect 20188 4116 20244 4126
rect 19740 3556 19796 3566
rect 19628 3554 19796 3556
rect 19628 3502 19742 3554
rect 19794 3502 19796 3554
rect 19628 3500 19796 3502
rect 19740 3490 19796 3500
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 800 20244 4060
rect 20860 3668 20916 3678
rect 20860 800 20916 3612
rect 21084 3554 21140 8372
rect 23772 8372 24164 8428
rect 23548 5236 23604 5246
rect 21420 4116 21476 4126
rect 21420 4022 21476 4060
rect 22092 3668 22148 3678
rect 22092 3574 22148 3612
rect 22876 3668 22932 3678
rect 21084 3502 21086 3554
rect 21138 3502 21140 3554
rect 21084 3490 21140 3502
rect 22876 800 22932 3612
rect 23548 800 23604 5180
rect 23772 5122 23828 8372
rect 24780 5236 24836 5246
rect 24780 5142 24836 5180
rect 23772 5070 23774 5122
rect 23826 5070 23828 5122
rect 23772 5058 23828 5070
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 25004 3556 25060 3566
rect 25004 3462 25060 3500
rect 25676 3556 25732 14588
rect 25788 4338 25844 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 25788 4286 25790 4338
rect 25842 4286 25844 4338
rect 25788 4274 25844 4286
rect 25676 3490 25732 3500
rect 25788 4116 25844 4126
rect 25788 980 25844 4060
rect 26796 4116 26852 4126
rect 26796 4022 26852 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 25564 924 25844 980
rect 25564 800 25620 924
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 22848 0 22960 800
rect 23520 0 23632 800
rect 25536 0 25648 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 17500 38220 17556 38276
rect 18620 38274 18676 38276
rect 18620 38222 18622 38274
rect 18622 38222 18674 38274
rect 18674 38222 18676 38274
rect 18620 38220 18676 38222
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 22876 38220 22932 38276
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 16828 37436 16884 37492
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4172 27580 4228 27636
rect 1932 26236 1988 26292
rect 1932 25564 1988 25620
rect 2044 24892 2100 24948
rect 1932 23548 1988 23604
rect 1932 22930 1988 22932
rect 1932 22878 1934 22930
rect 1934 22878 1986 22930
rect 1986 22878 1988 22930
rect 1932 22876 1988 22878
rect 1932 21532 1988 21588
rect 15148 27580 15204 27636
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4284 27074 4340 27076
rect 4284 27022 4286 27074
rect 4286 27022 4338 27074
rect 4338 27022 4340 27074
rect 4284 27020 4340 27022
rect 12124 27020 12180 27076
rect 4284 26290 4340 26292
rect 4284 26238 4286 26290
rect 4286 26238 4338 26290
rect 4338 26238 4340 26290
rect 4284 26236 4340 26238
rect 12124 26236 12180 26292
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4284 25506 4340 25508
rect 4284 25454 4286 25506
rect 4286 25454 4338 25506
rect 4338 25454 4340 25506
rect 4284 25452 4340 25454
rect 11676 25730 11732 25732
rect 11676 25678 11678 25730
rect 11678 25678 11730 25730
rect 11730 25678 11732 25730
rect 11676 25676 11732 25678
rect 10220 25452 10276 25508
rect 11676 25394 11732 25396
rect 11676 25342 11678 25394
rect 11678 25342 11730 25394
rect 11730 25342 11732 25394
rect 11676 25340 11732 25342
rect 12348 25676 12404 25732
rect 13132 26290 13188 26292
rect 13132 26238 13134 26290
rect 13134 26238 13186 26290
rect 13186 26238 13188 26290
rect 13132 26236 13188 26238
rect 13804 26290 13860 26292
rect 13804 26238 13806 26290
rect 13806 26238 13858 26290
rect 13858 26238 13860 26290
rect 13804 26236 13860 26238
rect 12348 25506 12404 25508
rect 12348 25454 12350 25506
rect 12350 25454 12402 25506
rect 12402 25454 12404 25506
rect 12348 25452 12404 25454
rect 13804 25116 13860 25172
rect 16828 26908 16884 26964
rect 16156 26236 16212 26292
rect 14476 26178 14532 26180
rect 14476 26126 14478 26178
rect 14478 26126 14530 26178
rect 14530 26126 14532 26178
rect 14476 26124 14532 26126
rect 16044 26124 16100 26180
rect 16604 26178 16660 26180
rect 16604 26126 16606 26178
rect 16606 26126 16658 26178
rect 16658 26126 16660 26178
rect 16604 26124 16660 26126
rect 16604 25564 16660 25620
rect 15932 25282 15988 25284
rect 15932 25230 15934 25282
rect 15934 25230 15986 25282
rect 15986 25230 15988 25282
rect 15932 25228 15988 25230
rect 14476 25116 14532 25172
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4284 23772 4340 23828
rect 13468 23772 13524 23828
rect 12684 23548 12740 23604
rect 13468 23436 13524 23492
rect 11004 23212 11060 23268
rect 4284 23154 4340 23156
rect 4284 23102 4286 23154
rect 4286 23102 4338 23154
rect 4338 23102 4340 23154
rect 4284 23100 4340 23102
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 13132 22540 13188 22596
rect 12908 21756 12964 21812
rect 4284 21420 4340 21476
rect 9996 21644 10052 21700
rect 13356 21698 13412 21700
rect 13356 21646 13358 21698
rect 13358 21646 13410 21698
rect 13410 21646 13412 21698
rect 13356 21644 13412 21646
rect 14252 23436 14308 23492
rect 15484 23548 15540 23604
rect 15372 23378 15428 23380
rect 15372 23326 15374 23378
rect 15374 23326 15426 23378
rect 15426 23326 15428 23378
rect 15372 23324 15428 23326
rect 14364 23266 14420 23268
rect 14364 23214 14366 23266
rect 14366 23214 14418 23266
rect 14418 23214 14420 23266
rect 14364 23212 14420 23214
rect 14812 23042 14868 23044
rect 14812 22990 14814 23042
rect 14814 22990 14866 23042
rect 14866 22990 14868 23042
rect 14812 22988 14868 22990
rect 15596 23042 15652 23044
rect 15596 22990 15598 23042
rect 15598 22990 15650 23042
rect 15650 22990 15652 23042
rect 15596 22988 15652 22990
rect 14364 22930 14420 22932
rect 14364 22878 14366 22930
rect 14366 22878 14418 22930
rect 14418 22878 14420 22930
rect 14364 22876 14420 22878
rect 15260 22876 15316 22932
rect 15484 22594 15540 22596
rect 15484 22542 15486 22594
rect 15486 22542 15538 22594
rect 15538 22542 15540 22594
rect 15484 22540 15540 22542
rect 13916 21810 13972 21812
rect 13916 21758 13918 21810
rect 13918 21758 13970 21810
rect 13970 21758 13972 21810
rect 13916 21756 13972 21758
rect 15596 21756 15652 21812
rect 16268 25116 16324 25172
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 18396 37490 18452 37492
rect 18396 37438 18398 37490
rect 18398 37438 18450 37490
rect 18450 37438 18452 37490
rect 18396 37436 18452 37438
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 17388 27634 17444 27636
rect 17388 27582 17390 27634
rect 17390 27582 17442 27634
rect 17442 27582 17444 27634
rect 17388 27580 17444 27582
rect 17612 26908 17668 26964
rect 17164 26796 17220 26852
rect 17500 26796 17556 26852
rect 17052 26124 17108 26180
rect 16940 25618 16996 25620
rect 16940 25566 16942 25618
rect 16942 25566 16994 25618
rect 16994 25566 16996 25618
rect 16940 25564 16996 25566
rect 17276 25394 17332 25396
rect 17276 25342 17278 25394
rect 17278 25342 17330 25394
rect 17330 25342 17332 25394
rect 17276 25340 17332 25342
rect 16828 25116 16884 25172
rect 16268 23938 16324 23940
rect 16268 23886 16270 23938
rect 16270 23886 16322 23938
rect 16322 23886 16324 23938
rect 16268 23884 16324 23886
rect 18284 27746 18340 27748
rect 18284 27694 18286 27746
rect 18286 27694 18338 27746
rect 18338 27694 18340 27746
rect 18284 27692 18340 27694
rect 20412 27746 20468 27748
rect 20412 27694 20414 27746
rect 20414 27694 20466 27746
rect 20466 27694 20468 27746
rect 20412 27692 20468 27694
rect 20412 27020 20468 27076
rect 18284 26908 18340 26964
rect 18732 26514 18788 26516
rect 18732 26462 18734 26514
rect 18734 26462 18786 26514
rect 18786 26462 18788 26514
rect 18732 26460 18788 26462
rect 20524 26796 20580 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20636 26684 20692 26740
rect 22764 27692 22820 27748
rect 21532 27074 21588 27076
rect 21532 27022 21534 27074
rect 21534 27022 21586 27074
rect 21586 27022 21588 27074
rect 21532 27020 21588 27022
rect 20044 26628 20100 26630
rect 19628 26514 19684 26516
rect 19628 26462 19630 26514
rect 19630 26462 19682 26514
rect 19682 26462 19684 26514
rect 19628 26460 19684 26462
rect 17500 25506 17556 25508
rect 17500 25454 17502 25506
rect 17502 25454 17554 25506
rect 17554 25454 17556 25506
rect 17500 25452 17556 25454
rect 17388 25228 17444 25284
rect 18956 26290 19012 26292
rect 18956 26238 18958 26290
rect 18958 26238 19010 26290
rect 19010 26238 19012 26290
rect 18956 26236 19012 26238
rect 18284 25340 18340 25396
rect 18396 24780 18452 24836
rect 17612 24108 17668 24164
rect 18172 24108 18228 24164
rect 17500 23938 17556 23940
rect 17500 23886 17502 23938
rect 17502 23886 17554 23938
rect 17554 23886 17556 23938
rect 17500 23884 17556 23886
rect 16940 23548 16996 23604
rect 17612 23660 17668 23716
rect 16716 23324 16772 23380
rect 15820 22258 15876 22260
rect 15820 22206 15822 22258
rect 15822 22206 15874 22258
rect 15874 22206 15876 22258
rect 15820 22204 15876 22206
rect 15708 22092 15764 22148
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 12460 21196 12516 21252
rect 15148 20748 15204 20804
rect 13020 20130 13076 20132
rect 13020 20078 13022 20130
rect 13022 20078 13074 20130
rect 13074 20078 13076 20130
rect 13020 20076 13076 20078
rect 4172 19964 4228 20020
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 15484 20076 15540 20132
rect 15484 19404 15540 19460
rect 12236 18956 12292 19012
rect 14028 18956 14084 19012
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 13804 18284 13860 18340
rect 15372 19010 15428 19012
rect 15372 18958 15374 19010
rect 15374 18958 15426 19010
rect 15426 18958 15428 19010
rect 15372 18956 15428 18958
rect 15036 18844 15092 18900
rect 15932 20748 15988 20804
rect 16156 22316 16212 22372
rect 17388 21196 17444 21252
rect 17500 21644 17556 21700
rect 16268 20748 16324 20804
rect 16156 20300 16212 20356
rect 16828 20802 16884 20804
rect 16828 20750 16830 20802
rect 16830 20750 16882 20802
rect 16882 20750 16884 20802
rect 16828 20748 16884 20750
rect 16940 20188 16996 20244
rect 15820 20130 15876 20132
rect 15820 20078 15822 20130
rect 15822 20078 15874 20130
rect 15874 20078 15876 20130
rect 15820 20076 15876 20078
rect 16604 19852 16660 19908
rect 15820 19458 15876 19460
rect 15820 19406 15822 19458
rect 15822 19406 15874 19458
rect 15874 19406 15876 19458
rect 15820 19404 15876 19406
rect 15932 19234 15988 19236
rect 15932 19182 15934 19234
rect 15934 19182 15986 19234
rect 15986 19182 15988 19234
rect 15932 19180 15988 19182
rect 16604 19234 16660 19236
rect 16604 19182 16606 19234
rect 16606 19182 16658 19234
rect 16658 19182 16660 19234
rect 16604 19180 16660 19182
rect 15708 18844 15764 18900
rect 16828 19010 16884 19012
rect 16828 18958 16830 19010
rect 16830 18958 16882 19010
rect 16882 18958 16884 19010
rect 16828 18956 16884 18958
rect 15932 18396 15988 18452
rect 17388 20300 17444 20356
rect 17500 20188 17556 20244
rect 17276 20076 17332 20132
rect 17164 18844 17220 18900
rect 15820 18338 15876 18340
rect 15820 18286 15822 18338
rect 15822 18286 15874 18338
rect 15874 18286 15876 18338
rect 15820 18284 15876 18286
rect 17948 22482 18004 22484
rect 17948 22430 17950 22482
rect 17950 22430 18002 22482
rect 18002 22430 18004 22482
rect 17948 22428 18004 22430
rect 17724 22204 17780 22260
rect 18060 21810 18116 21812
rect 18060 21758 18062 21810
rect 18062 21758 18114 21810
rect 18114 21758 18116 21810
rect 18060 21756 18116 21758
rect 18396 23660 18452 23716
rect 18844 25452 18900 25508
rect 21308 26460 21364 26516
rect 21644 26908 21700 26964
rect 22092 27074 22148 27076
rect 22092 27022 22094 27074
rect 22094 27022 22146 27074
rect 22146 27022 22148 27074
rect 22092 27020 22148 27022
rect 23548 27746 23604 27748
rect 23548 27694 23550 27746
rect 23550 27694 23602 27746
rect 23602 27694 23604 27746
rect 23548 27692 23604 27694
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 24556 27692 24612 27748
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 26908 27132 26964 27188
rect 22764 27020 22820 27076
rect 22540 26460 22596 26516
rect 21532 25564 21588 25620
rect 19292 25340 19348 25396
rect 22428 25506 22484 25508
rect 22428 25454 22430 25506
rect 22430 25454 22482 25506
rect 22482 25454 22484 25506
rect 22428 25452 22484 25454
rect 18956 24892 19012 24948
rect 19068 24108 19124 24164
rect 18732 23884 18788 23940
rect 18508 22370 18564 22372
rect 18508 22318 18510 22370
rect 18510 22318 18562 22370
rect 18562 22318 18564 22370
rect 18508 22316 18564 22318
rect 18620 23772 18676 23828
rect 21756 25228 21812 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19852 24834 19908 24836
rect 19852 24782 19854 24834
rect 19854 24782 19906 24834
rect 19906 24782 19908 24834
rect 19852 24780 19908 24782
rect 20636 24834 20692 24836
rect 20636 24782 20638 24834
rect 20638 24782 20690 24834
rect 20690 24782 20692 24834
rect 20636 24780 20692 24782
rect 21868 24834 21924 24836
rect 21868 24782 21870 24834
rect 21870 24782 21922 24834
rect 21922 24782 21924 24834
rect 21868 24780 21924 24782
rect 19740 24668 19796 24724
rect 19628 23938 19684 23940
rect 19628 23886 19630 23938
rect 19630 23886 19682 23938
rect 19682 23886 19684 23938
rect 19628 23884 19684 23886
rect 19180 23772 19236 23828
rect 19852 23996 19908 24052
rect 24220 26962 24276 26964
rect 24220 26910 24222 26962
rect 24222 26910 24274 26962
rect 24274 26910 24276 26962
rect 24220 26908 24276 26910
rect 24668 26908 24724 26964
rect 22876 26684 22932 26740
rect 20076 23884 20132 23940
rect 20524 23996 20580 24052
rect 18732 23660 18788 23716
rect 20188 23826 20244 23828
rect 20188 23774 20190 23826
rect 20190 23774 20242 23826
rect 20242 23774 20244 23826
rect 20188 23772 20244 23774
rect 19628 23548 19684 23604
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 18620 22428 18676 22484
rect 19628 22316 19684 22372
rect 17724 20076 17780 20132
rect 18060 21084 18116 21140
rect 18396 21026 18452 21028
rect 18396 20974 18398 21026
rect 18398 20974 18450 21026
rect 18450 20974 18452 21026
rect 18396 20972 18452 20974
rect 17836 19404 17892 19460
rect 18844 21308 18900 21364
rect 18620 20860 18676 20916
rect 17724 18508 17780 18564
rect 18060 20524 18116 20580
rect 18732 21084 18788 21140
rect 18396 20300 18452 20356
rect 18284 20076 18340 20132
rect 18060 18844 18116 18900
rect 18956 21196 19012 21252
rect 18956 20524 19012 20580
rect 18732 20018 18788 20020
rect 18732 19966 18734 20018
rect 18734 19966 18786 20018
rect 18786 19966 18788 20018
rect 18732 19964 18788 19966
rect 19180 19852 19236 19908
rect 18844 19122 18900 19124
rect 18844 19070 18846 19122
rect 18846 19070 18898 19122
rect 18898 19070 18900 19122
rect 18844 19068 18900 19070
rect 17724 17666 17780 17668
rect 17724 17614 17726 17666
rect 17726 17614 17778 17666
rect 17778 17614 17780 17666
rect 17724 17612 17780 17614
rect 19180 18620 19236 18676
rect 19292 20578 19348 20580
rect 19292 20526 19294 20578
rect 19294 20526 19346 20578
rect 19346 20526 19348 20578
rect 19292 20524 19348 20526
rect 14700 17276 14756 17332
rect 14028 16882 14084 16884
rect 14028 16830 14030 16882
rect 14030 16830 14082 16882
rect 14082 16830 14084 16882
rect 14028 16828 14084 16830
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 16044 16828 16100 16884
rect 14700 15260 14756 15316
rect 16828 15820 16884 15876
rect 16716 15148 16772 15204
rect 17500 16882 17556 16884
rect 17500 16830 17502 16882
rect 17502 16830 17554 16882
rect 17554 16830 17556 16882
rect 17500 16828 17556 16830
rect 17724 15874 17780 15876
rect 17724 15822 17726 15874
rect 17726 15822 17778 15874
rect 17778 15822 17780 15874
rect 17724 15820 17780 15822
rect 17612 15484 17668 15540
rect 17724 15314 17780 15316
rect 17724 15262 17726 15314
rect 17726 15262 17778 15314
rect 17778 15262 17780 15314
rect 17724 15260 17780 15262
rect 18508 17388 18564 17444
rect 18732 17276 18788 17332
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19628 20972 19684 21028
rect 21980 23938 22036 23940
rect 21980 23886 21982 23938
rect 21982 23886 22034 23938
rect 22034 23886 22036 23938
rect 21980 23884 22036 23886
rect 21420 22204 21476 22260
rect 22092 23660 22148 23716
rect 22316 25004 22372 25060
rect 20076 20914 20132 20916
rect 20076 20862 20078 20914
rect 20078 20862 20130 20914
rect 20130 20862 20132 20914
rect 20076 20860 20132 20862
rect 20524 21756 20580 21812
rect 21868 22146 21924 22148
rect 21868 22094 21870 22146
rect 21870 22094 21922 22146
rect 21922 22094 21924 22146
rect 21868 22092 21924 22094
rect 21868 21698 21924 21700
rect 21868 21646 21870 21698
rect 21870 21646 21922 21698
rect 21922 21646 21924 21698
rect 21868 21644 21924 21646
rect 21644 21532 21700 21588
rect 20972 21474 21028 21476
rect 20972 21422 20974 21474
rect 20974 21422 21026 21474
rect 21026 21422 21028 21474
rect 20972 21420 21028 21422
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19516 18844 19572 18900
rect 19292 17948 19348 18004
rect 19180 17554 19236 17556
rect 19180 17502 19182 17554
rect 19182 17502 19234 17554
rect 19234 17502 19236 17554
rect 19180 17500 19236 17502
rect 19068 17388 19124 17444
rect 19404 17836 19460 17892
rect 19516 18620 19572 18676
rect 21532 18956 21588 19012
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20972 18562 21028 18564
rect 20972 18510 20974 18562
rect 20974 18510 21026 18562
rect 21026 18510 21028 18562
rect 20972 18508 21028 18510
rect 21868 20690 21924 20692
rect 21868 20638 21870 20690
rect 21870 20638 21922 20690
rect 21922 20638 21924 20690
rect 21868 20636 21924 20638
rect 22652 24946 22708 24948
rect 22652 24894 22654 24946
rect 22654 24894 22706 24946
rect 22706 24894 22708 24946
rect 22652 24892 22708 24894
rect 27468 27186 27524 27188
rect 27468 27134 27470 27186
rect 27470 27134 27522 27186
rect 27522 27134 27524 27186
rect 27468 27132 27524 27134
rect 27916 27132 27972 27188
rect 37660 27074 37716 27076
rect 37660 27022 37662 27074
rect 37662 27022 37714 27074
rect 37714 27022 37716 27074
rect 37660 27020 37716 27022
rect 28140 26962 28196 26964
rect 28140 26910 28142 26962
rect 28142 26910 28194 26962
rect 28194 26910 28196 26962
rect 28140 26908 28196 26910
rect 37884 26908 37940 26964
rect 23884 24892 23940 24948
rect 23436 24780 23492 24836
rect 23100 23714 23156 23716
rect 23100 23662 23102 23714
rect 23102 23662 23154 23714
rect 23154 23662 23156 23714
rect 23100 23660 23156 23662
rect 22764 22258 22820 22260
rect 22764 22206 22766 22258
rect 22766 22206 22818 22258
rect 22818 22206 22820 22258
rect 22764 22204 22820 22206
rect 22540 22092 22596 22148
rect 22428 21420 22484 21476
rect 22540 20972 22596 21028
rect 22876 21196 22932 21252
rect 21756 18508 21812 18564
rect 19740 17948 19796 18004
rect 21644 18396 21700 18452
rect 20636 17778 20692 17780
rect 20636 17726 20638 17778
rect 20638 17726 20690 17778
rect 20690 17726 20692 17778
rect 20636 17724 20692 17726
rect 19740 17666 19796 17668
rect 19740 17614 19742 17666
rect 19742 17614 19794 17666
rect 19794 17614 19796 17666
rect 19740 17612 19796 17614
rect 21532 17778 21588 17780
rect 21532 17726 21534 17778
rect 21534 17726 21586 17778
rect 21586 17726 21588 17778
rect 21532 17724 21588 17726
rect 22988 20748 23044 20804
rect 22764 18508 22820 18564
rect 21868 17778 21924 17780
rect 21868 17726 21870 17778
rect 21870 17726 21922 17778
rect 21922 17726 21924 17778
rect 21868 17724 21924 17726
rect 22316 17666 22372 17668
rect 22316 17614 22318 17666
rect 22318 17614 22370 17666
rect 22370 17614 22372 17666
rect 22316 17612 22372 17614
rect 20748 17442 20804 17444
rect 20748 17390 20750 17442
rect 20750 17390 20802 17442
rect 20802 17390 20804 17442
rect 20748 17388 20804 17390
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19628 17052 19684 17108
rect 18508 15426 18564 15428
rect 18508 15374 18510 15426
rect 18510 15374 18562 15426
rect 18562 15374 18564 15426
rect 18508 15372 18564 15374
rect 18620 15202 18676 15204
rect 18620 15150 18622 15202
rect 18622 15150 18674 15202
rect 18674 15150 18676 15202
rect 18620 15148 18676 15150
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 18844 16658 18900 16660
rect 18844 16606 18846 16658
rect 18846 16606 18898 16658
rect 18898 16606 18900 16658
rect 18844 16604 18900 16606
rect 18956 16098 19012 16100
rect 18956 16046 18958 16098
rect 18958 16046 19010 16098
rect 19010 16046 19012 16098
rect 18956 16044 19012 16046
rect 18844 15820 18900 15876
rect 18508 13580 18564 13636
rect 18956 14476 19012 14532
rect 19292 15484 19348 15540
rect 19516 16828 19572 16884
rect 22204 17500 22260 17556
rect 21644 16604 21700 16660
rect 21756 16044 21812 16100
rect 20412 15874 20468 15876
rect 20412 15822 20414 15874
rect 20414 15822 20466 15874
rect 20466 15822 20468 15874
rect 20412 15820 20468 15822
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19628 15484 19684 15540
rect 19516 15148 19572 15204
rect 19852 15260 19908 15316
rect 21868 15484 21924 15540
rect 21420 15426 21476 15428
rect 21420 15374 21422 15426
rect 21422 15374 21474 15426
rect 21474 15374 21476 15426
rect 21420 15372 21476 15374
rect 19404 14476 19460 14532
rect 21196 15148 21252 15204
rect 19740 14306 19796 14308
rect 19740 14254 19742 14306
rect 19742 14254 19794 14306
rect 19794 14254 19796 14306
rect 19740 14252 19796 14254
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20412 14252 20468 14308
rect 20188 13634 20244 13636
rect 20188 13582 20190 13634
rect 20190 13582 20242 13634
rect 20242 13582 20244 13634
rect 20188 13580 20244 13582
rect 20076 13468 20132 13524
rect 20300 12908 20356 12964
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 17724 5180 17780 5236
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 18732 5234 18788 5236
rect 18732 5182 18734 5234
rect 18734 5182 18786 5234
rect 18786 5182 18788 5234
rect 18732 5180 18788 5182
rect 21532 14476 21588 14532
rect 21868 15260 21924 15316
rect 22092 15874 22148 15876
rect 22092 15822 22094 15874
rect 22094 15822 22146 15874
rect 22146 15822 22148 15874
rect 22092 15820 22148 15822
rect 22652 18450 22708 18452
rect 22652 18398 22654 18450
rect 22654 18398 22706 18450
rect 22706 18398 22708 18450
rect 22652 18396 22708 18398
rect 22540 17388 22596 17444
rect 25452 25452 25508 25508
rect 25228 24892 25284 24948
rect 24332 24780 24388 24836
rect 25788 24722 25844 24724
rect 25788 24670 25790 24722
rect 25790 24670 25842 24722
rect 25842 24670 25844 24722
rect 25788 24668 25844 24670
rect 23324 21756 23380 21812
rect 23212 21698 23268 21700
rect 23212 21646 23214 21698
rect 23214 21646 23266 21698
rect 23266 21646 23268 21698
rect 23212 21644 23268 21646
rect 23996 21586 24052 21588
rect 23996 21534 23998 21586
rect 23998 21534 24050 21586
rect 24050 21534 24052 21586
rect 23996 21532 24052 21534
rect 24332 23212 24388 23268
rect 24780 23548 24836 23604
rect 24108 21196 24164 21252
rect 24668 23436 24724 23492
rect 25228 23714 25284 23716
rect 25228 23662 25230 23714
rect 25230 23662 25282 23714
rect 25282 23662 25284 23714
rect 25228 23660 25284 23662
rect 25228 23436 25284 23492
rect 39900 26796 39956 26852
rect 40012 26236 40068 26292
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 26012 23714 26068 23716
rect 26012 23662 26014 23714
rect 26014 23662 26066 23714
rect 26066 23662 26068 23714
rect 26012 23660 26068 23662
rect 26124 23548 26180 23604
rect 26012 23266 26068 23268
rect 26012 23214 26014 23266
rect 26014 23214 26066 23266
rect 26066 23214 26068 23266
rect 26012 23212 26068 23214
rect 25004 22316 25060 22372
rect 28140 23884 28196 23940
rect 37660 23938 37716 23940
rect 37660 23886 37662 23938
rect 37662 23886 37714 23938
rect 37714 23886 37716 23938
rect 37660 23884 37716 23886
rect 28140 23548 28196 23604
rect 40012 23548 40068 23604
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 27020 22428 27076 22484
rect 27580 22482 27636 22484
rect 27580 22430 27582 22482
rect 27582 22430 27634 22482
rect 27634 22430 27636 22482
rect 27580 22428 27636 22430
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 37660 22428 37716 22484
rect 37324 21586 37380 21588
rect 37324 21534 37326 21586
rect 37326 21534 37378 21586
rect 37378 21534 37380 21586
rect 37324 21532 37380 21534
rect 37772 21586 37828 21588
rect 37772 21534 37774 21586
rect 37774 21534 37826 21586
rect 37826 21534 37828 21586
rect 37772 21532 37828 21534
rect 26572 21420 26628 21476
rect 27692 21420 27748 21476
rect 26348 20802 26404 20804
rect 26348 20750 26350 20802
rect 26350 20750 26402 20802
rect 26402 20750 26404 20802
rect 26348 20748 26404 20750
rect 24220 20636 24276 20692
rect 25900 20690 25956 20692
rect 25900 20638 25902 20690
rect 25902 20638 25954 20690
rect 25954 20638 25956 20690
rect 25900 20636 25956 20638
rect 26796 20690 26852 20692
rect 26796 20638 26798 20690
rect 26798 20638 26850 20690
rect 26850 20638 26852 20690
rect 26796 20636 26852 20638
rect 25676 20578 25732 20580
rect 25676 20526 25678 20578
rect 25678 20526 25730 20578
rect 25730 20526 25732 20578
rect 25676 20524 25732 20526
rect 22428 17052 22484 17108
rect 22988 17052 23044 17108
rect 24220 18956 24276 19012
rect 23212 17554 23268 17556
rect 23212 17502 23214 17554
rect 23214 17502 23266 17554
rect 23266 17502 23268 17554
rect 23212 17500 23268 17502
rect 23772 17500 23828 17556
rect 22876 16156 22932 16212
rect 22764 16098 22820 16100
rect 22764 16046 22766 16098
rect 22766 16046 22818 16098
rect 22818 16046 22820 16098
rect 22764 16044 22820 16046
rect 25004 19010 25060 19012
rect 25004 18958 25006 19010
rect 25006 18958 25058 19010
rect 25058 18958 25060 19010
rect 25004 18956 25060 18958
rect 25452 18956 25508 19012
rect 27356 20802 27412 20804
rect 27356 20750 27358 20802
rect 27358 20750 27410 20802
rect 27410 20750 27412 20802
rect 27356 20748 27412 20750
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 39900 20860 39956 20916
rect 37660 20802 37716 20804
rect 37660 20750 37662 20802
rect 37662 20750 37714 20802
rect 37714 20750 37716 20802
rect 37660 20748 37716 20750
rect 27580 20578 27636 20580
rect 27580 20526 27582 20578
rect 27582 20526 27634 20578
rect 27634 20526 27636 20578
rect 27580 20524 27636 20526
rect 27692 20412 27748 20468
rect 28364 20524 28420 20580
rect 27244 19740 27300 19796
rect 28252 20076 28308 20132
rect 28700 20412 28756 20468
rect 40012 20188 40068 20244
rect 28812 20130 28868 20132
rect 28812 20078 28814 20130
rect 28814 20078 28866 20130
rect 28866 20078 28868 20130
rect 28812 20076 28868 20078
rect 37660 20018 37716 20020
rect 37660 19966 37662 20018
rect 37662 19966 37714 20018
rect 37714 19966 37716 20018
rect 37660 19964 37716 19966
rect 28812 19794 28868 19796
rect 28812 19742 28814 19794
rect 28814 19742 28866 19794
rect 28866 19742 28868 19794
rect 28812 19740 28868 19742
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 40012 19516 40068 19572
rect 25900 18396 25956 18452
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 26012 17778 26068 17780
rect 26012 17726 26014 17778
rect 26014 17726 26066 17778
rect 26066 17726 26068 17778
rect 26012 17724 26068 17726
rect 26124 17666 26180 17668
rect 26124 17614 26126 17666
rect 26126 17614 26178 17666
rect 26178 17614 26180 17666
rect 26124 17612 26180 17614
rect 26908 17612 26964 17668
rect 24780 16210 24836 16212
rect 24780 16158 24782 16210
rect 24782 16158 24834 16210
rect 24834 16158 24836 16210
rect 24780 16156 24836 16158
rect 37660 17666 37716 17668
rect 37660 17614 37662 17666
rect 37662 17614 37714 17666
rect 37714 17614 37716 17666
rect 37660 17612 37716 17614
rect 40012 17500 40068 17556
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 22316 15820 22372 15876
rect 21980 14588 22036 14644
rect 22652 15484 22708 15540
rect 22540 15426 22596 15428
rect 22540 15374 22542 15426
rect 22542 15374 22594 15426
rect 22594 15374 22596 15426
rect 22540 15372 22596 15374
rect 22428 15314 22484 15316
rect 22428 15262 22430 15314
rect 22430 15262 22482 15314
rect 22482 15262 22484 15314
rect 22428 15260 22484 15262
rect 23548 14642 23604 14644
rect 23548 14590 23550 14642
rect 23550 14590 23602 14642
rect 23602 14590 23604 14642
rect 23548 14588 23604 14590
rect 22764 14530 22820 14532
rect 22764 14478 22766 14530
rect 22766 14478 22818 14530
rect 22818 14478 22820 14530
rect 22764 14476 22820 14478
rect 21868 13356 21924 13412
rect 21532 12962 21588 12964
rect 21532 12910 21534 12962
rect 21534 12910 21586 12962
rect 21586 12910 21588 12962
rect 21532 12908 21588 12910
rect 25228 15426 25284 15428
rect 25228 15374 25230 15426
rect 25230 15374 25282 15426
rect 25282 15374 25284 15426
rect 25228 15372 25284 15374
rect 23660 14252 23716 14308
rect 24556 14252 24612 14308
rect 22204 13580 22260 13636
rect 24108 13634 24164 13636
rect 24108 13582 24110 13634
rect 24110 13582 24162 13634
rect 24162 13582 24164 13634
rect 24108 13580 24164 13582
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20188 4060 20244 4116
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 20860 3612 20916 3668
rect 23548 5180 23604 5236
rect 21420 4114 21476 4116
rect 21420 4062 21422 4114
rect 21422 4062 21474 4114
rect 21474 4062 21476 4114
rect 21420 4060 21476 4062
rect 22092 3666 22148 3668
rect 22092 3614 22094 3666
rect 22094 3614 22146 3666
rect 22146 3614 22148 3666
rect 22092 3612 22148 3614
rect 22876 3612 22932 3668
rect 24780 5234 24836 5236
rect 24780 5182 24782 5234
rect 24782 5182 24834 5234
rect 24834 5182 24836 5234
rect 24780 5180 24836 5182
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
rect 25004 3554 25060 3556
rect 25004 3502 25006 3554
rect 25006 3502 25058 3554
rect 25058 3502 25060 3554
rect 25004 3500 25060 3502
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 25676 3500 25732 3556
rect 25788 4060 25844 4116
rect 26796 4114 26852 4116
rect 26796 4062 26798 4114
rect 26798 4062 26850 4114
rect 26850 4062 26852 4114
rect 26796 4060 26852 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 17490 38220 17500 38276
rect 17556 38220 18620 38276
rect 18676 38220 18686 38276
rect 22866 38220 22876 38276
rect 22932 38220 25564 38276
rect 25620 38220 25630 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 16818 37436 16828 37492
rect 16884 37436 18396 37492
rect 18452 37436 18462 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 18274 27692 18284 27748
rect 18340 27692 20412 27748
rect 20468 27692 20478 27748
rect 22754 27692 22764 27748
rect 22820 27692 23548 27748
rect 23604 27692 24556 27748
rect 24612 27692 24622 27748
rect 0 27636 800 27664
rect 0 27580 4172 27636
rect 4228 27580 4238 27636
rect 15138 27580 15148 27636
rect 15204 27580 17388 27636
rect 17444 27580 17454 27636
rect 0 27552 800 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 26898 27132 26908 27188
rect 26964 27132 27468 27188
rect 27524 27132 27916 27188
rect 27972 27132 31948 27188
rect 31892 27076 31948 27132
rect 4274 27020 4284 27076
rect 4340 27020 12124 27076
rect 12180 27020 12190 27076
rect 20402 27020 20412 27076
rect 20468 27020 21532 27076
rect 21588 27020 21598 27076
rect 22082 27020 22092 27076
rect 22148 27020 22764 27076
rect 22820 27020 22830 27076
rect 31892 27020 37660 27076
rect 37716 27020 37726 27076
rect 41200 26964 42000 26992
rect 16818 26908 16828 26964
rect 16884 26908 17612 26964
rect 17668 26908 18284 26964
rect 18340 26908 18350 26964
rect 21634 26908 21644 26964
rect 21700 26908 24220 26964
rect 24276 26908 24668 26964
rect 24724 26908 24734 26964
rect 28130 26908 28140 26964
rect 28196 26908 37884 26964
rect 37940 26908 37950 26964
rect 39900 26908 42000 26964
rect 39900 26852 39956 26908
rect 41200 26880 42000 26908
rect 17154 26796 17164 26852
rect 17220 26796 17500 26852
rect 17556 26796 20524 26852
rect 20580 26796 20590 26852
rect 39890 26796 39900 26852
rect 39956 26796 39966 26852
rect 20626 26684 20636 26740
rect 20692 26684 22876 26740
rect 22932 26684 22942 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 18722 26460 18732 26516
rect 18788 26460 19628 26516
rect 19684 26460 21308 26516
rect 21364 26460 22540 26516
rect 22596 26460 22606 26516
rect 0 26292 800 26320
rect 41200 26292 42000 26320
rect 0 26236 1932 26292
rect 1988 26236 1998 26292
rect 4274 26236 4284 26292
rect 4340 26236 12124 26292
rect 12180 26236 12190 26292
rect 13122 26236 13132 26292
rect 13188 26236 13804 26292
rect 13860 26236 13870 26292
rect 16146 26236 16156 26292
rect 16212 26236 18956 26292
rect 19012 26236 19022 26292
rect 40002 26236 40012 26292
rect 40068 26236 42000 26292
rect 0 26208 800 26236
rect 41200 26208 42000 26236
rect 14466 26124 14476 26180
rect 14532 26124 16044 26180
rect 16100 26124 16110 26180
rect 16594 26124 16604 26180
rect 16660 26124 17052 26180
rect 17108 26124 17118 26180
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 11666 25676 11676 25732
rect 11732 25676 12348 25732
rect 12404 25676 12414 25732
rect 0 25620 800 25648
rect 0 25564 1932 25620
rect 1988 25564 1998 25620
rect 16594 25564 16604 25620
rect 16660 25564 16940 25620
rect 16996 25564 17006 25620
rect 17276 25564 21532 25620
rect 21588 25564 21598 25620
rect 0 25536 800 25564
rect 17276 25508 17332 25564
rect 4274 25452 4284 25508
rect 4340 25452 10220 25508
rect 10276 25452 12348 25508
rect 12404 25452 12414 25508
rect 15092 25452 17332 25508
rect 17490 25452 17500 25508
rect 17556 25452 18844 25508
rect 18900 25452 18910 25508
rect 22418 25452 22428 25508
rect 22484 25452 25452 25508
rect 25508 25452 25518 25508
rect 15092 25396 15148 25452
rect 11666 25340 11676 25396
rect 11732 25340 15148 25396
rect 17266 25340 17276 25396
rect 17332 25340 18284 25396
rect 18340 25340 19292 25396
rect 19348 25340 19358 25396
rect 15922 25228 15932 25284
rect 15988 25228 17388 25284
rect 17444 25228 17454 25284
rect 21746 25228 21756 25284
rect 21812 25228 22372 25284
rect 13794 25116 13804 25172
rect 13860 25116 14476 25172
rect 14532 25116 16268 25172
rect 16324 25116 16828 25172
rect 16884 25116 16894 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 22316 25060 22372 25228
rect 22306 25004 22316 25060
rect 22372 25004 22382 25060
rect 0 24948 800 24976
rect 0 24892 2044 24948
rect 2100 24892 2110 24948
rect 18946 24892 18956 24948
rect 19012 24892 22652 24948
rect 22708 24892 23884 24948
rect 23940 24892 25228 24948
rect 25284 24892 25294 24948
rect 0 24864 800 24892
rect 18386 24780 18396 24836
rect 18452 24780 19852 24836
rect 19908 24780 19918 24836
rect 20626 24780 20636 24836
rect 20692 24780 21868 24836
rect 21924 24780 23436 24836
rect 23492 24780 24332 24836
rect 24388 24780 24398 24836
rect 19730 24668 19740 24724
rect 19796 24668 25788 24724
rect 25844 24668 25854 24724
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 17602 24108 17612 24164
rect 17668 24108 18172 24164
rect 18228 24108 19068 24164
rect 19124 24108 19134 24164
rect 19842 23996 19852 24052
rect 19908 23996 20524 24052
rect 20580 23996 20590 24052
rect 16258 23884 16268 23940
rect 16324 23884 17500 23940
rect 17556 23884 18732 23940
rect 18788 23884 18798 23940
rect 19618 23884 19628 23940
rect 19684 23884 20076 23940
rect 20132 23884 21980 23940
rect 22036 23884 22046 23940
rect 28130 23884 28140 23940
rect 28196 23884 37660 23940
rect 37716 23884 37726 23940
rect 4274 23772 4284 23828
rect 4340 23772 13468 23828
rect 13524 23772 13534 23828
rect 18610 23772 18620 23828
rect 18676 23772 19180 23828
rect 19236 23772 20188 23828
rect 20244 23772 20254 23828
rect 0 23604 800 23632
rect 13468 23604 13524 23772
rect 17602 23660 17612 23716
rect 17668 23660 18396 23716
rect 18452 23660 18462 23716
rect 18722 23660 18732 23716
rect 18788 23660 21588 23716
rect 22082 23660 22092 23716
rect 22148 23660 23100 23716
rect 23156 23660 25228 23716
rect 25284 23660 25294 23716
rect 26002 23660 26012 23716
rect 26068 23660 26908 23716
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 12674 23548 12684 23604
rect 12740 23548 13412 23604
rect 13468 23548 15484 23604
rect 15540 23548 15550 23604
rect 16930 23548 16940 23604
rect 16996 23548 19628 23604
rect 19684 23548 19694 23604
rect 0 23520 800 23548
rect 13356 23492 13412 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 21532 23492 21588 23660
rect 26852 23604 26908 23660
rect 41200 23604 42000 23632
rect 24770 23548 24780 23604
rect 24836 23548 26124 23604
rect 26180 23548 26190 23604
rect 26852 23548 28140 23604
rect 28196 23548 28206 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 41200 23520 42000 23548
rect 13356 23436 13468 23492
rect 13524 23436 14252 23492
rect 14308 23436 15148 23492
rect 21532 23436 24668 23492
rect 24724 23436 25228 23492
rect 25284 23436 25294 23492
rect 15092 23380 15148 23436
rect 15092 23324 15372 23380
rect 15428 23324 16716 23380
rect 16772 23324 16782 23380
rect 8372 23212 11004 23268
rect 11060 23212 14364 23268
rect 14420 23212 14430 23268
rect 24322 23212 24332 23268
rect 24388 23212 26012 23268
rect 26068 23212 26078 23268
rect 8372 23156 8428 23212
rect 4274 23100 4284 23156
rect 4340 23100 8428 23156
rect 14802 22988 14812 23044
rect 14868 22988 15596 23044
rect 15652 22988 15662 23044
rect 0 22932 800 22960
rect 41200 22932 42000 22960
rect 0 22876 1932 22932
rect 1988 22876 1998 22932
rect 14354 22876 14364 22932
rect 14420 22876 15260 22932
rect 15316 22876 15326 22932
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 0 22848 800 22876
rect 41200 22848 42000 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 13122 22540 13132 22596
rect 13188 22540 15484 22596
rect 15540 22540 15550 22596
rect 17938 22428 17948 22484
rect 18004 22428 18620 22484
rect 18676 22428 18686 22484
rect 27010 22428 27020 22484
rect 27076 22428 27580 22484
rect 27636 22428 37660 22484
rect 37716 22428 37726 22484
rect 16146 22316 16156 22372
rect 16212 22316 18508 22372
rect 18564 22316 18574 22372
rect 19618 22316 19628 22372
rect 19684 22316 25004 22372
rect 25060 22316 25070 22372
rect 19628 22260 19684 22316
rect 15810 22204 15820 22260
rect 15876 22204 17724 22260
rect 17780 22204 19684 22260
rect 21410 22204 21420 22260
rect 21476 22204 22764 22260
rect 22820 22204 22830 22260
rect 15698 22092 15708 22148
rect 15764 22092 21868 22148
rect 21924 22092 22540 22148
rect 22596 22092 22606 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 12898 21756 12908 21812
rect 12964 21756 13916 21812
rect 13972 21756 13982 21812
rect 15586 21756 15596 21812
rect 15652 21756 18060 21812
rect 18116 21756 18126 21812
rect 20514 21756 20524 21812
rect 20580 21756 23324 21812
rect 23380 21756 23390 21812
rect 8372 21644 9996 21700
rect 10052 21644 13356 21700
rect 13412 21644 13422 21700
rect 17490 21644 17500 21700
rect 17556 21644 21868 21700
rect 21924 21644 23212 21700
rect 23268 21644 23278 21700
rect 0 21588 800 21616
rect 0 21532 1932 21588
rect 1988 21532 1998 21588
rect 0 21504 800 21532
rect 8372 21476 8428 21644
rect 21634 21532 21644 21588
rect 21700 21532 23996 21588
rect 24052 21532 37324 21588
rect 37380 21532 37772 21588
rect 37828 21532 37838 21588
rect 4274 21420 4284 21476
rect 4340 21420 8428 21476
rect 20962 21420 20972 21476
rect 21028 21420 22428 21476
rect 22484 21420 22494 21476
rect 26562 21420 26572 21476
rect 26628 21420 27692 21476
rect 27748 21420 27758 21476
rect 17388 21308 18844 21364
rect 18900 21308 18910 21364
rect 17388 21252 17444 21308
rect 12450 21196 12460 21252
rect 12516 21196 17388 21252
rect 17444 21196 17454 21252
rect 18946 21196 18956 21252
rect 19012 21196 22876 21252
rect 22932 21196 24108 21252
rect 24164 21196 24174 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 18050 21084 18060 21140
rect 18116 21084 18732 21140
rect 18788 21084 18798 21140
rect 18386 20972 18396 21028
rect 18452 20972 19628 21028
rect 19684 20972 22540 21028
rect 22596 20972 22606 21028
rect 41200 20916 42000 20944
rect 18610 20860 18620 20916
rect 18676 20860 20076 20916
rect 20132 20860 20142 20916
rect 39890 20860 39900 20916
rect 39956 20860 42000 20916
rect 41200 20832 42000 20860
rect 15138 20748 15148 20804
rect 15204 20748 15932 20804
rect 15988 20748 16268 20804
rect 16324 20748 16828 20804
rect 16884 20748 16894 20804
rect 22978 20748 22988 20804
rect 23044 20748 23054 20804
rect 26338 20748 26348 20804
rect 26404 20748 27356 20804
rect 27412 20748 27422 20804
rect 31892 20748 37660 20804
rect 37716 20748 37726 20804
rect 22988 20692 23044 20748
rect 21858 20636 21868 20692
rect 21924 20636 24220 20692
rect 24276 20636 25900 20692
rect 25956 20636 26796 20692
rect 26852 20636 26862 20692
rect 31892 20580 31948 20748
rect 18050 20524 18060 20580
rect 18116 20524 18956 20580
rect 19012 20524 19022 20580
rect 19282 20524 19292 20580
rect 19348 20524 25676 20580
rect 25732 20524 25742 20580
rect 27570 20524 27580 20580
rect 27636 20524 28364 20580
rect 28420 20524 31948 20580
rect 27682 20412 27692 20468
rect 27748 20412 28700 20468
rect 28756 20412 28766 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 16146 20300 16156 20356
rect 16212 20300 17388 20356
rect 17444 20300 18396 20356
rect 18452 20300 18462 20356
rect 41200 20244 42000 20272
rect 16930 20188 16940 20244
rect 16996 20188 17500 20244
rect 17556 20188 18116 20244
rect 40002 20188 40012 20244
rect 40068 20188 42000 20244
rect 18060 20132 18116 20188
rect 41200 20160 42000 20188
rect 13010 20076 13020 20132
rect 13076 20076 15484 20132
rect 15540 20076 15550 20132
rect 15810 20076 15820 20132
rect 15876 20076 17276 20132
rect 17332 20076 17724 20132
rect 17780 20076 17790 20132
rect 18060 20076 18284 20132
rect 18340 20076 18350 20132
rect 28242 20076 28252 20132
rect 28308 20076 28812 20132
rect 28868 20076 31948 20132
rect 31892 20020 31948 20076
rect 4162 19964 4172 20020
rect 4228 19964 18732 20020
rect 18788 19964 18798 20020
rect 31892 19964 37660 20020
rect 37716 19964 37726 20020
rect 16594 19852 16604 19908
rect 16660 19852 19180 19908
rect 19236 19852 19246 19908
rect 27234 19740 27244 19796
rect 27300 19740 28812 19796
rect 28868 19740 28878 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 41200 19488 42000 19516
rect 15474 19404 15484 19460
rect 15540 19404 15820 19460
rect 15876 19404 17836 19460
rect 17892 19404 17902 19460
rect 15922 19180 15932 19236
rect 15988 19180 16604 19236
rect 16660 19180 16670 19236
rect 15372 19068 18844 19124
rect 18900 19068 18910 19124
rect 15372 19012 15428 19068
rect 12226 18956 12236 19012
rect 12292 18956 14028 19012
rect 14084 18956 15372 19012
rect 15428 18956 15438 19012
rect 16818 18956 16828 19012
rect 16884 18956 21532 19012
rect 21588 18956 21598 19012
rect 24210 18956 24220 19012
rect 24276 18956 25004 19012
rect 25060 18956 25452 19012
rect 25508 18956 25518 19012
rect 15026 18844 15036 18900
rect 15092 18844 15708 18900
rect 15764 18844 17164 18900
rect 17220 18844 18060 18900
rect 18116 18844 19516 18900
rect 19572 18844 19582 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 19170 18620 19180 18676
rect 19236 18620 19516 18676
rect 19572 18620 19582 18676
rect 17714 18508 17724 18564
rect 17780 18508 20972 18564
rect 21028 18508 21038 18564
rect 21746 18508 21756 18564
rect 21812 18508 22764 18564
rect 22820 18508 22830 18564
rect 15922 18396 15932 18452
rect 15988 18396 21644 18452
rect 21700 18396 22652 18452
rect 22708 18396 25900 18452
rect 25956 18396 25966 18452
rect 13794 18284 13804 18340
rect 13860 18284 15820 18340
rect 15876 18284 15886 18340
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 19282 17948 19292 18004
rect 19348 17948 19740 18004
rect 19796 17948 19806 18004
rect 19366 17836 19404 17892
rect 19460 17836 19470 17892
rect 20626 17724 20636 17780
rect 20692 17724 21532 17780
rect 21588 17724 21598 17780
rect 21858 17724 21868 17780
rect 21924 17724 26012 17780
rect 26068 17724 26078 17780
rect 17714 17612 17724 17668
rect 17780 17612 19740 17668
rect 19796 17612 22316 17668
rect 22372 17612 22382 17668
rect 26114 17612 26124 17668
rect 26180 17612 26908 17668
rect 26964 17612 37660 17668
rect 37716 17612 37726 17668
rect 41200 17556 42000 17584
rect 19170 17500 19180 17556
rect 19236 17500 22204 17556
rect 22260 17500 23212 17556
rect 23268 17500 23772 17556
rect 23828 17500 23838 17556
rect 40002 17500 40012 17556
rect 40068 17500 42000 17556
rect 41200 17472 42000 17500
rect 18498 17388 18508 17444
rect 18564 17388 19068 17444
rect 19124 17388 19134 17444
rect 20738 17388 20748 17444
rect 20804 17388 22540 17444
rect 22596 17388 22606 17444
rect 14690 17276 14700 17332
rect 14756 17276 18732 17332
rect 18788 17276 18798 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 19618 17052 19628 17108
rect 19684 17052 22428 17108
rect 22484 17052 22988 17108
rect 23044 17052 23054 17108
rect 14018 16828 14028 16884
rect 14084 16828 16044 16884
rect 16100 16828 17500 16884
rect 17556 16828 19516 16884
rect 19572 16828 19582 16884
rect 18834 16604 18844 16660
rect 18900 16604 21644 16660
rect 21700 16604 21710 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 22866 16156 22876 16212
rect 22932 16156 24780 16212
rect 24836 16156 24846 16212
rect 18946 16044 18956 16100
rect 19012 16044 19404 16100
rect 19460 16044 19470 16100
rect 21746 16044 21756 16100
rect 21812 16044 22764 16100
rect 22820 16044 22830 16100
rect 22316 15876 22372 16044
rect 16818 15820 16828 15876
rect 16884 15820 17724 15876
rect 17780 15820 17790 15876
rect 18834 15820 18844 15876
rect 18900 15820 20412 15876
rect 20468 15820 22092 15876
rect 22148 15820 22158 15876
rect 22306 15820 22316 15876
rect 22372 15820 22382 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 17602 15484 17612 15540
rect 17668 15484 19292 15540
rect 19348 15484 19628 15540
rect 19684 15484 19694 15540
rect 21858 15484 21868 15540
rect 21924 15484 22652 15540
rect 22708 15484 22718 15540
rect 18498 15372 18508 15428
rect 18564 15372 21420 15428
rect 21476 15372 21486 15428
rect 22530 15372 22540 15428
rect 22596 15372 25228 15428
rect 25284 15372 25294 15428
rect 14690 15260 14700 15316
rect 14756 15260 17724 15316
rect 17780 15260 17790 15316
rect 19842 15260 19852 15316
rect 19908 15260 21868 15316
rect 21924 15260 22428 15316
rect 22484 15260 22494 15316
rect 16706 15148 16716 15204
rect 16772 15148 18620 15204
rect 18676 15148 18686 15204
rect 19506 15148 19516 15204
rect 19572 15148 21196 15204
rect 21252 15148 21262 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 21970 14588 21980 14644
rect 22036 14588 23548 14644
rect 23604 14588 23614 14644
rect 18946 14476 18956 14532
rect 19012 14476 19404 14532
rect 19460 14476 19470 14532
rect 21522 14476 21532 14532
rect 21588 14476 22764 14532
rect 22820 14476 23548 14532
rect 23492 14308 23548 14476
rect 19730 14252 19740 14308
rect 19796 14252 20412 14308
rect 20468 14252 20478 14308
rect 23492 14252 23660 14308
rect 23716 14252 24556 14308
rect 24612 14252 24622 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 18498 13580 18508 13636
rect 18564 13580 20188 13636
rect 20244 13580 20254 13636
rect 22194 13580 22204 13636
rect 22260 13580 24108 13636
rect 24164 13580 24174 13636
rect 20066 13468 20076 13524
rect 20132 13468 20916 13524
rect 20860 13412 20916 13468
rect 20860 13356 21868 13412
rect 21924 13356 21934 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 20290 12908 20300 12964
rect 20356 12908 21532 12964
rect 21588 12908 21598 12964
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 17714 5180 17724 5236
rect 17780 5180 18732 5236
rect 18788 5180 18798 5236
rect 23538 5180 23548 5236
rect 23604 5180 24780 5236
rect 24836 5180 24846 5236
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 20178 4060 20188 4116
rect 20244 4060 21420 4116
rect 21476 4060 21486 4116
rect 25778 4060 25788 4116
rect 25844 4060 26796 4116
rect 26852 4060 26862 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 20850 3612 20860 3668
rect 20916 3612 22092 3668
rect 22148 3612 22158 3668
rect 22866 3612 22876 3668
rect 22932 3612 25564 3668
rect 25620 3612 25630 3668
rect 24994 3500 25004 3556
rect 25060 3500 25676 3556
rect 25732 3500 25742 3556
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19404 17836 19460 17892
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19404 16044 19460 16100
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 19404 17892 19460 17902
rect 19404 16100 19460 17836
rect 19404 16034 19460 16044
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _092_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22736 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _093_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20384 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _094_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _095_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23632 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _096_
timestamp 1698175906
transform -1 0 20832 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _097_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _098_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18592 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _099_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18592 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18368 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _101_
timestamp 1698175906
transform 1 0 16128 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19040 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19936 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _104_
timestamp 1698175906
transform 1 0 20272 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _105_
timestamp 1698175906
transform 1 0 22064 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_
timestamp 1698175906
transform -1 0 21952 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17472 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _108_
timestamp 1698175906
transform 1 0 15456 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_
timestamp 1698175906
transform 1 0 19152 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1698175906
transform -1 0 23632 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _111_
timestamp 1698175906
transform 1 0 22064 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _112_
timestamp 1698175906
transform -1 0 20832 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_
timestamp 1698175906
transform -1 0 20720 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20720 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform 1 0 25648 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _116_
timestamp 1698175906
transform -1 0 26880 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698175906
transform 1 0 16352 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform 1 0 21392 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _120_
timestamp 1698175906
transform 1 0 25760 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24864 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _122_
timestamp 1698175906
transform -1 0 16128 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _123_
timestamp 1698175906
transform 1 0 17024 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _124_
timestamp 1698175906
transform 1 0 17584 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17024 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14000 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _128_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22288 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _129_
timestamp 1698175906
transform -1 0 22624 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _130_
timestamp 1698175906
transform -1 0 22064 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _131_
timestamp 1698175906
transform 1 0 18144 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _132_
timestamp 1698175906
transform -1 0 19152 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _133_
timestamp 1698175906
transform -1 0 19936 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _134_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18144 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _135_
timestamp 1698175906
transform -1 0 17248 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _136_
timestamp 1698175906
transform -1 0 13664 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _137_
timestamp 1698175906
transform -1 0 12768 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _138_
timestamp 1698175906
transform -1 0 19376 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _139_
timestamp 1698175906
transform -1 0 20048 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _140_
timestamp 1698175906
transform 1 0 16464 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _141_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _142_
timestamp 1698175906
transform -1 0 17920 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _143_
timestamp 1698175906
transform -1 0 12880 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _144_
timestamp 1698175906
transform -1 0 11984 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform 1 0 15568 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _146_
timestamp 1698175906
transform 1 0 28560 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _147_
timestamp 1698175906
transform 1 0 26432 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_
timestamp 1698175906
transform -1 0 26992 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _149_
timestamp 1698175906
transform 1 0 24864 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _150_
timestamp 1698175906
transform -1 0 16128 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _151_
timestamp 1698175906
transform 1 0 14672 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _152_
timestamp 1698175906
transform 1 0 22512 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _153_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22288 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _154_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22288 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _155_
timestamp 1698175906
transform 1 0 23408 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _156_
timestamp 1698175906
transform -1 0 26320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _157_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22512 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _158_
timestamp 1698175906
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _159_
timestamp 1698175906
transform 1 0 22512 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _160_
timestamp 1698175906
transform -1 0 18480 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _161_
timestamp 1698175906
transform 1 0 18480 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _162_
timestamp 1698175906
transform -1 0 27888 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _163_
timestamp 1698175906
transform 1 0 25536 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _164_
timestamp 1698175906
transform -1 0 20944 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _165_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19600 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _166_
timestamp 1698175906
transform 1 0 18704 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _167_
timestamp 1698175906
transform 1 0 21728 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _168_
timestamp 1698175906
transform 1 0 21504 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _169_
timestamp 1698175906
transform 1 0 22288 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _170_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _171_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17584 0 -1 18816
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _172_
timestamp 1698175906
transform 1 0 18592 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _173_
timestamp 1698175906
transform 1 0 18368 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _174_
timestamp 1698175906
transform 1 0 19152 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _175_
timestamp 1698175906
transform -1 0 20496 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _176_
timestamp 1698175906
transform -1 0 18368 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform 1 0 14112 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _178_
timestamp 1698175906
transform 1 0 15232 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _179_
timestamp 1698175906
transform 1 0 22288 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _180_
timestamp 1698175906
transform -1 0 19152 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _181_
timestamp 1698175906
transform 1 0 21504 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _182_
timestamp 1698175906
transform -1 0 17696 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _183_
timestamp 1698175906
transform 1 0 15792 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _184_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13776 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _185_
timestamp 1698175906
transform 1 0 24416 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _186_
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _187_
timestamp 1698175906
transform 1 0 12096 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _188_
timestamp 1698175906
transform 1 0 11984 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _189_
timestamp 1698175906
transform 1 0 21280 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _190_
timestamp 1698175906
transform 1 0 17472 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _191_
timestamp 1698175906
transform -1 0 13104 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _192_
timestamp 1698175906
transform 1 0 14224 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _193_
timestamp 1698175906
transform -1 0 13328 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_
timestamp 1698175906
transform 1 0 25200 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1698175906
transform 1 0 24528 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _196_
timestamp 1698175906
transform -1 0 16576 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _197_
timestamp 1698175906
transform -1 0 24528 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _198_
timestamp 1698175906
transform 1 0 23856 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _199_
timestamp 1698175906
transform 1 0 13776 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _200_
timestamp 1698175906
transform 1 0 25312 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1698175906
transform 1 0 21056 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_
timestamp 1698175906
transform 1 0 20496 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform 1 0 15792 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform 1 0 17584 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform -1 0 14112 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform 1 0 22624 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform 1 0 13552 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _209_
timestamp 1698175906
transform -1 0 12656 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _210_
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _211_
timestamp 1698175906
transform 1 0 20160 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _212_
timestamp 1698175906
transform -1 0 12656 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _213_
timestamp 1698175906
transform 1 0 27664 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__153__C dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23968 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__CLK
timestamp 1698175906
transform 1 0 24192 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__CLK
timestamp 1698175906
transform 1 0 24640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__CLK
timestamp 1698175906
transform 1 0 15344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__CLK
timestamp 1698175906
transform 1 0 15456 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__CLK
timestamp 1698175906
transform 1 0 21056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__CLK
timestamp 1698175906
transform 1 0 20608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__CLK
timestamp 1698175906
transform 1 0 13888 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__CLK
timestamp 1698175906
transform -1 0 18368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__CLK
timestamp 1698175906
transform 1 0 13552 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__CLK
timestamp 1698175906
transform 1 0 24976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1698175906
transform 1 0 24304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__CLK
timestamp 1698175906
transform 1 0 17472 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__CLK
timestamp 1698175906
transform 1 0 18816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__CLK
timestamp 1698175906
transform 1 0 23632 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__CLK
timestamp 1698175906
transform -1 0 25312 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__CLK
timestamp 1698175906
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK
timestamp 1698175906
transform -1 0 20496 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1698175906
transform 1 0 19488 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform -1 0 21056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 14112 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 21504 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 18704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output5_I
timestamp 1698175906
transform 1 0 37296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18928 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 24752 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform -1 0 23968 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698175906
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698175906
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_195 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23184 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_203
timestamp 1698175906
transform 1 0 24080 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_216
timestamp 1698175906
transform 1 0 25536 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_243
timestamp 1698175906
transform 1 0 28560 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_275
timestamp 1698175906
transform 1 0 32144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698175906
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_139
timestamp 1698175906
transform 1 0 16912 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_143
timestamp 1698175906
transform 1 0 17360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_177 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_193
timestamp 1698175906
transform 1 0 22960 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_197
timestamp 1698175906
transform 1 0 23408 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_225
timestamp 1698175906
transform 1 0 26544 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_176
timestamp 1698175906
transform 1 0 21056 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698175906
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_139
timestamp 1698175906
transform 1 0 16912 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_143
timestamp 1698175906
transform 1 0 17360 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_179
timestamp 1698175906
transform 1 0 21392 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_188
timestamp 1698175906
transform 1 0 22400 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_220
timestamp 1698175906
transform 1 0 25984 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_236
timestamp 1698175906
transform 1 0 27776 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698175906
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_104
timestamp 1698175906
transform 1 0 12992 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_108
timestamp 1698175906
transform 1 0 13440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_110
timestamp 1698175906
transform 1 0 13664 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_146
timestamp 1698175906
transform 1 0 17696 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_171
timestamp 1698175906
transform 1 0 20496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_175
timestamp 1698175906
transform 1 0 20944 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_205
timestamp 1698175906
transform 1 0 24304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_127
timestamp 1698175906
transform 1 0 15568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_158
timestamp 1698175906
transform 1 0 19040 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_179
timestamp 1698175906
transform 1 0 21392 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_219
timestamp 1698175906
transform 1 0 25872 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_235
timestamp 1698175906
transform 1 0 27664 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698175906
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_160
timestamp 1698175906
transform 1 0 19264 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_164
timestamp 1698175906
transform 1 0 19712 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_172
timestamp 1698175906
transform 1 0 20608 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_176
timestamp 1698175906
transform 1 0 21056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_184
timestamp 1698175906
transform 1 0 21952 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_186
timestamp 1698175906
transform 1 0 22176 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_192
timestamp 1698175906
transform 1 0 22848 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698175906
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_218
timestamp 1698175906
transform 1 0 25760 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_250
timestamp 1698175906
transform 1 0 29344 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_266
timestamp 1698175906
transform 1 0 31136 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_274
timestamp 1698175906
transform 1 0 32032 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698175906
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_139
timestamp 1698175906
transform 1 0 16912 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_143
timestamp 1698175906
transform 1 0 17360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_152
timestamp 1698175906
transform 1 0 18368 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_154
timestamp 1698175906
transform 1 0 18592 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_161
timestamp 1698175906
transform 1 0 19376 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_179
timestamp 1698175906
transform 1 0 21392 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_195
timestamp 1698175906
transform 1 0 23184 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_230
timestamp 1698175906
transform 1 0 27104 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_238
timestamp 1698175906
transform 1 0 28000 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698175906
transform 1 0 28448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_104
timestamp 1698175906
transform 1 0 12992 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_108
timestamp 1698175906
transform 1 0 13440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_110
timestamp 1698175906
transform 1 0 13664 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_146
timestamp 1698175906
transform 1 0 17696 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_150
timestamp 1698175906
transform 1 0 18144 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_113
timestamp 1698175906
transform 1 0 14000 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_166
timestamp 1698175906
transform 1 0 19936 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_170
timestamp 1698175906
transform 1 0 20384 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_197
timestamp 1698175906
transform 1 0 23408 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_213
timestamp 1698175906
transform 1 0 25200 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_217
timestamp 1698175906
transform 1 0 25648 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_223
timestamp 1698175906
transform 1 0 26320 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_239
timestamp 1698175906
transform 1 0 28112 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698175906
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_88
timestamp 1698175906
transform 1 0 11200 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_92
timestamp 1698175906
transform 1 0 11648 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_94
timestamp 1698175906
transform 1 0 11872 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_124
timestamp 1698175906
transform 1 0 15232 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_144
timestamp 1698175906
transform 1 0 17472 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_185
timestamp 1698175906
transform 1 0 22064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_203
timestamp 1698175906
transform 1 0 24080 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698175906
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698175906
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 40320 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_123
timestamp 1698175906
transform 1 0 15120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_127
timestamp 1698175906
transform 1 0 15568 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_132
timestamp 1698175906
transform 1 0 16128 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_154
timestamp 1698175906
transform 1 0 18592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_172
timestamp 1698175906
transform 1 0 20608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698175906
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_207
timestamp 1698175906
transform 1 0 24528 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_242
timestamp 1698175906
transform 1 0 28448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_88
timestamp 1698175906
transform 1 0 11200 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_125
timestamp 1698175906
transform 1 0 15344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_138
timestamp 1698175906
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_144
timestamp 1698175906
transform 1 0 17472 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_153
timestamp 1698175906
transform 1 0 18480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_207
timestamp 1698175906
transform 1 0 24528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_248
timestamp 1698175906
transform 1 0 29120 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_69
timestamp 1698175906
transform 1 0 9072 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_85
timestamp 1698175906
transform 1 0 10864 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_93
timestamp 1698175906
transform 1 0 11760 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_102
timestamp 1698175906
transform 1 0 12768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698175906
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_123
timestamp 1698175906
transform 1 0 15120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_125
timestamp 1698175906
transform 1 0 15344 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_145
timestamp 1698175906
transform 1 0 17584 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_147
timestamp 1698175906
transform 1 0 17808 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_163
timestamp 1698175906
transform 1 0 19600 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_165
timestamp 1698175906
transform 1 0 19824 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698175906
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_199
timestamp 1698175906
transform 1 0 23632 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_207
timestamp 1698175906
transform 1 0 24528 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_211
timestamp 1698175906
transform 1 0 24976 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_214
timestamp 1698175906
transform 1 0 25312 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_237
timestamp 1698175906
transform 1 0 27888 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_110
timestamp 1698175906
transform 1 0 13664 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_114
timestamp 1698175906
transform 1 0 14112 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_130
timestamp 1698175906
transform 1 0 15904 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_138
timestamp 1698175906
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_152
timestamp 1698175906
transform 1 0 18368 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_166
timestamp 1698175906
transform 1 0 19936 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_168
timestamp 1698175906
transform 1 0 20160 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_200
timestamp 1698175906
transform 1 0 23744 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_204
timestamp 1698175906
transform 1 0 24192 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698175906
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698175906
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_318
timestamp 1698175906
transform 1 0 36960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_320
timestamp 1698175906
transform 1 0 37184 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 4480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_111
timestamp 1698175906
transform 1 0 13776 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_113
timestamp 1698175906
transform 1 0 14000 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_116
timestamp 1698175906
transform 1 0 14336 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_131
timestamp 1698175906
transform 1 0 16016 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_139
timestamp 1698175906
transform 1 0 16912 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_141
timestamp 1698175906
transform 1 0 17136 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_173
timestamp 1698175906
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_199
timestamp 1698175906
transform 1 0 23632 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_203
timestamp 1698175906
transform 1 0 24080 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_236
timestamp 1698175906
transform 1 0 27776 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 4480 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_80
timestamp 1698175906
transform 1 0 10304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_84
timestamp 1698175906
transform 1 0 10752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_132
timestamp 1698175906
transform 1 0 16128 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_150
timestamp 1698175906
transform 1 0 18144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_202
timestamp 1698175906
transform 1 0 23968 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_206
timestamp 1698175906
transform 1 0 24416 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_241
timestamp 1698175906
transform 1 0 28336 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698175906
transform 1 0 31920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_142
timestamp 1698175906
transform 1 0 17248 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_146
timestamp 1698175906
transform 1 0 17696 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_154
timestamp 1698175906
transform 1 0 18592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_156
timestamp 1698175906
transform 1 0 18816 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_173
timestamp 1698175906
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_181
timestamp 1698175906
transform 1 0 21616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_191
timestamp 1698175906
transform 1 0 22736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_223
timestamp 1698175906
transform 1 0 26320 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_229
timestamp 1698175906
transform 1 0 26992 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_88
timestamp 1698175906
transform 1 0 11200 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_96
timestamp 1698175906
transform 1 0 12096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_103
timestamp 1698175906
transform 1 0 12880 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_135
timestamp 1698175906
transform 1 0 16464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_137
timestamp 1698175906
transform 1 0 16688 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_158
timestamp 1698175906
transform 1 0 19040 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_162
timestamp 1698175906
transform 1 0 19488 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_174
timestamp 1698175906
transform 1 0 20832 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_176
timestamp 1698175906
transform 1 0 21056 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_194
timestamp 1698175906
transform 1 0 23072 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_216
timestamp 1698175906
transform 1 0 25536 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_223
timestamp 1698175906
transform 1 0 26320 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_255
timestamp 1698175906
transform 1 0 29904 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_271
timestamp 1698175906
transform 1 0 31696 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_69
timestamp 1698175906
transform 1 0 9072 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_85
timestamp 1698175906
transform 1 0 10864 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_89
timestamp 1698175906
transform 1 0 11312 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_111
timestamp 1698175906
transform 1 0 13776 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_127
timestamp 1698175906
transform 1 0 15568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_146
timestamp 1698175906
transform 1 0 17696 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_161
timestamp 1698175906
transform 1 0 19376 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_169
timestamp 1698175906
transform 1 0 20272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_173
timestamp 1698175906
transform 1 0 20720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_179
timestamp 1698175906
transform 1 0 21392 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_190
timestamp 1698175906
transform 1 0 22624 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_222
timestamp 1698175906
transform 1 0 26208 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_238
timestamp 1698175906
transform 1 0 28000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698175906
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 4480 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_76
timestamp 1698175906
transform 1 0 9856 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_107
timestamp 1698175906
transform 1 0 13328 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698175906
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_165
timestamp 1698175906
transform 1 0 19824 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_169
timestamp 1698175906
transform 1 0 20272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_171
timestamp 1698175906
transform 1 0 20496 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_174
timestamp 1698175906
transform 1 0 20832 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698175906
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_220
timestamp 1698175906
transform 1 0 25984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_222
timestamp 1698175906
transform 1 0 26208 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_228
timestamp 1698175906
transform 1 0 26880 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_260
timestamp 1698175906
transform 1 0 30464 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 36512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 37408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_69
timestamp 1698175906
transform 1 0 9072 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_85
timestamp 1698175906
transform 1 0 10864 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_93
timestamp 1698175906
transform 1 0 11760 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698175906
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_193
timestamp 1698175906
transform 1 0 22960 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_201
timestamp 1698175906
transform 1 0 23856 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_203
timestamp 1698175906
transform 1 0 24080 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698175906
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_148
timestamp 1698175906
transform 1 0 17920 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_152
timestamp 1698175906
transform 1 0 18368 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_168
timestamp 1698175906
transform 1 0 20160 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_200
timestamp 1698175906
transform 1 0 23744 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698175906
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_168
timestamp 1698175906
transform 1 0 20160 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_200
timestamp 1698175906
transform 1 0 23744 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_208
timestamp 1698175906
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita55_26 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17024 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17584 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform -1 0 4480 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 37520 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 4480 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform -1 0 20384 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 25648 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 20944 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 20272 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 23632 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 4480 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 37520 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 17360 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 18144 41200 18256 42000 0 FreeSans 448 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 16800 41200 16912 42000 0 FreeSans 448 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 41200 26208 42000 26320 0 FreeSans 448 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 41200 17472 42000 17584 0 FreeSans 448 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 22848 41200 22960 42000 0 FreeSans 448 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 17472 41200 17584 42000 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 41200 26880 42000 26992 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 41200 20160 42000 20272 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 12264 21112 12264 21112 0 _000_
rlabel metal2 15176 27384 15176 27384 0 _001_
rlabel metal3 12040 25704 12040 25704 0 _002_
rlabel metal2 26152 19544 26152 19544 0 _003_
rlabel metal2 25480 23184 25480 23184 0 _004_
rlabel metal2 14952 23576 14952 23576 0 _005_
rlabel metal2 23688 18872 23688 18872 0 _006_
rlabel metal3 23856 16184 23856 16184 0 _007_
rlabel metal2 14728 17136 14728 17136 0 _008_
rlabel metal2 26264 20160 26264 20160 0 _009_
rlabel metal2 21784 13328 21784 13328 0 _010_
rlabel metal2 21448 27440 21448 27440 0 _011_
rlabel metal3 17696 15176 17696 15176 0 _012_
rlabel metal2 18536 13328 18536 13328 0 _013_
rlabel metal2 13160 22792 13160 22792 0 _014_
rlabel metal3 22792 14616 22792 14616 0 _015_
rlabel metal2 16072 25872 16072 25872 0 _016_
rlabel metal2 14728 14560 14728 14560 0 _017_
rlabel metal2 25368 26712 25368 26712 0 _018_
rlabel metal2 24360 23520 24360 23520 0 _019_
rlabel metal3 16856 19432 16856 19432 0 _020_
rlabel metal2 13496 17920 13496 17920 0 _021_
rlabel metal2 21784 25928 21784 25928 0 _022_
rlabel metal2 18872 26684 18872 26684 0 _023_
rlabel metal2 12376 24976 12376 24976 0 _024_
rlabel metal2 21672 18032 21672 18032 0 _025_
rlabel metal3 28056 19768 28056 19768 0 _026_
rlabel metal2 25704 23968 25704 23968 0 _027_
rlabel metal3 15232 23016 15232 23016 0 _028_
rlabel metal3 21224 17528 21224 17528 0 _029_
rlabel metal2 22792 18480 22792 18480 0 _030_
rlabel metal2 23408 18200 23408 18200 0 _031_
rlabel metal3 23968 17752 23968 17752 0 _032_
rlabel metal3 21112 17752 21112 17752 0 _033_
rlabel metal2 22568 17528 22568 17528 0 _034_
rlabel metal2 18648 17696 18648 17696 0 _035_
rlabel metal3 26880 20776 26880 20776 0 _036_
rlabel metal2 21896 13160 21896 13160 0 _037_
rlabel metal2 19432 20272 19432 20272 0 _038_
rlabel metal2 19432 14000 19432 14000 0 _039_
rlabel metal2 22120 13608 22120 13608 0 _040_
rlabel metal2 22232 27272 22232 27272 0 _041_
rlabel metal2 19208 16856 19208 16856 0 _042_
rlabel metal2 19096 14616 19096 14616 0 _043_
rlabel metal2 19712 13832 19712 13832 0 _044_
rlabel metal3 16856 21784 16856 21784 0 _045_
rlabel metal2 15288 22624 15288 22624 0 _046_
rlabel metal2 22792 15456 22792 15456 0 _047_
rlabel metal2 21672 16352 21672 16352 0 _048_
rlabel metal2 16632 25536 16632 25536 0 _049_
rlabel metal2 21784 22008 21784 22008 0 _050_
rlabel metal2 18256 17528 18256 17528 0 _051_
rlabel metal2 22904 21000 22904 21000 0 _052_
rlabel metal2 20552 21672 20552 21672 0 _053_
rlabel metal2 18648 21056 18648 21056 0 _054_
rlabel metal3 19040 21000 19040 21000 0 _055_
rlabel metal2 18088 21056 18088 21056 0 _056_
rlabel metal2 18536 17248 18536 17248 0 _057_
rlabel metal2 17864 15736 17864 15736 0 _058_
rlabel metal2 16632 19992 16632 19992 0 _059_
rlabel metal3 21056 17640 21056 17640 0 _060_
rlabel metal3 18480 15512 18480 15512 0 _061_
rlabel metal2 22456 24976 22456 24976 0 _062_
rlabel metal2 22792 16856 22792 16856 0 _063_
rlabel metal2 20328 13328 20328 13328 0 _064_
rlabel metal3 17360 22344 17360 22344 0 _065_
rlabel metal3 23968 25480 23968 25480 0 _066_
rlabel metal3 22624 23688 22624 23688 0 _067_
rlabel metal3 17584 26264 17584 26264 0 _068_
rlabel metal2 20552 24192 20552 24192 0 _069_
rlabel metal3 19712 23800 19712 23800 0 _070_
rlabel metal2 16968 24584 16968 24584 0 _071_
rlabel metal2 27720 20552 27720 20552 0 _072_
rlabel metal2 26152 26264 26152 26264 0 _073_
rlabel metal2 21448 17808 21448 17808 0 _074_
rlabel metal3 26376 20664 26376 20664 0 _075_
rlabel metal2 26208 23688 26208 23688 0 _076_
rlabel metal2 17752 18872 17752 18872 0 _077_
rlabel metal2 18312 20048 18312 20048 0 _078_
rlabel metal2 13832 17976 13832 17976 0 _079_
rlabel metal2 15736 21616 15736 21616 0 _080_
rlabel metal3 13412 25368 13412 25368 0 _081_
rlabel metal2 22008 25368 22008 25368 0 _082_
rlabel metal2 18424 25984 18424 25984 0 _083_
rlabel metal2 19656 22064 19656 22064 0 _084_
rlabel metal2 12488 20944 12488 20944 0 _085_
rlabel metal2 14280 23352 14280 23352 0 _086_
rlabel metal2 12600 20888 12600 20888 0 _087_
rlabel metal3 18872 26824 18872 26824 0 _088_
rlabel metal2 19096 24080 19096 24080 0 _089_
rlabel metal2 17416 20496 17416 20496 0 _090_
rlabel metal2 17752 27048 17752 27048 0 _091_
rlabel metal3 2478 27608 2478 27608 0 clk
rlabel metal2 23128 18368 23128 18368 0 clknet_0_clk
rlabel metal2 24584 14112 24584 14112 0 clknet_1_0__leaf_clk
rlabel metal2 14392 26096 14392 26096 0 clknet_1_1__leaf_clk
rlabel metal2 15960 20720 15960 20720 0 dut55.count\[0\]
rlabel metal2 15064 18592 15064 18592 0 dut55.count\[1\]
rlabel metal2 23464 24360 23464 24360 0 dut55.count\[2\]
rlabel metal2 22568 24080 22568 24080 0 dut55.count\[3\]
rlabel metal2 17864 6748 17864 6748 0 net1
rlabel metal2 19712 3528 19712 3528 0 net10
rlabel metal2 25816 9716 25816 9716 0 net11
rlabel metal2 21112 5964 21112 5964 0 net12
rlabel metal2 20440 6356 20440 6356 0 net13
rlabel metal2 4312 23856 4312 23856 0 net14
rlabel metal2 23800 6748 23800 6748 0 net15
rlabel metal3 24080 27720 24080 27720 0 net16
rlabel metal2 26936 23016 26936 23016 0 net17
rlabel metal2 28280 19712 28280 19712 0 net18
rlabel metal2 12152 26992 12152 26992 0 net19
rlabel metal3 6356 23128 6356 23128 0 net2
rlabel metal2 17304 27272 17304 27272 0 net20
rlabel metal2 4312 21896 4312 21896 0 net21
rlabel metal2 28168 23464 28168 23464 0 net22
rlabel metal2 37912 26600 37912 26600 0 net23
rlabel metal3 28000 20552 28000 20552 0 net24
rlabel metal2 17528 6356 17528 6356 0 net25
rlabel metal2 17304 38248 17304 38248 0 net26
rlabel metal3 25368 3528 25368 3528 0 net3
rlabel metal3 16856 26152 16856 26152 0 net4
rlabel metal3 37576 21560 37576 21560 0 net5
rlabel metal2 27944 27104 27944 27104 0 net6
rlabel metal2 12152 25816 12152 25816 0 net7
rlabel metal2 26936 16912 26936 16912 0 net8
rlabel metal2 10248 25816 10248 25816 0 net9
rlabel metal2 17528 854 17528 854 0 segm[10]
rlabel metal3 1358 22904 1358 22904 0 segm[11]
rlabel metal2 22904 2198 22904 2198 0 segm[12]
rlabel metal3 17640 37464 17640 37464 0 segm[13]
rlabel metal2 39928 21168 39928 21168 0 segm[1]
rlabel metal2 40040 26712 40040 26712 0 segm[2]
rlabel metal3 1358 25592 1358 25592 0 segm[3]
rlabel metal2 40040 17640 40040 17640 0 segm[4]
rlabel metal3 1414 24920 1414 24920 0 segm[5]
rlabel metal2 18872 2198 18872 2198 0 segm[6]
rlabel metal2 25592 854 25592 854 0 segm[7]
rlabel metal2 20888 2198 20888 2198 0 segm[8]
rlabel metal2 20216 2422 20216 2422 0 segm[9]
rlabel metal3 1358 23576 1358 23576 0 sel[0]
rlabel metal2 23576 2982 23576 2982 0 sel[10]
rlabel metal3 24248 38248 24248 38248 0 sel[11]
rlabel metal3 40642 22904 40642 22904 0 sel[1]
rlabel metal2 40040 19656 40040 19656 0 sel[2]
rlabel metal3 1358 26264 1358 26264 0 sel[3]
rlabel metal3 18088 38248 18088 38248 0 sel[4]
rlabel metal3 1358 21560 1358 21560 0 sel[5]
rlabel metal2 40040 23800 40040 23800 0 sel[6]
rlabel metal2 39928 26488 39928 26488 0 sel[7]
rlabel metal2 40040 20552 40040 20552 0 sel[8]
rlabel metal2 18200 2422 18200 2422 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
