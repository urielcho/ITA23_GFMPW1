magic
tech gf180mcuD
magscale 1 10
timestamp 1699641798
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 22430 38274 22482 38286
rect 22430 38210 22482 38222
rect 26126 38274 26178 38286
rect 26126 38210 26178 38222
rect 18834 38110 18846 38162
rect 18898 38110 18910 38162
rect 17602 37998 17614 38050
rect 17666 37998 17678 38050
rect 21746 37998 21758 38050
rect 21810 37998 21822 38050
rect 25218 37998 25230 38050
rect 25282 37998 25294 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 22094 37490 22146 37502
rect 22094 37426 22146 37438
rect 40238 37378 40290 37390
rect 40238 37314 40290 37326
rect 21410 37214 21422 37266
rect 21474 37214 21486 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 19394 27806 19406 27858
rect 19458 27806 19470 27858
rect 37650 27806 37662 27858
rect 37714 27806 37726 27858
rect 22766 27746 22818 27758
rect 20066 27694 20078 27746
rect 20130 27694 20142 27746
rect 22194 27694 22206 27746
rect 22258 27694 22270 27746
rect 39890 27694 39902 27746
rect 39954 27694 39966 27746
rect 22766 27682 22818 27694
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 1934 27186 1986 27198
rect 40014 27186 40066 27198
rect 25218 27134 25230 27186
rect 25282 27134 25294 27186
rect 28466 27134 28478 27186
rect 28530 27134 28542 27186
rect 1934 27122 1986 27134
rect 40014 27122 40066 27134
rect 4274 27022 4286 27074
rect 4338 27022 4350 27074
rect 22306 27022 22318 27074
rect 22370 27022 22382 27074
rect 25554 27022 25566 27074
rect 25618 27022 25630 27074
rect 37650 27022 37662 27074
rect 37714 27022 37726 27074
rect 29262 26962 29314 26974
rect 23090 26910 23102 26962
rect 23154 26910 23166 26962
rect 26338 26910 26350 26962
rect 26402 26910 26414 26962
rect 29262 26898 29314 26910
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 23774 26514 23826 26526
rect 15362 26462 15374 26514
rect 15426 26462 15438 26514
rect 23774 26450 23826 26462
rect 27022 26514 27074 26526
rect 27022 26450 27074 26462
rect 17390 26402 17442 26414
rect 28242 26350 28254 26402
rect 28306 26350 28318 26402
rect 17390 26338 17442 26350
rect 17726 26290 17778 26302
rect 21870 26290 21922 26302
rect 4274 26238 4286 26290
rect 4338 26238 4350 26290
rect 14914 26238 14926 26290
rect 14978 26238 14990 26290
rect 15586 26238 15598 26290
rect 15650 26238 15662 26290
rect 18610 26238 18622 26290
rect 18674 26238 18686 26290
rect 17726 26226 17778 26238
rect 21870 26226 21922 26238
rect 27134 26290 27186 26302
rect 28018 26238 28030 26290
rect 28082 26238 28094 26290
rect 37874 26238 37886 26290
rect 37938 26238 37950 26290
rect 27134 26226 27186 26238
rect 23886 26178 23938 26190
rect 12114 26126 12126 26178
rect 12178 26126 12190 26178
rect 14242 26126 14254 26178
rect 14306 26126 14318 26178
rect 19282 26126 19294 26178
rect 19346 26126 19358 26178
rect 21410 26126 21422 26178
rect 21474 26126 21486 26178
rect 23886 26114 23938 26126
rect 25454 26178 25506 26190
rect 39890 26126 39902 26178
rect 39954 26126 39966 26178
rect 25454 26114 25506 26126
rect 1934 26066 1986 26078
rect 1934 26002 1986 26014
rect 27022 26066 27074 26078
rect 27022 26002 27074 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 20190 25730 20242 25742
rect 20190 25666 20242 25678
rect 20302 25730 20354 25742
rect 20302 25666 20354 25678
rect 19406 25618 19458 25630
rect 2034 25566 2046 25618
rect 2098 25566 2110 25618
rect 9986 25566 9998 25618
rect 10050 25566 10062 25618
rect 16370 25566 16382 25618
rect 16434 25566 16446 25618
rect 18498 25566 18510 25618
rect 18562 25566 18574 25618
rect 19406 25554 19458 25566
rect 21422 25618 21474 25630
rect 40014 25618 40066 25630
rect 23986 25566 23998 25618
rect 24050 25566 24062 25618
rect 28578 25566 28590 25618
rect 28642 25566 28654 25618
rect 21422 25554 21474 25566
rect 40014 25554 40066 25566
rect 19742 25506 19794 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 12786 25454 12798 25506
rect 12850 25454 12862 25506
rect 15586 25454 15598 25506
rect 15650 25454 15662 25506
rect 19742 25442 19794 25454
rect 20526 25506 20578 25518
rect 21870 25506 21922 25518
rect 20738 25454 20750 25506
rect 20802 25454 20814 25506
rect 20526 25442 20578 25454
rect 21870 25442 21922 25454
rect 24446 25506 24498 25518
rect 25666 25454 25678 25506
rect 25730 25454 25742 25506
rect 29250 25454 29262 25506
rect 29314 25454 29326 25506
rect 37650 25454 37662 25506
rect 37714 25454 37726 25506
rect 24446 25442 24498 25454
rect 14702 25394 14754 25406
rect 12114 25342 12126 25394
rect 12178 25342 12190 25394
rect 14702 25330 14754 25342
rect 14814 25394 14866 25406
rect 14814 25330 14866 25342
rect 19294 25394 19346 25406
rect 19294 25330 19346 25342
rect 19630 25394 19682 25406
rect 19630 25330 19682 25342
rect 21310 25394 21362 25406
rect 21310 25330 21362 25342
rect 21646 25394 21698 25406
rect 21646 25330 21698 25342
rect 23998 25394 24050 25406
rect 26450 25342 26462 25394
rect 26514 25342 26526 25394
rect 23998 25330 24050 25342
rect 15038 25282 15090 25294
rect 15038 25218 15090 25230
rect 24110 25282 24162 25294
rect 24110 25218 24162 25230
rect 24334 25282 24386 25294
rect 29474 25230 29486 25282
rect 29538 25230 29550 25282
rect 24334 25218 24386 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 12462 24946 12514 24958
rect 12462 24882 12514 24894
rect 20414 24946 20466 24958
rect 20414 24882 20466 24894
rect 20526 24946 20578 24958
rect 26798 24946 26850 24958
rect 23762 24894 23774 24946
rect 23826 24894 23838 24946
rect 20526 24882 20578 24894
rect 26798 24882 26850 24894
rect 27694 24946 27746 24958
rect 27694 24882 27746 24894
rect 13470 24834 13522 24846
rect 13470 24770 13522 24782
rect 15150 24834 15202 24846
rect 15150 24770 15202 24782
rect 15486 24834 15538 24846
rect 15486 24770 15538 24782
rect 26126 24834 26178 24846
rect 26126 24770 26178 24782
rect 26238 24834 26290 24846
rect 26238 24770 26290 24782
rect 27022 24834 27074 24846
rect 27022 24770 27074 24782
rect 13694 24722 13746 24734
rect 13694 24658 13746 24670
rect 13918 24722 13970 24734
rect 15374 24722 15426 24734
rect 14130 24670 14142 24722
rect 14194 24670 14206 24722
rect 13918 24658 13970 24670
rect 15374 24658 15426 24670
rect 15710 24722 15762 24734
rect 15710 24658 15762 24670
rect 20302 24722 20354 24734
rect 27134 24722 27186 24734
rect 20850 24670 20862 24722
rect 20914 24670 20926 24722
rect 23538 24670 23550 24722
rect 23602 24670 23614 24722
rect 20302 24658 20354 24670
rect 27134 24658 27186 24670
rect 27582 24722 27634 24734
rect 37650 24670 37662 24722
rect 37714 24670 37726 24722
rect 27582 24658 27634 24670
rect 12574 24610 12626 24622
rect 12574 24546 12626 24558
rect 13806 24610 13858 24622
rect 13806 24546 13858 24558
rect 28814 24610 28866 24622
rect 28814 24546 28866 24558
rect 15934 24498 15986 24510
rect 15934 24434 15986 24446
rect 26126 24498 26178 24510
rect 26126 24434 26178 24446
rect 27694 24498 27746 24510
rect 27694 24434 27746 24446
rect 40014 24498 40066 24510
rect 40014 24434 40066 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 27694 24162 27746 24174
rect 18162 24110 18174 24162
rect 18226 24110 18238 24162
rect 22082 24110 22094 24162
rect 22146 24110 22158 24162
rect 27694 24098 27746 24110
rect 40014 24050 40066 24062
rect 40014 23986 40066 23998
rect 13918 23938 13970 23950
rect 13918 23874 13970 23886
rect 15598 23938 15650 23950
rect 15598 23874 15650 23886
rect 15822 23938 15874 23950
rect 27582 23938 27634 23950
rect 18050 23886 18062 23938
rect 18114 23886 18126 23938
rect 22082 23886 22094 23938
rect 22146 23886 22158 23938
rect 22978 23886 22990 23938
rect 23042 23886 23054 23938
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 15822 23874 15874 23886
rect 27582 23874 27634 23886
rect 18734 23826 18786 23838
rect 18498 23774 18510 23826
rect 18562 23774 18574 23826
rect 18734 23762 18786 23774
rect 21534 23826 21586 23838
rect 23550 23826 23602 23838
rect 21746 23774 21758 23826
rect 21810 23774 21822 23826
rect 22754 23774 22766 23826
rect 22818 23774 22830 23826
rect 21534 23762 21586 23774
rect 23550 23762 23602 23774
rect 23662 23826 23714 23838
rect 23662 23762 23714 23774
rect 22318 23714 22370 23726
rect 13570 23662 13582 23714
rect 13634 23662 13646 23714
rect 16146 23662 16158 23714
rect 16210 23662 16222 23714
rect 18386 23662 18398 23714
rect 18450 23662 18462 23714
rect 22318 23650 22370 23662
rect 23326 23714 23378 23726
rect 23326 23650 23378 23662
rect 24894 23714 24946 23726
rect 24894 23650 24946 23662
rect 27694 23714 27746 23726
rect 27694 23650 27746 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 15934 23378 15986 23390
rect 15934 23314 15986 23326
rect 19742 23378 19794 23390
rect 19742 23314 19794 23326
rect 19966 23378 20018 23390
rect 19966 23314 20018 23326
rect 20862 23378 20914 23390
rect 20862 23314 20914 23326
rect 20974 23378 21026 23390
rect 20974 23314 21026 23326
rect 17838 23266 17890 23278
rect 25678 23266 25730 23278
rect 15362 23214 15374 23266
rect 15426 23263 15438 23266
rect 15698 23263 15710 23266
rect 15426 23217 15710 23263
rect 15426 23214 15438 23217
rect 15698 23214 15710 23217
rect 15762 23214 15774 23266
rect 16482 23214 16494 23266
rect 16546 23214 16558 23266
rect 22530 23214 22542 23266
rect 22594 23214 22606 23266
rect 17838 23202 17890 23214
rect 25678 23202 25730 23214
rect 25790 23266 25842 23278
rect 25790 23202 25842 23214
rect 27022 23266 27074 23278
rect 27022 23202 27074 23214
rect 27134 23266 27186 23278
rect 28242 23214 28254 23266
rect 28306 23214 28318 23266
rect 29362 23214 29374 23266
rect 29426 23214 29438 23266
rect 27134 23202 27186 23214
rect 17950 23154 18002 23166
rect 12338 23102 12350 23154
rect 12402 23102 12414 23154
rect 16706 23102 16718 23154
rect 16770 23102 16782 23154
rect 17950 23090 18002 23102
rect 18174 23154 18226 23166
rect 18174 23090 18226 23102
rect 18510 23154 18562 23166
rect 18510 23090 18562 23102
rect 19630 23154 19682 23166
rect 19630 23090 19682 23102
rect 21086 23154 21138 23166
rect 21086 23090 21138 23102
rect 21534 23154 21586 23166
rect 25566 23154 25618 23166
rect 21858 23102 21870 23154
rect 21922 23102 21934 23154
rect 26002 23102 26014 23154
rect 26066 23102 26078 23154
rect 28018 23102 28030 23154
rect 28082 23102 28094 23154
rect 29138 23102 29150 23154
rect 29202 23102 29214 23154
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 21534 23090 21586 23102
rect 25566 23090 25618 23102
rect 13010 22990 13022 23042
rect 13074 22990 13086 23042
rect 15138 22990 15150 23042
rect 15202 22990 15214 23042
rect 24658 22990 24670 23042
rect 24722 22990 24734 23042
rect 15822 22930 15874 22942
rect 15822 22866 15874 22878
rect 16158 22930 16210 22942
rect 16158 22866 16210 22878
rect 18398 22930 18450 22942
rect 18398 22866 18450 22878
rect 26462 22930 26514 22942
rect 26462 22866 26514 22878
rect 27022 22930 27074 22942
rect 27022 22866 27074 22878
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 16718 22594 16770 22606
rect 16718 22530 16770 22542
rect 17390 22594 17442 22606
rect 17390 22530 17442 22542
rect 17726 22594 17778 22606
rect 17726 22530 17778 22542
rect 19854 22594 19906 22606
rect 19854 22530 19906 22542
rect 21646 22594 21698 22606
rect 21646 22530 21698 22542
rect 1934 22482 1986 22494
rect 1934 22418 1986 22430
rect 16606 22482 16658 22494
rect 40014 22482 40066 22494
rect 25330 22430 25342 22482
rect 25394 22430 25406 22482
rect 16606 22418 16658 22430
rect 40014 22418 40066 22430
rect 13694 22370 13746 22382
rect 4162 22318 4174 22370
rect 4226 22318 4238 22370
rect 13694 22306 13746 22318
rect 14030 22370 14082 22382
rect 18734 22370 18786 22382
rect 17714 22318 17726 22370
rect 17778 22318 17790 22370
rect 18498 22318 18510 22370
rect 18562 22318 18574 22370
rect 19842 22318 19854 22370
rect 19906 22318 19918 22370
rect 22306 22318 22318 22370
rect 22370 22318 22382 22370
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 14030 22306 14082 22318
rect 18734 22306 18786 22318
rect 20190 22258 20242 22270
rect 20190 22194 20242 22206
rect 21758 22258 21810 22270
rect 21758 22194 21810 22206
rect 13918 22146 13970 22158
rect 16270 22146 16322 22158
rect 15922 22094 15934 22146
rect 15986 22094 15998 22146
rect 13918 22082 13970 22094
rect 16270 22082 16322 22094
rect 18286 22146 18338 22158
rect 18286 22082 18338 22094
rect 19406 22146 19458 22158
rect 19406 22082 19458 22094
rect 21310 22146 21362 22158
rect 21310 22082 21362 22094
rect 21534 22146 21586 22158
rect 21534 22082 21586 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 28926 21810 28978 21822
rect 28926 21746 28978 21758
rect 12910 21698 12962 21710
rect 17390 21698 17442 21710
rect 15810 21646 15822 21698
rect 15874 21646 15886 21698
rect 12910 21634 12962 21646
rect 17390 21634 17442 21646
rect 17502 21698 17554 21710
rect 18622 21698 18674 21710
rect 18274 21646 18286 21698
rect 18338 21646 18350 21698
rect 17502 21634 17554 21646
rect 18622 21634 18674 21646
rect 18846 21698 18898 21710
rect 22306 21646 22318 21698
rect 22370 21646 22382 21698
rect 18846 21634 18898 21646
rect 13022 21586 13074 21598
rect 11666 21534 11678 21586
rect 11730 21534 11742 21586
rect 12450 21534 12462 21586
rect 12514 21534 12526 21586
rect 13022 21522 13074 21534
rect 16158 21586 16210 21598
rect 16158 21522 16210 21534
rect 16718 21586 16770 21598
rect 16718 21522 16770 21534
rect 16830 21586 16882 21598
rect 16830 21522 16882 21534
rect 17950 21586 18002 21598
rect 17950 21522 18002 21534
rect 19182 21586 19234 21598
rect 19394 21534 19406 21586
rect 19458 21534 19470 21586
rect 25554 21534 25566 21586
rect 25618 21534 25630 21586
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 19182 21522 19234 21534
rect 18958 21474 19010 21486
rect 40014 21474 40066 21486
rect 9538 21422 9550 21474
rect 9602 21422 9614 21474
rect 26338 21422 26350 21474
rect 26402 21422 26414 21474
rect 28466 21422 28478 21474
rect 28530 21422 28542 21474
rect 18958 21410 19010 21422
rect 40014 21410 40066 21422
rect 12910 21362 12962 21374
rect 12910 21298 12962 21310
rect 17502 21362 17554 21374
rect 17502 21298 17554 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 14254 21026 14306 21038
rect 14254 20962 14306 20974
rect 26238 21026 26290 21038
rect 26238 20962 26290 20974
rect 11006 20914 11058 20926
rect 11006 20850 11058 20862
rect 22542 20914 22594 20926
rect 22542 20850 22594 20862
rect 26126 20914 26178 20926
rect 26126 20850 26178 20862
rect 11118 20802 11170 20814
rect 11118 20738 11170 20750
rect 11566 20802 11618 20814
rect 22990 20802 23042 20814
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 21298 20750 21310 20802
rect 21362 20750 21374 20802
rect 22754 20750 22766 20802
rect 22818 20750 22830 20802
rect 11566 20738 11618 20750
rect 22990 20738 23042 20750
rect 25678 20802 25730 20814
rect 25678 20738 25730 20750
rect 14142 20690 14194 20702
rect 23102 20690 23154 20702
rect 17378 20638 17390 20690
rect 17442 20638 17454 20690
rect 21410 20638 21422 20690
rect 21474 20638 21486 20690
rect 22194 20638 22206 20690
rect 22258 20638 22270 20690
rect 14142 20626 14194 20638
rect 23102 20626 23154 20638
rect 25342 20690 25394 20702
rect 25342 20626 25394 20638
rect 25454 20690 25506 20702
rect 25454 20626 25506 20638
rect 26014 20690 26066 20702
rect 26014 20626 26066 20638
rect 10894 20578 10946 20590
rect 13806 20578 13858 20590
rect 13458 20526 13470 20578
rect 13522 20526 13534 20578
rect 10894 20514 10946 20526
rect 13806 20514 13858 20526
rect 14254 20578 14306 20590
rect 23538 20526 23550 20578
rect 23602 20526 23614 20578
rect 14254 20514 14306 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 11454 20242 11506 20254
rect 20078 20242 20130 20254
rect 16594 20190 16606 20242
rect 16658 20190 16670 20242
rect 11454 20178 11506 20190
rect 20078 20178 20130 20190
rect 26238 20242 26290 20254
rect 26238 20178 26290 20190
rect 15150 20130 15202 20142
rect 17502 20130 17554 20142
rect 19406 20130 19458 20142
rect 15922 20078 15934 20130
rect 15986 20078 15998 20130
rect 18834 20078 18846 20130
rect 18898 20078 18910 20130
rect 15150 20066 15202 20078
rect 17502 20066 17554 20078
rect 19406 20066 19458 20078
rect 19630 20130 19682 20142
rect 19630 20066 19682 20078
rect 19742 20130 19794 20142
rect 20402 20078 20414 20130
rect 20466 20078 20478 20130
rect 20738 20078 20750 20130
rect 20802 20078 20814 20130
rect 21746 20078 21758 20130
rect 21810 20078 21822 20130
rect 27346 20078 27358 20130
rect 27410 20078 27422 20130
rect 19742 20066 19794 20078
rect 11230 20018 11282 20030
rect 14926 20018 14978 20030
rect 4274 19966 4286 20018
rect 4338 19966 4350 20018
rect 10882 19966 10894 20018
rect 10946 19966 10958 20018
rect 11778 19966 11790 20018
rect 11842 19966 11854 20018
rect 11230 19954 11282 19966
rect 14926 19954 14978 19966
rect 15262 20018 15314 20030
rect 17614 20018 17666 20030
rect 21086 20018 21138 20030
rect 15698 19966 15710 20018
rect 15762 19966 15774 20018
rect 16370 19966 16382 20018
rect 16434 19966 16446 20018
rect 17938 19966 17950 20018
rect 18002 19966 18014 20018
rect 19058 19966 19070 20018
rect 19122 19966 19134 20018
rect 21522 19966 21534 20018
rect 21586 19966 21598 20018
rect 26562 19966 26574 20018
rect 26626 19966 26638 20018
rect 37874 19966 37886 20018
rect 37938 19966 37950 20018
rect 15262 19954 15314 19966
rect 17614 19954 17666 19966
rect 21086 19954 21138 19966
rect 11342 19906 11394 19918
rect 12562 19854 12574 19906
rect 12626 19854 12638 19906
rect 14690 19854 14702 19906
rect 14754 19854 14766 19906
rect 29474 19854 29486 19906
rect 29538 19854 29550 19906
rect 11342 19842 11394 19854
rect 1934 19794 1986 19806
rect 1934 19730 1986 19742
rect 40014 19794 40066 19806
rect 40014 19730 40066 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 20178 19406 20190 19458
rect 20242 19406 20254 19458
rect 13582 19346 13634 19358
rect 8866 19294 8878 19346
rect 8930 19294 8942 19346
rect 10994 19294 11006 19346
rect 11058 19294 11070 19346
rect 13582 19282 13634 19294
rect 22542 19346 22594 19358
rect 40014 19346 40066 19358
rect 23762 19294 23774 19346
rect 23826 19294 23838 19346
rect 24994 19294 25006 19346
rect 25058 19294 25070 19346
rect 22542 19282 22594 19294
rect 40014 19282 40066 19294
rect 13470 19234 13522 19246
rect 11778 19182 11790 19234
rect 11842 19182 11854 19234
rect 13470 19170 13522 19182
rect 13694 19234 13746 19246
rect 14254 19234 14306 19246
rect 14018 19182 14030 19234
rect 14082 19182 14094 19234
rect 13694 19170 13746 19182
rect 14254 19170 14306 19182
rect 14590 19234 14642 19246
rect 14590 19170 14642 19182
rect 16158 19234 16210 19246
rect 16158 19170 16210 19182
rect 16494 19234 16546 19246
rect 17278 19234 17330 19246
rect 17950 19234 18002 19246
rect 16706 19182 16718 19234
rect 16770 19182 16782 19234
rect 17714 19182 17726 19234
rect 17778 19182 17790 19234
rect 16494 19170 16546 19182
rect 17278 19170 17330 19182
rect 17950 19170 18002 19182
rect 19070 19234 19122 19246
rect 20526 19234 20578 19246
rect 24894 19234 24946 19246
rect 19618 19182 19630 19234
rect 19682 19182 19694 19234
rect 20066 19182 20078 19234
rect 20130 19182 20142 19234
rect 21298 19182 21310 19234
rect 21362 19182 21374 19234
rect 23202 19182 23214 19234
rect 23266 19182 23278 19234
rect 24434 19182 24446 19234
rect 24498 19182 24510 19234
rect 19070 19170 19122 19182
rect 20526 19170 20578 19182
rect 24894 19170 24946 19182
rect 25454 19234 25506 19246
rect 25454 19170 25506 19182
rect 25790 19234 25842 19246
rect 25790 19170 25842 19182
rect 26014 19234 26066 19246
rect 27234 19182 27246 19234
rect 27298 19182 27310 19234
rect 37650 19182 37662 19234
rect 37714 19182 37726 19234
rect 26014 19170 26066 19182
rect 15598 19122 15650 19134
rect 15598 19058 15650 19070
rect 15934 19122 15986 19134
rect 23662 19122 23714 19134
rect 21410 19070 21422 19122
rect 21474 19070 21486 19122
rect 21970 19070 21982 19122
rect 22034 19070 22046 19122
rect 15934 19058 15986 19070
rect 23662 19058 23714 19070
rect 14478 19010 14530 19022
rect 14478 18946 14530 18958
rect 15710 19010 15762 19022
rect 15710 18946 15762 18958
rect 18286 19010 18338 19022
rect 23438 19010 23490 19022
rect 18722 18958 18734 19010
rect 18786 18958 18798 19010
rect 18286 18946 18338 18958
rect 23438 18946 23490 18958
rect 23774 19010 23826 19022
rect 23774 18946 23826 18958
rect 24670 19010 24722 19022
rect 24670 18946 24722 18958
rect 25006 19010 25058 19022
rect 25006 18946 25058 18958
rect 25790 19010 25842 19022
rect 27458 18958 27470 19010
rect 27522 18958 27534 19010
rect 25790 18946 25842 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 10894 18674 10946 18686
rect 10894 18610 10946 18622
rect 11118 18674 11170 18686
rect 11118 18610 11170 18622
rect 12910 18674 12962 18686
rect 12910 18610 12962 18622
rect 18958 18674 19010 18686
rect 18958 18610 19010 18622
rect 20638 18674 20690 18686
rect 21870 18674 21922 18686
rect 21410 18622 21422 18674
rect 21474 18622 21486 18674
rect 20638 18610 20690 18622
rect 21870 18610 21922 18622
rect 11230 18562 11282 18574
rect 11230 18498 11282 18510
rect 12686 18562 12738 18574
rect 12686 18498 12738 18510
rect 15822 18562 15874 18574
rect 15822 18498 15874 18510
rect 16382 18562 16434 18574
rect 16382 18498 16434 18510
rect 19182 18562 19234 18574
rect 19182 18498 19234 18510
rect 19294 18562 19346 18574
rect 19294 18498 19346 18510
rect 21086 18562 21138 18574
rect 21086 18498 21138 18510
rect 23550 18562 23602 18574
rect 23550 18498 23602 18510
rect 23774 18562 23826 18574
rect 23774 18498 23826 18510
rect 16046 18450 16098 18462
rect 12450 18398 12462 18450
rect 12514 18398 12526 18450
rect 13122 18398 13134 18450
rect 13186 18398 13198 18450
rect 16046 18386 16098 18398
rect 20302 18450 20354 18462
rect 20302 18386 20354 18398
rect 20750 18450 20802 18462
rect 20750 18386 20802 18398
rect 21758 18450 21810 18462
rect 21758 18386 21810 18398
rect 22094 18450 22146 18462
rect 23998 18450 24050 18462
rect 23314 18398 23326 18450
rect 23378 18398 23390 18450
rect 22094 18386 22146 18398
rect 23998 18386 24050 18398
rect 24334 18450 24386 18462
rect 24334 18386 24386 18398
rect 24670 18450 24722 18462
rect 28590 18450 28642 18462
rect 25330 18398 25342 18450
rect 25394 18398 25406 18450
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 24670 18386 24722 18398
rect 28590 18386 28642 18398
rect 12798 18338 12850 18350
rect 12798 18274 12850 18286
rect 15934 18338 15986 18350
rect 15934 18274 15986 18286
rect 24222 18338 24274 18350
rect 26002 18286 26014 18338
rect 26066 18286 26078 18338
rect 28130 18286 28142 18338
rect 28194 18286 28206 18338
rect 24222 18274 24274 18286
rect 23438 18226 23490 18238
rect 23438 18162 23490 18174
rect 40014 18226 40066 18238
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 15822 17890 15874 17902
rect 21646 17890 21698 17902
rect 21298 17838 21310 17890
rect 21362 17838 21374 17890
rect 15822 17826 15874 17838
rect 21646 17826 21698 17838
rect 1934 17778 1986 17790
rect 20302 17778 20354 17790
rect 9314 17726 9326 17778
rect 9378 17726 9390 17778
rect 1934 17714 1986 17726
rect 20302 17714 20354 17726
rect 21870 17778 21922 17790
rect 29262 17778 29314 17790
rect 26226 17726 26238 17778
rect 26290 17726 26302 17778
rect 28354 17726 28366 17778
rect 28418 17726 28430 17778
rect 21870 17714 21922 17726
rect 29262 17714 29314 17726
rect 40014 17778 40066 17790
rect 40014 17714 40066 17726
rect 14478 17666 14530 17678
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 12226 17614 12238 17666
rect 12290 17614 12302 17666
rect 14478 17602 14530 17614
rect 14814 17666 14866 17678
rect 14814 17602 14866 17614
rect 14926 17666 14978 17678
rect 14926 17602 14978 17614
rect 15598 17666 15650 17678
rect 15598 17602 15650 17614
rect 15934 17666 15986 17678
rect 15934 17602 15986 17614
rect 16382 17666 16434 17678
rect 16382 17602 16434 17614
rect 18622 17666 18674 17678
rect 18622 17602 18674 17614
rect 18958 17666 19010 17678
rect 22542 17666 22594 17678
rect 19842 17614 19854 17666
rect 19906 17614 19918 17666
rect 22306 17614 22318 17666
rect 22370 17614 22382 17666
rect 18958 17602 19010 17614
rect 22542 17602 22594 17614
rect 22766 17666 22818 17678
rect 22766 17602 22818 17614
rect 22878 17666 22930 17678
rect 25442 17614 25454 17666
rect 25506 17614 25518 17666
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 22878 17602 22930 17614
rect 15374 17554 15426 17566
rect 11442 17502 11454 17554
rect 11506 17502 11518 17554
rect 15374 17490 15426 17502
rect 14590 17442 14642 17454
rect 14590 17378 14642 17390
rect 14702 17442 14754 17454
rect 14702 17378 14754 17390
rect 15262 17442 15314 17454
rect 15262 17378 15314 17390
rect 18846 17442 18898 17454
rect 18846 17378 18898 17390
rect 22654 17442 22706 17454
rect 22654 17378 22706 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 11118 17106 11170 17118
rect 11118 17042 11170 17054
rect 15038 17106 15090 17118
rect 15038 17042 15090 17054
rect 25342 17106 25394 17118
rect 25342 17042 25394 17054
rect 11230 16994 11282 17006
rect 11230 16930 11282 16942
rect 14814 16994 14866 17006
rect 14814 16930 14866 16942
rect 20862 16994 20914 17006
rect 22530 16942 22542 16994
rect 22594 16942 22606 16994
rect 20862 16930 20914 16942
rect 19182 16882 19234 16894
rect 4274 16830 4286 16882
rect 4338 16830 4350 16882
rect 19182 16818 19234 16830
rect 19742 16882 19794 16894
rect 20290 16830 20302 16882
rect 20354 16830 20366 16882
rect 21858 16830 21870 16882
rect 21922 16830 21934 16882
rect 19742 16818 19794 16830
rect 1934 16770 1986 16782
rect 15026 16718 15038 16770
rect 15090 16718 15102 16770
rect 20178 16718 20190 16770
rect 20242 16718 20254 16770
rect 24658 16718 24670 16770
rect 24722 16718 24734 16770
rect 1934 16706 1986 16718
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 21422 16322 21474 16334
rect 21422 16258 21474 16270
rect 21310 16210 21362 16222
rect 14690 16158 14702 16210
rect 14754 16158 14766 16210
rect 16818 16158 16830 16210
rect 16882 16158 16894 16210
rect 21310 16146 21362 16158
rect 20302 16098 20354 16110
rect 14018 16046 14030 16098
rect 14082 16046 14094 16098
rect 19842 16046 19854 16098
rect 19906 16046 19918 16098
rect 20302 16034 20354 16046
rect 17166 15986 17218 15998
rect 17166 15922 17218 15934
rect 17278 15986 17330 15998
rect 17278 15922 17330 15934
rect 18734 15986 18786 15998
rect 18734 15922 18786 15934
rect 19070 15986 19122 15998
rect 19070 15922 19122 15934
rect 19406 15986 19458 15998
rect 19406 15922 19458 15934
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 21870 15538 21922 15550
rect 21870 15474 21922 15486
rect 15026 15374 15038 15426
rect 15090 15374 15102 15426
rect 20626 15374 20638 15426
rect 20690 15374 20702 15426
rect 15810 15262 15822 15314
rect 15874 15262 15886 15314
rect 21410 15262 21422 15314
rect 21474 15262 21486 15314
rect 12898 15150 12910 15202
rect 12962 15150 12974 15202
rect 18498 15150 18510 15202
rect 18562 15150 18574 15202
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 18274 14590 18286 14642
rect 18338 14590 18350 14642
rect 20402 14590 20414 14642
rect 20466 14590 20478 14642
rect 17490 14478 17502 14530
rect 17554 14478 17566 14530
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 17042 3502 17054 3554
rect 17106 3502 17118 3554
rect 18062 3330 18114 3342
rect 18062 3266 18114 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 22430 38222 22482 38274
rect 26126 38222 26178 38274
rect 18846 38110 18898 38162
rect 17614 37998 17666 38050
rect 21758 37998 21810 38050
rect 25230 37998 25282 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 22094 37438 22146 37490
rect 40238 37326 40290 37378
rect 21422 37214 21474 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 19406 27806 19458 27858
rect 37662 27806 37714 27858
rect 20078 27694 20130 27746
rect 22206 27694 22258 27746
rect 22766 27694 22818 27746
rect 39902 27694 39954 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 1934 27134 1986 27186
rect 25230 27134 25282 27186
rect 28478 27134 28530 27186
rect 40014 27134 40066 27186
rect 4286 27022 4338 27074
rect 22318 27022 22370 27074
rect 25566 27022 25618 27074
rect 37662 27022 37714 27074
rect 23102 26910 23154 26962
rect 26350 26910 26402 26962
rect 29262 26910 29314 26962
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 15374 26462 15426 26514
rect 23774 26462 23826 26514
rect 27022 26462 27074 26514
rect 17390 26350 17442 26402
rect 28254 26350 28306 26402
rect 4286 26238 4338 26290
rect 14926 26238 14978 26290
rect 15598 26238 15650 26290
rect 17726 26238 17778 26290
rect 18622 26238 18674 26290
rect 21870 26238 21922 26290
rect 27134 26238 27186 26290
rect 28030 26238 28082 26290
rect 37886 26238 37938 26290
rect 12126 26126 12178 26178
rect 14254 26126 14306 26178
rect 19294 26126 19346 26178
rect 21422 26126 21474 26178
rect 23886 26126 23938 26178
rect 25454 26126 25506 26178
rect 39902 26126 39954 26178
rect 1934 26014 1986 26066
rect 27022 26014 27074 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 20190 25678 20242 25730
rect 20302 25678 20354 25730
rect 2046 25566 2098 25618
rect 9998 25566 10050 25618
rect 16382 25566 16434 25618
rect 18510 25566 18562 25618
rect 19406 25566 19458 25618
rect 21422 25566 21474 25618
rect 23998 25566 24050 25618
rect 28590 25566 28642 25618
rect 40014 25566 40066 25618
rect 4286 25454 4338 25506
rect 12798 25454 12850 25506
rect 15598 25454 15650 25506
rect 19742 25454 19794 25506
rect 20526 25454 20578 25506
rect 20750 25454 20802 25506
rect 21870 25454 21922 25506
rect 24446 25454 24498 25506
rect 25678 25454 25730 25506
rect 29262 25454 29314 25506
rect 37662 25454 37714 25506
rect 12126 25342 12178 25394
rect 14702 25342 14754 25394
rect 14814 25342 14866 25394
rect 19294 25342 19346 25394
rect 19630 25342 19682 25394
rect 21310 25342 21362 25394
rect 21646 25342 21698 25394
rect 23998 25342 24050 25394
rect 26462 25342 26514 25394
rect 15038 25230 15090 25282
rect 24110 25230 24162 25282
rect 24334 25230 24386 25282
rect 29486 25230 29538 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 12462 24894 12514 24946
rect 20414 24894 20466 24946
rect 20526 24894 20578 24946
rect 23774 24894 23826 24946
rect 26798 24894 26850 24946
rect 27694 24894 27746 24946
rect 13470 24782 13522 24834
rect 15150 24782 15202 24834
rect 15486 24782 15538 24834
rect 26126 24782 26178 24834
rect 26238 24782 26290 24834
rect 27022 24782 27074 24834
rect 13694 24670 13746 24722
rect 13918 24670 13970 24722
rect 14142 24670 14194 24722
rect 15374 24670 15426 24722
rect 15710 24670 15762 24722
rect 20302 24670 20354 24722
rect 20862 24670 20914 24722
rect 23550 24670 23602 24722
rect 27134 24670 27186 24722
rect 27582 24670 27634 24722
rect 37662 24670 37714 24722
rect 12574 24558 12626 24610
rect 13806 24558 13858 24610
rect 28814 24558 28866 24610
rect 15934 24446 15986 24498
rect 26126 24446 26178 24498
rect 27694 24446 27746 24498
rect 40014 24446 40066 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 18174 24110 18226 24162
rect 22094 24110 22146 24162
rect 27694 24110 27746 24162
rect 40014 23998 40066 24050
rect 13918 23886 13970 23938
rect 15598 23886 15650 23938
rect 15822 23886 15874 23938
rect 18062 23886 18114 23938
rect 22094 23886 22146 23938
rect 22990 23886 23042 23938
rect 27582 23886 27634 23938
rect 37662 23886 37714 23938
rect 18510 23774 18562 23826
rect 18734 23774 18786 23826
rect 21534 23774 21586 23826
rect 21758 23774 21810 23826
rect 22766 23774 22818 23826
rect 23550 23774 23602 23826
rect 23662 23774 23714 23826
rect 13582 23662 13634 23714
rect 16158 23662 16210 23714
rect 18398 23662 18450 23714
rect 22318 23662 22370 23714
rect 23326 23662 23378 23714
rect 24894 23662 24946 23714
rect 27694 23662 27746 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 15934 23326 15986 23378
rect 19742 23326 19794 23378
rect 19966 23326 20018 23378
rect 20862 23326 20914 23378
rect 20974 23326 21026 23378
rect 15374 23214 15426 23266
rect 15710 23214 15762 23266
rect 16494 23214 16546 23266
rect 17838 23214 17890 23266
rect 22542 23214 22594 23266
rect 25678 23214 25730 23266
rect 25790 23214 25842 23266
rect 27022 23214 27074 23266
rect 27134 23214 27186 23266
rect 28254 23214 28306 23266
rect 29374 23214 29426 23266
rect 12350 23102 12402 23154
rect 16718 23102 16770 23154
rect 17950 23102 18002 23154
rect 18174 23102 18226 23154
rect 18510 23102 18562 23154
rect 19630 23102 19682 23154
rect 21086 23102 21138 23154
rect 21534 23102 21586 23154
rect 21870 23102 21922 23154
rect 25566 23102 25618 23154
rect 26014 23102 26066 23154
rect 28030 23102 28082 23154
rect 29150 23102 29202 23154
rect 37662 23102 37714 23154
rect 13022 22990 13074 23042
rect 15150 22990 15202 23042
rect 24670 22990 24722 23042
rect 15822 22878 15874 22930
rect 16158 22878 16210 22930
rect 18398 22878 18450 22930
rect 26462 22878 26514 22930
rect 27022 22878 27074 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 16718 22542 16770 22594
rect 17390 22542 17442 22594
rect 17726 22542 17778 22594
rect 19854 22542 19906 22594
rect 21646 22542 21698 22594
rect 1934 22430 1986 22482
rect 16606 22430 16658 22482
rect 25342 22430 25394 22482
rect 40014 22430 40066 22482
rect 4174 22318 4226 22370
rect 13694 22318 13746 22370
rect 14030 22318 14082 22370
rect 17726 22318 17778 22370
rect 18510 22318 18562 22370
rect 18734 22318 18786 22370
rect 19854 22318 19906 22370
rect 22318 22318 22370 22370
rect 37662 22318 37714 22370
rect 20190 22206 20242 22258
rect 21758 22206 21810 22258
rect 13918 22094 13970 22146
rect 15934 22094 15986 22146
rect 16270 22094 16322 22146
rect 18286 22094 18338 22146
rect 19406 22094 19458 22146
rect 21310 22094 21362 22146
rect 21534 22094 21586 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 28926 21758 28978 21810
rect 12910 21646 12962 21698
rect 15822 21646 15874 21698
rect 17390 21646 17442 21698
rect 17502 21646 17554 21698
rect 18286 21646 18338 21698
rect 18622 21646 18674 21698
rect 18846 21646 18898 21698
rect 22318 21646 22370 21698
rect 11678 21534 11730 21586
rect 12462 21534 12514 21586
rect 13022 21534 13074 21586
rect 16158 21534 16210 21586
rect 16718 21534 16770 21586
rect 16830 21534 16882 21586
rect 17950 21534 18002 21586
rect 19182 21534 19234 21586
rect 19406 21534 19458 21586
rect 25566 21534 25618 21586
rect 37662 21534 37714 21586
rect 9550 21422 9602 21474
rect 18958 21422 19010 21474
rect 26350 21422 26402 21474
rect 28478 21422 28530 21474
rect 40014 21422 40066 21474
rect 12910 21310 12962 21362
rect 17502 21310 17554 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 14254 20974 14306 21026
rect 26238 20974 26290 21026
rect 11006 20862 11058 20914
rect 22542 20862 22594 20914
rect 26126 20862 26178 20914
rect 11118 20750 11170 20802
rect 11566 20750 11618 20802
rect 20078 20750 20130 20802
rect 21310 20750 21362 20802
rect 22766 20750 22818 20802
rect 22990 20750 23042 20802
rect 25678 20750 25730 20802
rect 14142 20638 14194 20690
rect 17390 20638 17442 20690
rect 21422 20638 21474 20690
rect 22206 20638 22258 20690
rect 23102 20638 23154 20690
rect 25342 20638 25394 20690
rect 25454 20638 25506 20690
rect 26014 20638 26066 20690
rect 10894 20526 10946 20578
rect 13470 20526 13522 20578
rect 13806 20526 13858 20578
rect 14254 20526 14306 20578
rect 23550 20526 23602 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 11454 20190 11506 20242
rect 16606 20190 16658 20242
rect 20078 20190 20130 20242
rect 26238 20190 26290 20242
rect 15150 20078 15202 20130
rect 15934 20078 15986 20130
rect 17502 20078 17554 20130
rect 18846 20078 18898 20130
rect 19406 20078 19458 20130
rect 19630 20078 19682 20130
rect 19742 20078 19794 20130
rect 20414 20078 20466 20130
rect 20750 20078 20802 20130
rect 21758 20078 21810 20130
rect 27358 20078 27410 20130
rect 4286 19966 4338 20018
rect 10894 19966 10946 20018
rect 11230 19966 11282 20018
rect 11790 19966 11842 20018
rect 14926 19966 14978 20018
rect 15262 19966 15314 20018
rect 15710 19966 15762 20018
rect 16382 19966 16434 20018
rect 17614 19966 17666 20018
rect 17950 19966 18002 20018
rect 19070 19966 19122 20018
rect 21086 19966 21138 20018
rect 21534 19966 21586 20018
rect 26574 19966 26626 20018
rect 37886 19966 37938 20018
rect 11342 19854 11394 19906
rect 12574 19854 12626 19906
rect 14702 19854 14754 19906
rect 29486 19854 29538 19906
rect 1934 19742 1986 19794
rect 40014 19742 40066 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 20190 19406 20242 19458
rect 8878 19294 8930 19346
rect 11006 19294 11058 19346
rect 13582 19294 13634 19346
rect 22542 19294 22594 19346
rect 23774 19294 23826 19346
rect 25006 19294 25058 19346
rect 40014 19294 40066 19346
rect 11790 19182 11842 19234
rect 13470 19182 13522 19234
rect 13694 19182 13746 19234
rect 14030 19182 14082 19234
rect 14254 19182 14306 19234
rect 14590 19182 14642 19234
rect 16158 19182 16210 19234
rect 16494 19182 16546 19234
rect 16718 19182 16770 19234
rect 17278 19182 17330 19234
rect 17726 19182 17778 19234
rect 17950 19182 18002 19234
rect 19070 19182 19122 19234
rect 19630 19182 19682 19234
rect 20078 19182 20130 19234
rect 20526 19182 20578 19234
rect 21310 19182 21362 19234
rect 23214 19182 23266 19234
rect 24446 19182 24498 19234
rect 24894 19182 24946 19234
rect 25454 19182 25506 19234
rect 25790 19182 25842 19234
rect 26014 19182 26066 19234
rect 27246 19182 27298 19234
rect 37662 19182 37714 19234
rect 15598 19070 15650 19122
rect 15934 19070 15986 19122
rect 21422 19070 21474 19122
rect 21982 19070 22034 19122
rect 23662 19070 23714 19122
rect 14478 18958 14530 19010
rect 15710 18958 15762 19010
rect 18286 18958 18338 19010
rect 18734 18958 18786 19010
rect 23438 18958 23490 19010
rect 23774 18958 23826 19010
rect 24670 18958 24722 19010
rect 25006 18958 25058 19010
rect 25790 18958 25842 19010
rect 27470 18958 27522 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 10894 18622 10946 18674
rect 11118 18622 11170 18674
rect 12910 18622 12962 18674
rect 18958 18622 19010 18674
rect 20638 18622 20690 18674
rect 21422 18622 21474 18674
rect 21870 18622 21922 18674
rect 11230 18510 11282 18562
rect 12686 18510 12738 18562
rect 15822 18510 15874 18562
rect 16382 18510 16434 18562
rect 19182 18510 19234 18562
rect 19294 18510 19346 18562
rect 21086 18510 21138 18562
rect 23550 18510 23602 18562
rect 23774 18510 23826 18562
rect 12462 18398 12514 18450
rect 13134 18398 13186 18450
rect 16046 18398 16098 18450
rect 20302 18398 20354 18450
rect 20750 18398 20802 18450
rect 21758 18398 21810 18450
rect 22094 18398 22146 18450
rect 23326 18398 23378 18450
rect 23998 18398 24050 18450
rect 24334 18398 24386 18450
rect 24670 18398 24722 18450
rect 25342 18398 25394 18450
rect 28590 18398 28642 18450
rect 37662 18398 37714 18450
rect 12798 18286 12850 18338
rect 15934 18286 15986 18338
rect 24222 18286 24274 18338
rect 26014 18286 26066 18338
rect 28142 18286 28194 18338
rect 23438 18174 23490 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 15822 17838 15874 17890
rect 21310 17838 21362 17890
rect 21646 17838 21698 17890
rect 1934 17726 1986 17778
rect 9326 17726 9378 17778
rect 20302 17726 20354 17778
rect 21870 17726 21922 17778
rect 26238 17726 26290 17778
rect 28366 17726 28418 17778
rect 29262 17726 29314 17778
rect 40014 17726 40066 17778
rect 4286 17614 4338 17666
rect 12238 17614 12290 17666
rect 14478 17614 14530 17666
rect 14814 17614 14866 17666
rect 14926 17614 14978 17666
rect 15598 17614 15650 17666
rect 15934 17614 15986 17666
rect 16382 17614 16434 17666
rect 18622 17614 18674 17666
rect 18958 17614 19010 17666
rect 19854 17614 19906 17666
rect 22318 17614 22370 17666
rect 22542 17614 22594 17666
rect 22766 17614 22818 17666
rect 22878 17614 22930 17666
rect 25454 17614 25506 17666
rect 37662 17614 37714 17666
rect 11454 17502 11506 17554
rect 15374 17502 15426 17554
rect 14590 17390 14642 17442
rect 14702 17390 14754 17442
rect 15262 17390 15314 17442
rect 18846 17390 18898 17442
rect 22654 17390 22706 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 11118 17054 11170 17106
rect 15038 17054 15090 17106
rect 25342 17054 25394 17106
rect 11230 16942 11282 16994
rect 14814 16942 14866 16994
rect 20862 16942 20914 16994
rect 22542 16942 22594 16994
rect 4286 16830 4338 16882
rect 19182 16830 19234 16882
rect 19742 16830 19794 16882
rect 20302 16830 20354 16882
rect 21870 16830 21922 16882
rect 1934 16718 1986 16770
rect 15038 16718 15090 16770
rect 20190 16718 20242 16770
rect 24670 16718 24722 16770
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 21422 16270 21474 16322
rect 14702 16158 14754 16210
rect 16830 16158 16882 16210
rect 21310 16158 21362 16210
rect 14030 16046 14082 16098
rect 19854 16046 19906 16098
rect 20302 16046 20354 16098
rect 17166 15934 17218 15986
rect 17278 15934 17330 15986
rect 18734 15934 18786 15986
rect 19070 15934 19122 15986
rect 19406 15934 19458 15986
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 21870 15486 21922 15538
rect 15038 15374 15090 15426
rect 20638 15374 20690 15426
rect 15822 15262 15874 15314
rect 21422 15262 21474 15314
rect 12910 15150 12962 15202
rect 18510 15150 18562 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 18286 14590 18338 14642
rect 20414 14590 20466 14642
rect 17502 14478 17554 14530
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 17054 3502 17106 3554
rect 18062 3278 18114 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 18816 41200 18928 42000
rect 20832 41200 20944 42000
rect 22176 41200 22288 42000
rect 24864 41200 24976 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 18844 38162 18900 41200
rect 18844 38110 18846 38162
rect 18898 38110 18900 38162
rect 18844 38098 18900 38110
rect 17612 38050 17668 38062
rect 17612 37998 17614 38050
rect 17666 37998 17668 38050
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 1932 27186 1988 27198
rect 1932 27134 1934 27186
rect 1986 27134 1988 27186
rect 1932 26292 1988 27134
rect 4284 27076 4340 27086
rect 4284 26982 4340 27020
rect 15372 27076 15428 27086
rect 15372 26514 15428 27020
rect 15372 26462 15374 26514
rect 15426 26462 15428 26514
rect 15372 26450 15428 26462
rect 16380 26404 16436 26414
rect 1932 26226 1988 26236
rect 4284 26292 4340 26302
rect 4284 26198 4340 26236
rect 12124 26292 12180 26302
rect 12124 26178 12180 26236
rect 14812 26292 14868 26302
rect 12124 26126 12126 26178
rect 12178 26126 12180 26178
rect 12124 26114 12180 26126
rect 14252 26178 14308 26190
rect 14252 26126 14254 26178
rect 14306 26126 14308 26178
rect 1932 26066 1988 26078
rect 1932 26014 1934 26066
rect 1986 26014 1988 26066
rect 1932 25620 1988 26014
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 1932 25554 1988 25564
rect 2044 25618 2100 25630
rect 2044 25566 2046 25618
rect 2098 25566 2100 25618
rect 2044 24948 2100 25566
rect 9996 25618 10052 25630
rect 9996 25566 9998 25618
rect 10050 25566 10052 25618
rect 4284 25508 4340 25518
rect 4284 25414 4340 25452
rect 9996 25508 10052 25566
rect 9996 25442 10052 25452
rect 12796 25508 12852 25518
rect 12124 25396 12180 25406
rect 12124 25394 12516 25396
rect 12124 25342 12126 25394
rect 12178 25342 12516 25394
rect 12124 25340 12516 25342
rect 12124 25330 12180 25340
rect 2044 24882 2100 24892
rect 12460 24946 12516 25340
rect 12460 24894 12462 24946
rect 12514 24894 12516 24946
rect 12460 24882 12516 24894
rect 12572 24612 12628 24622
rect 12572 24518 12628 24556
rect 4476 24332 4740 24342
rect 4284 24276 4340 24286
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 1932 22482 1988 22494
rect 1932 22430 1934 22482
rect 1986 22430 1988 22482
rect 1932 21588 1988 22430
rect 1932 21522 1988 21532
rect 4172 22370 4228 22382
rect 4172 22318 4174 22370
rect 4226 22318 4228 22370
rect 4172 21476 4228 22318
rect 4284 22148 4340 24220
rect 12348 23156 12404 23166
rect 12796 23156 12852 25452
rect 13468 25396 13524 25406
rect 13468 24834 13524 25340
rect 13468 24782 13470 24834
rect 13522 24782 13524 24834
rect 13468 24770 13524 24782
rect 14252 24836 14308 26126
rect 14252 24770 14308 24780
rect 14700 25394 14756 25406
rect 14700 25342 14702 25394
rect 14754 25342 14756 25394
rect 13692 24724 13748 24734
rect 12348 23154 12852 23156
rect 12348 23102 12350 23154
rect 12402 23102 12852 23154
rect 12348 23100 12852 23102
rect 13580 24722 13748 24724
rect 13580 24670 13694 24722
rect 13746 24670 13748 24722
rect 13580 24668 13748 24670
rect 13580 23714 13636 24668
rect 13692 24658 13748 24668
rect 13916 24724 13972 24734
rect 13916 24630 13972 24668
rect 14140 24722 14196 24734
rect 14140 24670 14142 24722
rect 14194 24670 14196 24722
rect 13804 24612 13860 24622
rect 13804 24518 13860 24556
rect 13916 24500 13972 24510
rect 13916 23938 13972 24444
rect 14140 24388 14196 24670
rect 14700 24500 14756 25342
rect 14812 25394 14868 26236
rect 14924 26290 14980 26302
rect 14924 26238 14926 26290
rect 14978 26238 14980 26290
rect 14924 25508 14980 26238
rect 15596 26292 15652 26302
rect 15596 26198 15652 26236
rect 16380 25618 16436 26348
rect 17388 26404 17444 26414
rect 17388 26310 17444 26348
rect 17612 25732 17668 37998
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20860 37492 20916 41200
rect 22204 38276 22260 41200
rect 22428 38276 22484 38286
rect 22204 38274 22484 38276
rect 22204 38222 22430 38274
rect 22482 38222 22484 38274
rect 22204 38220 22484 38222
rect 22428 38210 22484 38220
rect 24892 38276 24948 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 24892 38210 24948 38220
rect 26124 38276 26180 38286
rect 26124 38182 26180 38220
rect 21756 38052 21812 38062
rect 21756 38050 21924 38052
rect 21756 37998 21758 38050
rect 21810 37998 21924 38050
rect 21756 37996 21924 37998
rect 21756 37986 21812 37996
rect 20860 37426 20916 37436
rect 21420 37266 21476 37278
rect 21420 37214 21422 37266
rect 21474 37214 21476 37266
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19404 27858 19460 27870
rect 19404 27806 19406 27858
rect 19458 27806 19460 27858
rect 17724 26292 17780 26302
rect 18620 26292 18676 26302
rect 17724 26290 17892 26292
rect 17724 26238 17726 26290
rect 17778 26238 17892 26290
rect 17724 26236 17892 26238
rect 17724 26226 17780 26236
rect 17612 25666 17668 25676
rect 16380 25566 16382 25618
rect 16434 25566 16436 25618
rect 16380 25554 16436 25566
rect 14924 25442 14980 25452
rect 15596 25508 15652 25518
rect 15596 25414 15652 25452
rect 14812 25342 14814 25394
rect 14866 25342 14868 25394
rect 14812 25330 14868 25342
rect 15036 25282 15092 25294
rect 15036 25230 15038 25282
rect 15090 25230 15092 25282
rect 15036 24836 15092 25230
rect 15148 24836 15204 24846
rect 15036 24834 15204 24836
rect 15036 24782 15150 24834
rect 15202 24782 15204 24834
rect 15036 24780 15204 24782
rect 15148 24770 15204 24780
rect 15484 24836 15540 24846
rect 15484 24742 15540 24780
rect 15708 24836 15764 24846
rect 14700 24434 14756 24444
rect 15372 24722 15428 24734
rect 15372 24670 15374 24722
rect 15426 24670 15428 24722
rect 14140 24322 14196 24332
rect 13916 23886 13918 23938
rect 13970 23886 13972 23938
rect 13916 23874 13972 23886
rect 14028 23940 14084 23950
rect 13580 23662 13582 23714
rect 13634 23662 13636 23714
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4284 22082 4340 22092
rect 11676 21588 11732 21598
rect 11004 21586 11732 21588
rect 11004 21534 11678 21586
rect 11730 21534 11732 21586
rect 11004 21532 11732 21534
rect 4172 21410 4228 21420
rect 9548 21476 9604 21486
rect 9548 21382 9604 21420
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 11004 20914 11060 21532
rect 11676 21522 11732 21532
rect 11788 21588 11844 21598
rect 12348 21588 12404 23100
rect 13020 23042 13076 23054
rect 13020 22990 13022 23042
rect 13074 22990 13076 23042
rect 13020 22596 13076 22990
rect 13020 22530 13076 22540
rect 13580 21924 13636 23662
rect 13692 22596 13748 22606
rect 13692 22370 13748 22540
rect 13692 22318 13694 22370
rect 13746 22318 13748 22370
rect 13692 22306 13748 22318
rect 14028 22370 14084 23884
rect 15372 23266 15428 24670
rect 15372 23214 15374 23266
rect 15426 23214 15428 23266
rect 15372 23202 15428 23214
rect 15596 24724 15652 24734
rect 15596 23938 15652 24668
rect 15708 24722 15764 24780
rect 15708 24670 15710 24722
rect 15762 24670 15764 24722
rect 15708 24658 15764 24670
rect 17724 24724 17780 24734
rect 15932 24498 15988 24510
rect 15932 24446 15934 24498
rect 15986 24446 15988 24498
rect 15596 23886 15598 23938
rect 15650 23886 15652 23938
rect 15148 23044 15204 23054
rect 15148 22950 15204 22988
rect 15596 22932 15652 23886
rect 15820 24388 15876 24398
rect 15820 23938 15876 24332
rect 15820 23886 15822 23938
rect 15874 23886 15876 23938
rect 15820 23604 15876 23886
rect 15932 23716 15988 24446
rect 16156 23716 16212 23726
rect 15932 23714 16548 23716
rect 15932 23662 16158 23714
rect 16210 23662 16548 23714
rect 15932 23660 16548 23662
rect 16156 23650 16212 23660
rect 15820 23538 15876 23548
rect 16492 23492 16548 23660
rect 16604 23492 16660 23502
rect 15932 23436 16436 23492
rect 16492 23436 16604 23492
rect 15932 23378 15988 23436
rect 15932 23326 15934 23378
rect 15986 23326 15988 23378
rect 15932 23314 15988 23326
rect 15708 23266 15764 23278
rect 15708 23214 15710 23266
rect 15762 23214 15764 23266
rect 15708 23156 15764 23214
rect 16044 23268 16100 23278
rect 15708 23100 15988 23156
rect 15820 22932 15876 22942
rect 15596 22930 15876 22932
rect 15596 22878 15822 22930
rect 15874 22878 15876 22930
rect 15596 22876 15876 22878
rect 14028 22318 14030 22370
rect 14082 22318 14084 22370
rect 14028 22306 14084 22318
rect 13916 22148 13972 22158
rect 13916 22146 14308 22148
rect 13916 22094 13918 22146
rect 13970 22094 14308 22146
rect 13916 22092 14308 22094
rect 13916 22082 13972 22092
rect 13356 21868 13636 21924
rect 12908 21700 12964 21710
rect 12796 21698 12964 21700
rect 12796 21646 12910 21698
rect 12962 21646 12964 21698
rect 12796 21644 12964 21646
rect 12460 21588 12516 21598
rect 12348 21532 12460 21588
rect 11004 20862 11006 20914
rect 11058 20862 11060 20914
rect 11004 20850 11060 20862
rect 11564 21364 11620 21374
rect 11116 20804 11172 20814
rect 11116 20710 11172 20748
rect 11564 20802 11620 21308
rect 11564 20750 11566 20802
rect 11618 20750 11620 20802
rect 11564 20738 11620 20750
rect 10892 20580 10948 20590
rect 11452 20580 11508 20590
rect 10892 20578 11452 20580
rect 10892 20526 10894 20578
rect 10946 20526 11452 20578
rect 10892 20524 11452 20526
rect 10892 20514 10948 20524
rect 11452 20242 11508 20524
rect 11452 20190 11454 20242
rect 11506 20190 11508 20242
rect 11452 20178 11508 20190
rect 4284 20020 4340 20030
rect 4284 19926 4340 19964
rect 8876 20020 8932 20030
rect 1932 19796 1988 19806
rect 1932 19702 1988 19740
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 8876 19346 8932 19964
rect 8876 19294 8878 19346
rect 8930 19294 8932 19346
rect 8876 18676 8932 19294
rect 8876 18610 8932 18620
rect 10892 20018 10948 20030
rect 10892 19966 10894 20018
rect 10946 19966 10948 20018
rect 10892 18674 10948 19966
rect 11228 20020 11284 20030
rect 11228 19926 11284 19964
rect 11788 20018 11844 21532
rect 12460 21494 12516 21532
rect 12796 21476 12852 21644
rect 12908 21634 12964 21644
rect 12796 21410 12852 21420
rect 13020 21588 13076 21598
rect 13356 21588 13412 21868
rect 13020 21586 13412 21588
rect 13020 21534 13022 21586
rect 13074 21534 13412 21586
rect 13020 21532 13412 21534
rect 12908 21364 12964 21374
rect 12908 21270 12964 21308
rect 13020 21140 13076 21532
rect 11788 19966 11790 20018
rect 11842 19966 11844 20018
rect 11340 19906 11396 19918
rect 11340 19854 11342 19906
rect 11394 19854 11396 19906
rect 11004 19348 11060 19358
rect 11340 19348 11396 19854
rect 11004 19346 11396 19348
rect 11004 19294 11006 19346
rect 11058 19294 11396 19346
rect 11004 19292 11396 19294
rect 11004 19282 11060 19292
rect 11788 19234 11844 19966
rect 12796 21084 13076 21140
rect 12572 19908 12628 19918
rect 12572 19814 12628 19852
rect 11788 19182 11790 19234
rect 11842 19182 11844 19234
rect 10892 18622 10894 18674
rect 10946 18622 10948 18674
rect 10892 18610 10948 18622
rect 11116 18676 11172 18686
rect 11116 18582 11172 18620
rect 11228 18564 11284 18574
rect 11228 18470 11284 18508
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1932 17780 1988 17790
rect 1932 17686 1988 17724
rect 9324 17778 9380 17790
rect 9324 17726 9326 17778
rect 9378 17726 9380 17778
rect 4284 17668 4340 17678
rect 4284 17574 4340 17612
rect 9324 17668 9380 17726
rect 11788 17668 11844 19182
rect 12684 18564 12740 18574
rect 12796 18564 12852 21084
rect 14252 21026 14308 22092
rect 14252 20974 14254 21026
rect 14306 20974 14308 21026
rect 14252 20962 14308 20974
rect 14140 20690 14196 20702
rect 14140 20638 14142 20690
rect 14194 20638 14196 20690
rect 13468 20580 13524 20590
rect 13468 19234 13524 20524
rect 13804 20578 13860 20590
rect 13804 20526 13806 20578
rect 13858 20526 13860 20578
rect 13692 20020 13748 20030
rect 13580 19908 13636 19918
rect 13580 19346 13636 19852
rect 13580 19294 13582 19346
rect 13634 19294 13636 19346
rect 13580 19282 13636 19294
rect 13468 19182 13470 19234
rect 13522 19182 13524 19234
rect 13468 19170 13524 19182
rect 13692 19234 13748 19964
rect 13692 19182 13694 19234
rect 13746 19182 13748 19234
rect 13692 19170 13748 19182
rect 13804 19236 13860 20526
rect 13916 20580 13972 20590
rect 14140 20580 14196 20638
rect 13972 20524 14196 20580
rect 14252 20580 14308 20590
rect 13916 20514 13972 20524
rect 14252 20486 14308 20524
rect 15708 20356 15764 22876
rect 15820 22866 15876 22876
rect 15932 22146 15988 23100
rect 16044 22932 16100 23212
rect 16156 22932 16212 22942
rect 16044 22930 16212 22932
rect 16044 22878 16158 22930
rect 16210 22878 16212 22930
rect 16044 22876 16212 22878
rect 16156 22866 16212 22876
rect 15932 22094 15934 22146
rect 15986 22094 15988 22146
rect 15036 20300 15764 20356
rect 15820 21698 15876 21710
rect 15820 21646 15822 21698
rect 15874 21646 15876 21698
rect 15820 20580 15876 21646
rect 15932 21364 15988 22094
rect 16268 22148 16324 22158
rect 16380 22148 16436 23436
rect 16604 23426 16660 23436
rect 16492 23268 16548 23278
rect 16492 23174 16548 23212
rect 16716 23154 16772 23166
rect 16716 23102 16718 23154
rect 16770 23102 16772 23154
rect 16492 23044 16548 23054
rect 16548 22988 16660 23044
rect 16492 22978 16548 22988
rect 16604 22484 16660 22988
rect 16716 22596 16772 23102
rect 16716 22502 16772 22540
rect 17388 22596 17444 22606
rect 16268 22146 16436 22148
rect 16268 22094 16270 22146
rect 16322 22094 16436 22146
rect 16268 22092 16436 22094
rect 16492 22482 16660 22484
rect 16492 22430 16606 22482
rect 16658 22430 16660 22482
rect 16492 22428 16660 22430
rect 16156 21588 16212 21598
rect 16156 21494 16212 21532
rect 15932 21308 16212 21364
rect 14924 20020 14980 20030
rect 14924 19926 14980 19964
rect 14700 19908 14756 19918
rect 14700 19814 14756 19852
rect 13804 19170 13860 19180
rect 14028 19236 14084 19246
rect 14252 19236 14308 19246
rect 14028 19234 14308 19236
rect 14028 19182 14030 19234
rect 14082 19182 14254 19234
rect 14306 19182 14308 19234
rect 14028 19180 14308 19182
rect 14028 19170 14084 19180
rect 14252 19170 14308 19180
rect 14588 19236 14644 19246
rect 14588 19142 14644 19180
rect 14476 19010 14532 19022
rect 14476 18958 14478 19010
rect 14530 18958 14532 19010
rect 12908 18788 12964 18798
rect 12908 18674 12964 18732
rect 12908 18622 12910 18674
rect 12962 18622 12964 18674
rect 12908 18610 12964 18622
rect 12740 18508 12852 18564
rect 13132 18564 13188 18574
rect 12684 18470 12740 18508
rect 12460 18450 12516 18462
rect 12460 18398 12462 18450
rect 12514 18398 12516 18450
rect 12236 17668 12292 17678
rect 11788 17666 12292 17668
rect 11788 17614 12238 17666
rect 12290 17614 12292 17666
rect 11788 17612 12292 17614
rect 9324 17602 9380 17612
rect 11452 17556 11508 17566
rect 11116 17554 11508 17556
rect 11116 17502 11454 17554
rect 11506 17502 11508 17554
rect 11116 17500 11508 17502
rect 11116 17106 11172 17500
rect 11452 17490 11508 17500
rect 11116 17054 11118 17106
rect 11170 17054 11172 17106
rect 11116 17042 11172 17054
rect 11228 16996 11284 17006
rect 11228 16902 11284 16940
rect 1932 16884 1988 16894
rect 1932 16770 1988 16828
rect 4284 16884 4340 16894
rect 4284 16790 4340 16828
rect 1932 16718 1934 16770
rect 1986 16718 1988 16770
rect 1932 16706 1988 16718
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 12236 16100 12292 17612
rect 12460 17668 12516 18398
rect 13132 18450 13188 18508
rect 13132 18398 13134 18450
rect 13186 18398 13188 18450
rect 13132 18386 13188 18398
rect 14476 18452 14532 18958
rect 15036 18900 15092 20300
rect 15148 20130 15204 20142
rect 15148 20078 15150 20130
rect 15202 20078 15204 20130
rect 15148 19796 15204 20078
rect 15708 20132 15764 20142
rect 15260 20018 15316 20030
rect 15260 19966 15262 20018
rect 15314 19966 15316 20018
rect 15260 19796 15316 19966
rect 15708 20018 15764 20076
rect 15708 19966 15710 20018
rect 15762 19966 15764 20018
rect 15708 19954 15764 19966
rect 15820 19796 15876 20524
rect 15260 19740 15876 19796
rect 15148 19730 15204 19740
rect 12460 17602 12516 17612
rect 12796 18338 12852 18350
rect 12796 18286 12798 18338
rect 12850 18286 12852 18338
rect 12796 16996 12852 18286
rect 14476 17668 14532 18396
rect 14476 17574 14532 17612
rect 14812 18844 15092 18900
rect 15596 19124 15652 19134
rect 15820 19124 15876 19740
rect 15932 20130 15988 20142
rect 15932 20078 15934 20130
rect 15986 20078 15988 20130
rect 15932 19684 15988 20078
rect 16156 19908 16212 21308
rect 16268 20692 16324 22092
rect 16268 20626 16324 20636
rect 16380 20020 16436 20030
rect 16492 20020 16548 22428
rect 16604 22418 16660 22428
rect 17388 21698 17444 22540
rect 17724 22594 17780 24668
rect 17836 23266 17892 26236
rect 18620 26198 18676 26236
rect 19404 26292 19460 27806
rect 20076 27746 20132 27758
rect 20076 27694 20078 27746
rect 20130 27694 20132 27746
rect 20076 26908 20132 27694
rect 20076 26852 20244 26908
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19404 26226 19460 26236
rect 19292 26178 19348 26190
rect 19292 26126 19294 26178
rect 19346 26126 19348 26178
rect 18172 25732 18228 25742
rect 18172 24162 18228 25676
rect 18508 25732 18564 25742
rect 18508 25618 18564 25676
rect 18508 25566 18510 25618
rect 18562 25566 18564 25618
rect 18508 25554 18564 25566
rect 19292 25620 19348 26126
rect 19740 25732 19796 25742
rect 19404 25620 19460 25630
rect 19740 25620 19796 25676
rect 20188 25730 20244 26852
rect 21420 26178 21476 37214
rect 21868 31948 21924 37996
rect 25228 38050 25284 38062
rect 25228 37998 25230 38050
rect 25282 37998 25284 38050
rect 22092 37492 22148 37502
rect 22092 37398 22148 37436
rect 21868 31892 22260 31948
rect 22204 27748 22260 31892
rect 22092 27746 22260 27748
rect 22092 27694 22206 27746
rect 22258 27694 22260 27746
rect 22092 27692 22260 27694
rect 22092 26908 22148 27692
rect 22204 27682 22260 27692
rect 22764 27746 22820 27758
rect 22764 27694 22766 27746
rect 22818 27694 22820 27746
rect 21868 26852 22148 26908
rect 22316 27076 22372 27086
rect 22764 27076 22820 27694
rect 25228 27186 25284 37998
rect 40236 37378 40292 37390
rect 40236 37326 40238 37378
rect 40290 37326 40292 37378
rect 40236 37044 40292 37326
rect 40236 36978 40292 36988
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 28476 27860 28532 27870
rect 28476 27188 28532 27804
rect 37660 27860 37716 27870
rect 37660 27766 37716 27804
rect 39900 27746 39956 27758
rect 39900 27694 39902 27746
rect 39954 27694 39956 27746
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 25228 27134 25230 27186
rect 25282 27134 25284 27186
rect 25228 27076 25284 27134
rect 28028 27186 28532 27188
rect 28028 27134 28478 27186
rect 28530 27134 28532 27186
rect 28028 27132 28532 27134
rect 25564 27076 25620 27086
rect 22316 27074 22820 27076
rect 22316 27022 22318 27074
rect 22370 27022 22820 27074
rect 22316 27020 22820 27022
rect 25116 27020 25284 27076
rect 25452 27074 25620 27076
rect 25452 27022 25566 27074
rect 25618 27022 25620 27074
rect 25452 27020 25620 27022
rect 21868 26516 21924 26852
rect 21420 26126 21422 26178
rect 21474 26126 21476 26178
rect 21420 25956 21476 26126
rect 21756 26460 21924 26516
rect 21756 26068 21812 26460
rect 21868 26292 21924 26302
rect 22316 26292 22372 27020
rect 23100 26962 23156 26974
rect 23100 26910 23102 26962
rect 23154 26910 23156 26962
rect 23100 26516 23156 26910
rect 23100 26450 23156 26460
rect 23772 26516 23828 26526
rect 23772 26422 23828 26460
rect 21924 26236 22372 26292
rect 21868 26198 21924 26236
rect 21756 26012 21924 26068
rect 20636 25900 21476 25956
rect 20188 25678 20190 25730
rect 20242 25678 20244 25730
rect 20188 25666 20244 25678
rect 20300 25732 20356 25742
rect 20300 25638 20356 25676
rect 19292 25618 19460 25620
rect 19292 25566 19406 25618
rect 19458 25566 19460 25618
rect 19292 25564 19460 25566
rect 19404 25554 19460 25564
rect 19516 25564 19796 25620
rect 18172 24110 18174 24162
rect 18226 24110 18228 24162
rect 18172 24098 18228 24110
rect 18732 25396 18788 25406
rect 18060 23938 18116 23950
rect 18060 23886 18062 23938
rect 18114 23886 18116 23938
rect 17836 23214 17838 23266
rect 17890 23214 17892 23266
rect 17836 23202 17892 23214
rect 17948 23716 18004 23726
rect 17948 23154 18004 23660
rect 17948 23102 17950 23154
rect 18002 23102 18004 23154
rect 17948 23090 18004 23102
rect 18060 23380 18116 23886
rect 18508 23828 18564 23838
rect 18508 23826 18676 23828
rect 18508 23774 18510 23826
rect 18562 23774 18676 23826
rect 18508 23772 18676 23774
rect 18508 23762 18564 23772
rect 18396 23714 18452 23726
rect 18396 23662 18398 23714
rect 18450 23662 18452 23714
rect 17724 22542 17726 22594
rect 17778 22542 17780 22594
rect 17724 22530 17780 22542
rect 17724 22370 17780 22382
rect 17724 22318 17726 22370
rect 17778 22318 17780 22370
rect 17388 21646 17390 21698
rect 17442 21646 17444 21698
rect 17388 21634 17444 21646
rect 17500 21700 17556 21710
rect 17500 21698 17668 21700
rect 17500 21646 17502 21698
rect 17554 21646 17668 21698
rect 17500 21644 17668 21646
rect 17500 21634 17556 21644
rect 16380 20018 16548 20020
rect 16380 19966 16382 20018
rect 16434 19966 16548 20018
rect 16380 19964 16548 19966
rect 16380 19954 16436 19964
rect 16156 19852 16324 19908
rect 15932 19618 15988 19628
rect 16156 19572 16212 19582
rect 16156 19234 16212 19516
rect 16156 19182 16158 19234
rect 16210 19182 16212 19234
rect 16156 19170 16212 19182
rect 15932 19124 15988 19134
rect 15820 19122 16100 19124
rect 15820 19070 15934 19122
rect 15986 19070 16100 19122
rect 15820 19068 16100 19070
rect 14812 17666 14868 18844
rect 15596 18676 15652 19068
rect 15932 19058 15988 19068
rect 15596 18610 15652 18620
rect 15708 19010 15764 19022
rect 15708 18958 15710 19010
rect 15762 18958 15764 19010
rect 14812 17614 14814 17666
rect 14866 17614 14868 17666
rect 14812 17602 14868 17614
rect 14924 18564 14980 18574
rect 14924 17666 14980 18508
rect 15708 17892 15764 18958
rect 15820 18900 15876 18910
rect 15820 18564 15876 18844
rect 15820 18470 15876 18508
rect 16044 18450 16100 19068
rect 16044 18398 16046 18450
rect 16098 18398 16100 18450
rect 16044 18386 16100 18398
rect 16156 18452 16212 18462
rect 16268 18452 16324 19852
rect 16492 19234 16548 19964
rect 16604 21588 16660 21598
rect 16604 20242 16660 21532
rect 16604 20190 16606 20242
rect 16658 20190 16660 20242
rect 16604 20020 16660 20190
rect 16604 19954 16660 19964
rect 16716 21586 16772 21598
rect 16716 21534 16718 21586
rect 16770 21534 16772 21586
rect 16716 20132 16772 21534
rect 16828 21588 16884 21598
rect 16828 21494 16884 21532
rect 17612 21476 17668 21644
rect 17724 21588 17780 22318
rect 18060 21700 18116 23324
rect 18172 23492 18228 23502
rect 18172 23154 18228 23436
rect 18172 23102 18174 23154
rect 18226 23102 18228 23154
rect 18172 23090 18228 23102
rect 18396 23156 18452 23662
rect 18620 23268 18676 23772
rect 18508 23156 18564 23166
rect 18396 23154 18564 23156
rect 18396 23102 18510 23154
rect 18562 23102 18564 23154
rect 18396 23100 18564 23102
rect 18508 23090 18564 23100
rect 18396 22930 18452 22942
rect 18396 22878 18398 22930
rect 18450 22878 18452 22930
rect 18396 22260 18452 22878
rect 18620 22820 18676 23212
rect 18620 22754 18676 22764
rect 18732 23826 18788 25340
rect 19292 25394 19348 25406
rect 19292 25342 19294 25394
rect 19346 25342 19348 25394
rect 19292 24948 19348 25342
rect 19292 24882 19348 24892
rect 19404 23828 19460 23838
rect 18732 23774 18734 23826
rect 18786 23774 18788 23826
rect 18284 22148 18340 22158
rect 18396 22148 18452 22204
rect 18284 22146 18452 22148
rect 18284 22094 18286 22146
rect 18338 22094 18452 22146
rect 18284 22092 18452 22094
rect 18508 22370 18564 22382
rect 18508 22318 18510 22370
rect 18562 22318 18564 22370
rect 18284 22082 18340 22092
rect 18284 21700 18340 21710
rect 18060 21698 18340 21700
rect 18060 21646 18286 21698
rect 18338 21646 18340 21698
rect 18060 21644 18340 21646
rect 17948 21588 18004 21598
rect 17724 21532 17948 21588
rect 17612 21420 17892 21476
rect 17500 21364 17556 21374
rect 17500 20804 17556 21308
rect 17500 20738 17556 20748
rect 16492 19182 16494 19234
rect 16546 19182 16548 19234
rect 16492 19170 16548 19182
rect 16716 19234 16772 20076
rect 17388 20690 17444 20702
rect 17388 20638 17390 20690
rect 17442 20638 17444 20690
rect 16716 19182 16718 19234
rect 16770 19182 16772 19234
rect 16716 19170 16772 19182
rect 17276 19236 17332 19246
rect 17276 19142 17332 19180
rect 16380 18564 16436 18574
rect 16380 18470 16436 18508
rect 16212 18396 16324 18452
rect 16156 18386 16212 18396
rect 15932 18338 15988 18350
rect 15932 18286 15934 18338
rect 15986 18286 15988 18338
rect 15820 17892 15876 17902
rect 14924 17614 14926 17666
rect 14978 17614 14980 17666
rect 14924 17602 14980 17614
rect 15036 17890 15876 17892
rect 15036 17838 15822 17890
rect 15874 17838 15876 17890
rect 15036 17836 15876 17838
rect 12796 16930 12852 16940
rect 14588 17442 14644 17454
rect 14588 17390 14590 17442
rect 14642 17390 14644 17442
rect 12236 16034 12292 16044
rect 12908 16884 12964 16894
rect 12908 15202 12964 16828
rect 14588 16884 14644 17390
rect 14700 17442 14756 17454
rect 14700 17390 14702 17442
rect 14754 17390 14756 17442
rect 14700 16996 14756 17390
rect 15036 17106 15092 17836
rect 15820 17826 15876 17836
rect 15596 17668 15652 17678
rect 15596 17574 15652 17612
rect 15932 17666 15988 18286
rect 15932 17614 15934 17666
rect 15986 17614 15988 17666
rect 15932 17602 15988 17614
rect 16380 17668 16436 17678
rect 16380 17574 16436 17612
rect 15372 17554 15428 17566
rect 15372 17502 15374 17554
rect 15426 17502 15428 17554
rect 15036 17054 15038 17106
rect 15090 17054 15092 17106
rect 15036 17042 15092 17054
rect 15260 17442 15316 17454
rect 15260 17390 15262 17442
rect 15314 17390 15316 17442
rect 14812 16996 14868 17006
rect 14700 16994 14868 16996
rect 14700 16942 14814 16994
rect 14866 16942 14868 16994
rect 14700 16940 14868 16942
rect 14812 16930 14868 16940
rect 14588 16818 14644 16828
rect 15036 16770 15092 16782
rect 15036 16718 15038 16770
rect 15090 16718 15092 16770
rect 14700 16212 14756 16222
rect 14700 16118 14756 16156
rect 14028 16100 14084 16110
rect 14028 15316 14084 16044
rect 15036 15426 15092 16718
rect 15260 16212 15316 17390
rect 15372 17332 15428 17502
rect 15372 17276 15876 17332
rect 15260 16146 15316 16156
rect 15820 15988 15876 17276
rect 16828 16212 16884 16222
rect 16828 16210 17332 16212
rect 16828 16158 16830 16210
rect 16882 16158 17332 16210
rect 16828 16156 17332 16158
rect 16828 16146 16884 16156
rect 15820 15922 15876 15932
rect 17164 15988 17220 15998
rect 17164 15894 17220 15932
rect 17276 15986 17332 16156
rect 17276 15934 17278 15986
rect 17330 15934 17332 15986
rect 15036 15374 15038 15426
rect 15090 15374 15092 15426
rect 15036 15362 15092 15374
rect 14028 15250 14084 15260
rect 15820 15316 15876 15326
rect 15820 15222 15876 15260
rect 12908 15150 12910 15202
rect 12962 15150 12964 15202
rect 12908 15138 12964 15150
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 17276 8428 17332 15934
rect 17388 15316 17444 20638
rect 17500 20132 17556 20142
rect 17500 19572 17556 20076
rect 17500 19506 17556 19516
rect 17612 20020 17668 20030
rect 17612 19236 17668 19964
rect 17836 20020 17892 21420
rect 17836 19684 17892 19964
rect 17948 20018 18004 21532
rect 17948 19966 17950 20018
rect 18002 19966 18004 20018
rect 17948 19954 18004 19966
rect 17836 19618 17892 19628
rect 17948 19796 18004 19806
rect 18284 19796 18340 21644
rect 18508 21588 18564 22318
rect 18732 22370 18788 23774
rect 19292 23772 19404 23828
rect 18732 22318 18734 22370
rect 18786 22318 18788 22370
rect 18396 21532 18564 21588
rect 18620 21698 18676 21710
rect 18620 21646 18622 21698
rect 18674 21646 18676 21698
rect 18620 21588 18676 21646
rect 18396 21364 18452 21532
rect 18620 21522 18676 21532
rect 18396 21298 18452 21308
rect 18004 19740 18340 19796
rect 18620 20580 18676 20590
rect 17724 19236 17780 19246
rect 17612 19234 17780 19236
rect 17612 19182 17726 19234
rect 17778 19182 17780 19234
rect 17612 19180 17780 19182
rect 17724 19170 17780 19180
rect 17948 19234 18004 19740
rect 17948 19182 17950 19234
rect 18002 19182 18004 19234
rect 17948 19170 18004 19182
rect 18060 19572 18116 19582
rect 18060 18900 18116 19516
rect 18060 18834 18116 18844
rect 18284 19010 18340 19022
rect 18284 18958 18286 19010
rect 18338 18958 18340 19010
rect 18284 18788 18340 18958
rect 18284 18722 18340 18732
rect 18620 17668 18676 20524
rect 18732 19908 18788 22318
rect 19068 23604 19124 23614
rect 18844 21700 18900 21710
rect 18844 21606 18900 21644
rect 18956 21588 19012 21598
rect 18956 21474 19012 21532
rect 18956 21422 18958 21474
rect 19010 21422 19012 21474
rect 18956 21410 19012 21422
rect 19068 21252 19124 23548
rect 18956 21196 19124 21252
rect 19180 21586 19236 21598
rect 19180 21534 19182 21586
rect 19234 21534 19236 21586
rect 18844 20692 18900 20702
rect 18844 20130 18900 20636
rect 18844 20078 18846 20130
rect 18898 20078 18900 20130
rect 18844 20066 18900 20078
rect 18844 19908 18900 19918
rect 18732 19852 18844 19908
rect 18844 19842 18900 19852
rect 18956 19460 19012 21196
rect 19180 20244 19236 21534
rect 19180 20178 19236 20188
rect 19292 20132 19348 23772
rect 19404 23762 19460 23772
rect 19516 22596 19572 25564
rect 19740 25506 19796 25564
rect 19740 25454 19742 25506
rect 19794 25454 19796 25506
rect 19740 25442 19796 25454
rect 20524 25506 20580 25518
rect 20524 25454 20526 25506
rect 20578 25454 20580 25506
rect 19628 25394 19684 25406
rect 19628 25342 19630 25394
rect 19682 25342 19684 25394
rect 19628 23940 19684 25342
rect 20524 25172 20580 25454
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20524 25106 20580 25116
rect 19836 25050 20100 25060
rect 20412 24948 20468 24958
rect 20412 24854 20468 24892
rect 20524 24948 20580 24958
rect 20636 24948 20692 25900
rect 21420 25620 21476 25630
rect 21196 25618 21476 25620
rect 21196 25566 21422 25618
rect 21474 25566 21476 25618
rect 21196 25564 21476 25566
rect 20748 25508 20804 25518
rect 21196 25508 21252 25564
rect 21420 25554 21476 25564
rect 20748 25506 21252 25508
rect 20748 25454 20750 25506
rect 20802 25454 21252 25506
rect 20748 25452 21252 25454
rect 21868 25506 21924 26012
rect 21868 25454 21870 25506
rect 21922 25454 21924 25506
rect 20748 25442 20804 25452
rect 21868 25442 21924 25454
rect 21308 25396 21364 25406
rect 21308 25302 21364 25340
rect 21644 25396 21700 25406
rect 21644 25302 21700 25340
rect 20524 24946 20692 24948
rect 20524 24894 20526 24946
rect 20578 24894 20692 24946
rect 20524 24892 20692 24894
rect 20748 25284 20804 25294
rect 20524 24882 20580 24892
rect 20300 24724 20356 24734
rect 19628 23874 19684 23884
rect 20188 24722 20356 24724
rect 20188 24670 20302 24722
rect 20354 24670 20356 24722
rect 20188 24668 20356 24670
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19740 23380 19796 23390
rect 19740 23286 19796 23324
rect 19964 23380 20020 23390
rect 19964 23286 20020 23324
rect 19628 23154 19684 23166
rect 19628 23102 19630 23154
rect 19682 23102 19684 23154
rect 19628 22820 19684 23102
rect 19628 22754 19684 22764
rect 19852 22596 19908 22606
rect 19516 22594 19908 22596
rect 19516 22542 19854 22594
rect 19906 22542 19908 22594
rect 19516 22540 19908 22542
rect 19852 22530 19908 22540
rect 19852 22372 19908 22382
rect 19516 22370 19908 22372
rect 19516 22318 19854 22370
rect 19906 22318 19908 22370
rect 19516 22316 19908 22318
rect 19404 22148 19460 22158
rect 19404 21586 19460 22092
rect 19404 21534 19406 21586
rect 19458 21534 19460 21586
rect 19404 21522 19460 21534
rect 19404 20132 19460 20142
rect 19292 20130 19460 20132
rect 19292 20078 19406 20130
rect 19458 20078 19460 20130
rect 19292 20076 19460 20078
rect 19404 20066 19460 20076
rect 19516 20132 19572 22316
rect 19852 22306 19908 22316
rect 20188 22258 20244 24668
rect 20300 24658 20356 24668
rect 20188 22206 20190 22258
rect 20242 22206 20244 22258
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20076 21700 20132 21710
rect 20076 20802 20132 21644
rect 20076 20750 20078 20802
rect 20130 20750 20132 20802
rect 20076 20738 20132 20750
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20076 20244 20132 20254
rect 20076 20150 20132 20188
rect 19516 20066 19572 20076
rect 19628 20130 19684 20142
rect 19628 20078 19630 20130
rect 19682 20078 19684 20130
rect 18956 19394 19012 19404
rect 19068 20020 19124 20030
rect 18956 19236 19012 19246
rect 18844 19180 18956 19236
rect 18732 19010 18788 19022
rect 18732 18958 18734 19010
rect 18786 18958 18788 19010
rect 18732 18564 18788 18958
rect 18732 18498 18788 18508
rect 18844 17668 18900 19180
rect 18956 19170 19012 19180
rect 19068 19236 19124 19964
rect 19628 19572 19684 20078
rect 19740 20132 19796 20142
rect 19740 20038 19796 20076
rect 19628 19506 19684 19516
rect 20188 19458 20244 22206
rect 20188 19406 20190 19458
rect 20242 19406 20244 19458
rect 20188 19394 20244 19406
rect 20300 20244 20356 20254
rect 19628 19236 19684 19246
rect 19068 19234 19684 19236
rect 19068 19182 19070 19234
rect 19122 19182 19630 19234
rect 19682 19182 19684 19234
rect 19068 19180 19684 19182
rect 19068 19170 19124 19180
rect 19628 19170 19684 19180
rect 20076 19234 20132 19246
rect 20300 19236 20356 20188
rect 20412 20130 20468 20142
rect 20412 20078 20414 20130
rect 20466 20078 20468 20130
rect 20412 20020 20468 20078
rect 20748 20132 20804 25228
rect 21644 24836 21700 24846
rect 20860 24722 20916 24734
rect 20860 24670 20862 24722
rect 20914 24670 20916 24722
rect 20860 23380 20916 24670
rect 21532 23828 21588 23838
rect 20860 23286 20916 23324
rect 20972 23826 21588 23828
rect 20972 23774 21534 23826
rect 21586 23774 21588 23826
rect 20972 23772 21588 23774
rect 20972 23378 21028 23772
rect 21532 23762 21588 23772
rect 20972 23326 20974 23378
rect 21026 23326 21028 23378
rect 20972 23314 21028 23326
rect 21084 23156 21140 23166
rect 20748 20038 20804 20076
rect 20972 23154 21140 23156
rect 20972 23102 21086 23154
rect 21138 23102 21140 23154
rect 20972 23100 21140 23102
rect 20412 19954 20468 19964
rect 20636 19460 20692 19470
rect 20076 19182 20078 19234
rect 20130 19182 20132 19234
rect 19852 19124 19908 19134
rect 19180 19012 19236 19022
rect 19852 19012 19908 19068
rect 18956 18676 19012 18686
rect 18956 18582 19012 18620
rect 19180 18562 19236 18956
rect 19180 18510 19182 18562
rect 19234 18510 19236 18562
rect 18956 17668 19012 17678
rect 18844 17666 19012 17668
rect 18844 17614 18958 17666
rect 19010 17614 19012 17666
rect 18844 17612 19012 17614
rect 18620 17574 18676 17612
rect 18956 17602 19012 17612
rect 18844 17442 18900 17454
rect 18844 17390 18846 17442
rect 18898 17390 18900 17442
rect 18732 15988 18788 15998
rect 18844 15988 18900 17390
rect 19180 16882 19236 18510
rect 19292 18956 19908 19012
rect 20076 19012 20132 19182
rect 19292 18562 19348 18956
rect 20076 18946 20132 18956
rect 20188 19180 20356 19236
rect 20524 19234 20580 19246
rect 20524 19182 20526 19234
rect 20578 19182 20580 19234
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19292 18510 19294 18562
rect 19346 18510 19348 18562
rect 19292 18498 19348 18510
rect 19852 17666 19908 17678
rect 19852 17614 19854 17666
rect 19906 17614 19908 17666
rect 19852 17444 19908 17614
rect 20188 17556 20244 19180
rect 20300 18450 20356 18462
rect 20524 18452 20580 19182
rect 20636 18900 20692 19404
rect 20636 18674 20692 18844
rect 20972 19124 21028 23100
rect 21084 23090 21140 23100
rect 21532 23156 21588 23166
rect 21532 23062 21588 23100
rect 21420 22820 21476 22830
rect 21308 22148 21364 22158
rect 21308 22054 21364 22092
rect 21308 20802 21364 20814
rect 21308 20750 21310 20802
rect 21362 20750 21364 20802
rect 21308 20244 21364 20750
rect 21420 20690 21476 22764
rect 21644 22594 21700 24780
rect 21980 24164 22036 26236
rect 23884 26178 23940 26190
rect 23884 26126 23886 26178
rect 23938 26126 23940 26178
rect 21868 24108 22036 24164
rect 22092 25732 22148 25742
rect 22092 24162 22148 25676
rect 23884 25620 23940 26126
rect 23996 25620 24052 25630
rect 23884 25618 24052 25620
rect 23884 25566 23998 25618
rect 24050 25566 24052 25618
rect 23884 25564 24052 25566
rect 23996 25554 24052 25564
rect 24444 25508 24500 25518
rect 24444 25414 24500 25452
rect 25116 25508 25172 27020
rect 25116 25442 25172 25452
rect 25452 26964 25508 27020
rect 25564 27010 25620 27020
rect 27020 27076 27076 27086
rect 25452 26178 25508 26908
rect 25452 26126 25454 26178
rect 25506 26126 25508 26178
rect 25452 25508 25508 26126
rect 26348 26962 26404 26974
rect 26348 26910 26350 26962
rect 26402 26910 26404 26962
rect 26236 26068 26292 26078
rect 25676 25508 25732 25518
rect 25452 25506 25732 25508
rect 25452 25454 25678 25506
rect 25730 25454 25732 25506
rect 25452 25452 25732 25454
rect 23996 25396 24052 25406
rect 23996 25302 24052 25340
rect 24108 25282 24164 25294
rect 24108 25230 24110 25282
rect 24162 25230 24164 25282
rect 23772 25172 23828 25182
rect 23772 24946 23828 25116
rect 23772 24894 23774 24946
rect 23826 24894 23828 24946
rect 23772 24882 23828 24894
rect 23548 24724 23604 24734
rect 23548 24630 23604 24668
rect 22092 24110 22094 24162
rect 22146 24110 22148 24162
rect 21756 23828 21812 23838
rect 21756 23734 21812 23772
rect 21868 23492 21924 24108
rect 22092 24098 22148 24110
rect 22092 23938 22148 23950
rect 22092 23886 22094 23938
rect 22146 23886 22148 23938
rect 22092 23716 22148 23886
rect 22764 23940 22820 23950
rect 22764 23826 22820 23884
rect 22764 23774 22766 23826
rect 22818 23774 22820 23826
rect 22764 23762 22820 23774
rect 22988 23940 23044 23950
rect 22988 23938 23604 23940
rect 22988 23886 22990 23938
rect 23042 23886 23604 23938
rect 22988 23884 23604 23886
rect 22092 23650 22148 23660
rect 22316 23716 22372 23726
rect 22316 23714 22596 23716
rect 22316 23662 22318 23714
rect 22370 23662 22596 23714
rect 22316 23660 22596 23662
rect 22316 23650 22372 23660
rect 21868 23154 21924 23436
rect 22540 23266 22596 23660
rect 22540 23214 22542 23266
rect 22594 23214 22596 23266
rect 22540 23202 22596 23214
rect 21868 23102 21870 23154
rect 21922 23102 21924 23154
rect 21868 23090 21924 23102
rect 21644 22542 21646 22594
rect 21698 22542 21700 22594
rect 21644 22530 21700 22542
rect 22316 22370 22372 22382
rect 22316 22318 22318 22370
rect 22370 22318 22372 22370
rect 21756 22258 21812 22270
rect 21756 22206 21758 22258
rect 21810 22206 21812 22258
rect 21420 20638 21422 20690
rect 21474 20638 21476 20690
rect 21420 20626 21476 20638
rect 21532 22146 21588 22158
rect 21532 22094 21534 22146
rect 21586 22094 21588 22146
rect 21532 21588 21588 22094
rect 21308 20178 21364 20188
rect 21084 20018 21140 20030
rect 21084 19966 21086 20018
rect 21138 19966 21140 20018
rect 21084 19236 21140 19966
rect 21532 20018 21588 21532
rect 21756 21028 21812 22206
rect 22316 21700 22372 22318
rect 22764 22148 22820 22158
rect 22988 22148 23044 23884
rect 23548 23826 23604 23884
rect 23548 23774 23550 23826
rect 23602 23774 23604 23826
rect 23548 23762 23604 23774
rect 23660 23828 23716 23838
rect 23660 23734 23716 23772
rect 23324 23716 23380 23726
rect 23324 23622 23380 23660
rect 22820 22092 23044 22148
rect 24108 22148 24164 25230
rect 24332 25282 24388 25294
rect 24332 25230 24334 25282
rect 24386 25230 24388 25282
rect 24332 25172 24388 25230
rect 24332 25106 24388 25116
rect 24892 23714 24948 23726
rect 24892 23662 24894 23714
rect 24946 23662 24948 23714
rect 24892 23492 24948 23662
rect 25452 23492 25508 25452
rect 25676 25442 25732 25452
rect 25676 24836 25732 24846
rect 26124 24836 26180 24846
rect 24892 23426 24948 23436
rect 25340 23436 25452 23492
rect 24668 23156 24724 23166
rect 24668 23042 24724 23100
rect 24668 22990 24670 23042
rect 24722 22990 24724 23042
rect 24668 22978 24724 22990
rect 25340 22484 25396 23436
rect 25452 23426 25508 23436
rect 25564 23940 25620 23950
rect 25564 23154 25620 23884
rect 25564 23102 25566 23154
rect 25618 23102 25620 23154
rect 25564 23090 25620 23102
rect 25676 23828 25732 24780
rect 26012 24834 26180 24836
rect 26012 24782 26126 24834
rect 26178 24782 26180 24834
rect 26012 24780 26180 24782
rect 26012 23940 26068 24780
rect 26124 24770 26180 24780
rect 26236 24834 26292 26012
rect 26236 24782 26238 24834
rect 26290 24782 26292 24834
rect 26236 24770 26292 24782
rect 26124 24500 26180 24510
rect 26348 24500 26404 26910
rect 27020 26514 27076 27020
rect 27020 26462 27022 26514
rect 27074 26462 27076 26514
rect 27020 26450 27076 26462
rect 28028 27076 28084 27132
rect 28476 27122 28532 27132
rect 27132 26292 27188 26302
rect 27132 26290 27300 26292
rect 27132 26238 27134 26290
rect 27186 26238 27300 26290
rect 27132 26236 27300 26238
rect 27132 26226 27188 26236
rect 27020 26068 27076 26078
rect 27020 25974 27076 26012
rect 26460 25396 26516 25406
rect 26460 25394 26852 25396
rect 26460 25342 26462 25394
rect 26514 25342 26852 25394
rect 26460 25340 26852 25342
rect 26460 25330 26516 25340
rect 26796 24946 26852 25340
rect 26796 24894 26798 24946
rect 26850 24894 26852 24946
rect 26796 24882 26852 24894
rect 27244 25172 27300 26236
rect 28028 26290 28084 27020
rect 37660 27074 37716 27086
rect 37660 27022 37662 27074
rect 37714 27022 37716 27074
rect 29260 26964 29316 26974
rect 29260 26870 29316 26908
rect 37660 26516 37716 27022
rect 39900 26964 39956 27694
rect 39900 26898 39956 26908
rect 40012 27186 40068 27198
rect 40012 27134 40014 27186
rect 40066 27134 40068 27186
rect 37660 26450 37716 26460
rect 28252 26404 28308 26414
rect 28252 26310 28308 26348
rect 28028 26238 28030 26290
rect 28082 26238 28084 26290
rect 28028 26226 28084 26238
rect 37884 26290 37940 26302
rect 37884 26238 37886 26290
rect 37938 26238 37940 26290
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 27020 24836 27076 24846
rect 27020 24742 27076 24780
rect 26124 24498 26404 24500
rect 26124 24446 26126 24498
rect 26178 24446 26404 24498
rect 26124 24444 26404 24446
rect 27132 24722 27188 24734
rect 27132 24670 27134 24722
rect 27186 24670 27188 24722
rect 27132 24500 27188 24670
rect 27244 24724 27300 25116
rect 27692 25620 27748 25630
rect 27692 24946 27748 25564
rect 28588 25620 28644 25630
rect 28588 25526 28644 25564
rect 29260 25620 29316 25630
rect 29260 25506 29316 25564
rect 29260 25454 29262 25506
rect 29314 25454 29316 25506
rect 29260 25442 29316 25454
rect 37660 25508 37716 25518
rect 37660 25414 37716 25452
rect 29484 25284 29540 25294
rect 29484 25190 29540 25228
rect 37884 25284 37940 26238
rect 40012 26292 40068 27134
rect 40012 26226 40068 26236
rect 39900 26178 39956 26190
rect 39900 26126 39902 26178
rect 39954 26126 39956 26178
rect 39900 25620 39956 26126
rect 39900 25554 39956 25564
rect 40012 25618 40068 25630
rect 40012 25566 40014 25618
rect 40066 25566 40068 25618
rect 37884 25218 37940 25228
rect 27692 24894 27694 24946
rect 27746 24894 27748 24946
rect 27692 24882 27748 24894
rect 40012 24948 40068 25566
rect 40012 24882 40068 24892
rect 27580 24724 27636 24734
rect 29148 24724 29204 24734
rect 27244 24722 27860 24724
rect 27244 24670 27582 24722
rect 27634 24670 27860 24722
rect 27244 24668 27860 24670
rect 27580 24658 27636 24668
rect 27692 24500 27748 24510
rect 27132 24498 27748 24500
rect 27132 24446 27694 24498
rect 27746 24446 27748 24498
rect 27132 24444 27748 24446
rect 26124 24434 26180 24444
rect 27692 24434 27748 24444
rect 27692 24164 27748 24174
rect 26012 23874 26068 23884
rect 27132 24162 27748 24164
rect 27132 24110 27694 24162
rect 27746 24110 27748 24162
rect 27132 24108 27748 24110
rect 25676 23266 25732 23772
rect 25676 23214 25678 23266
rect 25730 23214 25732 23266
rect 25340 22482 25620 22484
rect 25340 22430 25342 22482
rect 25394 22430 25620 22482
rect 25340 22428 25620 22430
rect 25340 22418 25396 22428
rect 24108 22092 24612 22148
rect 22316 21606 22372 21644
rect 22540 21924 22596 21934
rect 21756 20972 21924 21028
rect 21756 20804 21812 20814
rect 21756 20130 21812 20748
rect 21868 20580 21924 20972
rect 22540 20914 22596 21868
rect 22540 20862 22542 20914
rect 22594 20862 22596 20914
rect 22540 20850 22596 20862
rect 22764 20802 22820 22092
rect 23324 21924 23380 21934
rect 22764 20750 22766 20802
rect 22818 20750 22820 20802
rect 22204 20692 22260 20702
rect 22204 20598 22260 20636
rect 21868 20514 21924 20524
rect 21756 20078 21758 20130
rect 21810 20078 21812 20130
rect 21756 20066 21812 20078
rect 21532 19966 21534 20018
rect 21586 19966 21588 20018
rect 21532 19954 21588 19966
rect 22540 19348 22596 19358
rect 22764 19348 22820 20750
rect 22988 21812 23044 21822
rect 22988 20804 23044 21756
rect 22988 20710 23044 20748
rect 23100 20690 23156 20702
rect 23100 20638 23102 20690
rect 23154 20638 23156 20690
rect 23100 20580 23156 20638
rect 23100 20514 23156 20524
rect 22540 19346 22820 19348
rect 22540 19294 22542 19346
rect 22594 19294 22820 19346
rect 22540 19292 22820 19294
rect 23212 20020 23268 20030
rect 22540 19282 22596 19292
rect 21308 19236 21364 19246
rect 21140 19234 21364 19236
rect 21140 19182 21310 19234
rect 21362 19182 21364 19234
rect 21140 19180 21364 19182
rect 21084 19142 21140 19180
rect 21308 19170 21364 19180
rect 23212 19234 23268 19964
rect 23212 19182 23214 19234
rect 23266 19182 23268 19234
rect 23212 19170 23268 19182
rect 20972 18788 21028 19068
rect 21420 19122 21476 19134
rect 21420 19070 21422 19122
rect 21474 19070 21476 19122
rect 21420 19012 21476 19070
rect 21980 19122 22036 19134
rect 21980 19070 21982 19122
rect 22034 19070 22036 19122
rect 20972 18722 21028 18732
rect 21084 18956 21476 19012
rect 21644 19012 21700 19022
rect 21700 18956 21812 19012
rect 20636 18622 20638 18674
rect 20690 18622 20692 18674
rect 20636 18610 20692 18622
rect 21084 18564 21140 18956
rect 21644 18946 21700 18956
rect 21420 18788 21476 18798
rect 21420 18676 21476 18732
rect 21644 18676 21700 18686
rect 21420 18674 21588 18676
rect 21420 18622 21422 18674
rect 21474 18622 21588 18674
rect 21420 18620 21588 18622
rect 21420 18610 21476 18620
rect 20748 18562 21140 18564
rect 20748 18510 21086 18562
rect 21138 18510 21140 18562
rect 20748 18508 21140 18510
rect 20748 18452 20804 18508
rect 21084 18498 21140 18508
rect 20300 18398 20302 18450
rect 20354 18398 20356 18450
rect 20300 18004 20356 18398
rect 20300 17938 20356 17948
rect 20412 18450 20804 18452
rect 20412 18398 20750 18450
rect 20802 18398 20804 18450
rect 20412 18396 20804 18398
rect 20300 17780 20356 17790
rect 20412 17780 20468 18396
rect 20748 18386 20804 18396
rect 21420 18004 21476 18014
rect 21308 17892 21364 17902
rect 21308 17798 21364 17836
rect 20300 17778 20468 17780
rect 20300 17726 20302 17778
rect 20354 17726 20468 17778
rect 20300 17724 20468 17726
rect 20300 17714 20356 17724
rect 20188 17500 20468 17556
rect 19852 17388 20244 17444
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19180 16830 19182 16882
rect 19234 16830 19236 16882
rect 19180 16818 19236 16830
rect 19740 16884 19796 16894
rect 17388 15148 17444 15260
rect 18284 15986 18900 15988
rect 18284 15934 18734 15986
rect 18786 15934 18900 15986
rect 18284 15932 18900 15934
rect 19068 15988 19124 15998
rect 19404 15988 19460 15998
rect 19740 15988 19796 16828
rect 20188 16770 20244 17388
rect 20412 16996 20468 17500
rect 20860 16996 20916 17006
rect 20412 16994 20916 16996
rect 20412 16942 20862 16994
rect 20914 16942 20916 16994
rect 20412 16940 20916 16942
rect 20860 16930 20916 16940
rect 20300 16884 20356 16894
rect 20300 16790 20356 16828
rect 21308 16884 21364 16894
rect 20188 16718 20190 16770
rect 20242 16718 20244 16770
rect 19852 16098 19908 16110
rect 19852 16046 19854 16098
rect 19906 16046 19908 16098
rect 19852 15988 19908 16046
rect 20188 16100 20244 16718
rect 21308 16210 21364 16828
rect 21308 16158 21310 16210
rect 21362 16158 21364 16210
rect 21308 16146 21364 16158
rect 21420 16322 21476 17948
rect 21532 17892 21588 18620
rect 21756 18676 21812 18956
rect 21868 18676 21924 18686
rect 21980 18676 22036 19070
rect 21756 18674 22036 18676
rect 21756 18622 21870 18674
rect 21922 18622 22036 18674
rect 21756 18620 22036 18622
rect 22876 18676 22932 18686
rect 21644 18564 21700 18620
rect 21868 18610 21924 18620
rect 21644 18508 21812 18564
rect 21756 18450 21812 18508
rect 21756 18398 21758 18450
rect 21810 18398 21812 18450
rect 21756 18386 21812 18398
rect 22092 18452 22148 18462
rect 22092 18450 22372 18452
rect 22092 18398 22094 18450
rect 22146 18398 22372 18450
rect 22092 18396 22372 18398
rect 22092 18386 22148 18396
rect 21868 18004 21924 18014
rect 21644 17892 21700 17902
rect 21532 17836 21644 17892
rect 21644 17798 21700 17836
rect 21868 17778 21924 17948
rect 21868 17726 21870 17778
rect 21922 17726 21924 17778
rect 21868 17714 21924 17726
rect 22316 17666 22372 18396
rect 22316 17614 22318 17666
rect 22370 17614 22372 17666
rect 22316 17602 22372 17614
rect 22540 18228 22596 18238
rect 22540 17666 22596 18172
rect 22540 17614 22542 17666
rect 22594 17614 22596 17666
rect 22540 17602 22596 17614
rect 22764 17892 22820 17902
rect 22764 17666 22820 17836
rect 22764 17614 22766 17666
rect 22818 17614 22820 17666
rect 22764 17602 22820 17614
rect 22876 17666 22932 18620
rect 23324 18450 23380 21868
rect 23548 20580 23604 20590
rect 23548 20578 24388 20580
rect 23548 20526 23550 20578
rect 23602 20526 24388 20578
rect 23548 20524 24388 20526
rect 23548 20514 23604 20524
rect 23772 19348 23828 19358
rect 23772 19346 24052 19348
rect 23772 19294 23774 19346
rect 23826 19294 24052 19346
rect 23772 19292 24052 19294
rect 23772 19282 23828 19292
rect 23660 19124 23716 19134
rect 23660 19030 23716 19068
rect 23436 19010 23492 19022
rect 23436 18958 23438 19010
rect 23490 18958 23492 19010
rect 23436 18676 23492 18958
rect 23772 19012 23828 19022
rect 23772 18900 23828 18956
rect 23436 18610 23492 18620
rect 23548 18844 23828 18900
rect 23548 18564 23604 18844
rect 23548 18470 23604 18508
rect 23772 18562 23828 18574
rect 23772 18510 23774 18562
rect 23826 18510 23828 18562
rect 23324 18398 23326 18450
rect 23378 18398 23380 18450
rect 23324 18386 23380 18398
rect 23436 18228 23492 18238
rect 23436 18134 23492 18172
rect 22876 17614 22878 17666
rect 22930 17614 22932 17666
rect 22876 17602 22932 17614
rect 23772 17668 23828 18510
rect 23996 18450 24052 19292
rect 23996 18398 23998 18450
rect 24050 18398 24052 18450
rect 23996 18386 24052 18398
rect 24332 18450 24388 20524
rect 24444 20132 24500 20142
rect 24444 19234 24500 20076
rect 24444 19182 24446 19234
rect 24498 19182 24500 19234
rect 24444 19170 24500 19182
rect 24556 19012 24612 22092
rect 25564 21586 25620 22428
rect 25676 21812 25732 23214
rect 25676 21746 25732 21756
rect 25788 23268 25844 23278
rect 25788 21924 25844 23212
rect 27020 23268 27076 23278
rect 27020 23174 27076 23212
rect 27132 23266 27188 24108
rect 27692 24098 27748 24108
rect 27580 23940 27636 23950
rect 27804 23940 27860 24668
rect 27580 23938 27860 23940
rect 27580 23886 27582 23938
rect 27634 23886 27860 23938
rect 27580 23884 27860 23886
rect 28812 24610 28868 24622
rect 28812 24558 28814 24610
rect 28866 24558 28868 24610
rect 27580 23874 27636 23884
rect 27692 23716 27748 23726
rect 27692 23622 27748 23660
rect 27132 23214 27134 23266
rect 27186 23214 27188 23266
rect 27132 23202 27188 23214
rect 28252 23268 28308 23278
rect 28252 23174 28308 23212
rect 26012 23156 26068 23166
rect 25564 21534 25566 21586
rect 25618 21534 25620 21586
rect 25452 21364 25508 21374
rect 25340 20692 25396 20702
rect 25340 20598 25396 20636
rect 25452 20690 25508 21308
rect 25452 20638 25454 20690
rect 25506 20638 25508 20690
rect 25452 20626 25508 20638
rect 25564 20244 25620 21534
rect 25788 21140 25844 21868
rect 25788 21074 25844 21084
rect 25900 23154 26068 23156
rect 25900 23102 26014 23154
rect 26066 23102 26068 23154
rect 25900 23100 26068 23102
rect 25676 20804 25732 20814
rect 25900 20804 25956 23100
rect 26012 23090 26068 23100
rect 28028 23154 28084 23166
rect 28028 23102 28030 23154
rect 28082 23102 28084 23154
rect 26460 22930 26516 22942
rect 26460 22878 26462 22930
rect 26514 22878 26516 22930
rect 25676 20802 25956 20804
rect 25676 20750 25678 20802
rect 25730 20750 25956 20802
rect 25676 20748 25956 20750
rect 26012 22260 26068 22270
rect 25676 20738 25732 20748
rect 26012 20690 26068 22204
rect 26348 21476 26404 21486
rect 26124 21474 26404 21476
rect 26124 21422 26350 21474
rect 26402 21422 26404 21474
rect 26124 21420 26404 21422
rect 26124 20914 26180 21420
rect 26348 21410 26404 21420
rect 26236 21028 26292 21038
rect 26460 21028 26516 22878
rect 26236 21026 26516 21028
rect 26236 20974 26238 21026
rect 26290 20974 26516 21026
rect 26236 20972 26516 20974
rect 27020 22930 27076 22942
rect 27020 22878 27022 22930
rect 27074 22878 27076 22930
rect 26236 20962 26292 20972
rect 26124 20862 26126 20914
rect 26178 20862 26180 20914
rect 26124 20850 26180 20862
rect 26012 20638 26014 20690
rect 26066 20638 26068 20690
rect 25340 20188 25564 20244
rect 25004 19348 25060 19358
rect 25004 19254 25060 19292
rect 24892 19236 24948 19246
rect 24892 19142 24948 19180
rect 24668 19012 24724 19022
rect 24556 19010 24724 19012
rect 24556 18958 24670 19010
rect 24722 18958 24724 19010
rect 24556 18956 24724 18958
rect 24556 18900 24612 18956
rect 24668 18946 24724 18956
rect 25004 19012 25060 19022
rect 25004 18918 25060 18956
rect 24556 18834 24612 18844
rect 24332 18398 24334 18450
rect 24386 18398 24388 18450
rect 24332 18386 24388 18398
rect 24668 18788 24724 18798
rect 24668 18450 24724 18732
rect 24668 18398 24670 18450
rect 24722 18398 24724 18450
rect 24668 18386 24724 18398
rect 25340 18450 25396 20188
rect 25564 20178 25620 20188
rect 25788 20580 25844 20590
rect 25452 19348 25508 19358
rect 25452 19234 25508 19292
rect 25452 19182 25454 19234
rect 25506 19182 25508 19234
rect 25452 19170 25508 19182
rect 25788 19234 25844 20524
rect 25788 19182 25790 19234
rect 25842 19182 25844 19234
rect 25788 19170 25844 19182
rect 26012 19234 26068 20638
rect 26236 20244 26292 20254
rect 26236 20150 26292 20188
rect 26572 20244 26628 20254
rect 26572 20018 26628 20188
rect 27020 20188 27076 22878
rect 28028 21364 28084 23102
rect 28812 21812 28868 24558
rect 29148 23716 29204 24668
rect 37660 24724 37716 24734
rect 37660 24630 37716 24668
rect 40012 24498 40068 24510
rect 40012 24446 40014 24498
rect 40066 24446 40068 24498
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 40012 24276 40068 24446
rect 40012 24210 40068 24220
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 37660 23940 37716 23950
rect 29148 23154 29204 23660
rect 37436 23938 37716 23940
rect 37436 23886 37662 23938
rect 37714 23886 37716 23938
rect 37436 23884 37716 23886
rect 29372 23268 29428 23278
rect 29372 23174 29428 23212
rect 29148 23102 29150 23154
rect 29202 23102 29204 23154
rect 28924 21812 28980 21822
rect 28812 21810 28980 21812
rect 28812 21758 28926 21810
rect 28978 21758 28980 21810
rect 28812 21756 28980 21758
rect 28028 21298 28084 21308
rect 28476 21474 28532 21486
rect 28476 21422 28478 21474
rect 28530 21422 28532 21474
rect 28476 21364 28532 21422
rect 28476 21298 28532 21308
rect 28588 20244 28644 20254
rect 28812 20244 28868 21756
rect 28924 21746 28980 21756
rect 28644 20188 28868 20244
rect 29148 20188 29204 23102
rect 37436 22932 37492 23884
rect 37660 23874 37716 23884
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 37660 23156 37716 23166
rect 37660 23062 37716 23100
rect 37436 22866 37492 22876
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 37660 22820 37716 22830
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 37660 22370 37716 22764
rect 37660 22318 37662 22370
rect 37714 22318 37716 22370
rect 37660 22306 37716 22318
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 37660 21588 37716 21598
rect 37660 21494 37716 21532
rect 40012 21588 40068 21598
rect 40012 21474 40068 21532
rect 40012 21422 40014 21474
rect 40066 21422 40068 21474
rect 40012 21410 40068 21422
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 27020 20132 27412 20188
rect 27356 20130 27412 20132
rect 27356 20078 27358 20130
rect 27410 20078 27412 20130
rect 27356 20066 27412 20078
rect 26572 19966 26574 20018
rect 26626 19966 26628 20018
rect 26572 19954 26628 19966
rect 26012 19182 26014 19234
rect 26066 19182 26068 19234
rect 25788 19010 25844 19022
rect 25788 18958 25790 19010
rect 25842 18958 25844 19010
rect 25788 18564 25844 18958
rect 26012 18788 26068 19182
rect 27244 19234 27300 19246
rect 27244 19182 27246 19234
rect 27298 19182 27300 19234
rect 27244 19124 27300 19182
rect 28364 19236 28420 19246
rect 27244 19058 27300 19068
rect 28140 19124 28196 19134
rect 27468 19012 27524 19022
rect 27468 18918 27524 18956
rect 26012 18722 26068 18732
rect 25788 18508 26292 18564
rect 25340 18398 25342 18450
rect 25394 18398 25396 18450
rect 24220 18340 24276 18350
rect 24220 18246 24276 18284
rect 23772 17602 23828 17612
rect 24668 17668 24724 17678
rect 22652 17442 22708 17454
rect 22652 17390 22654 17442
rect 22706 17390 22708 17442
rect 21420 16270 21422 16322
rect 21474 16270 21476 16322
rect 20300 16100 20356 16110
rect 20188 16098 20356 16100
rect 20188 16046 20302 16098
rect 20354 16046 20356 16098
rect 20188 16044 20356 16046
rect 19068 15986 19460 15988
rect 19068 15934 19070 15986
rect 19122 15934 19406 15986
rect 19458 15934 19460 15986
rect 19068 15932 19460 15934
rect 17388 15092 17556 15148
rect 17500 14530 17556 15092
rect 18284 14642 18340 15932
rect 18732 15922 18788 15932
rect 19068 15922 19124 15932
rect 19404 15922 19460 15932
rect 19628 15932 19908 15988
rect 18508 15204 18564 15242
rect 18508 15138 18564 15148
rect 19628 15204 19684 15932
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19628 15138 19684 15148
rect 18284 14590 18286 14642
rect 18338 14590 18340 14642
rect 18284 14578 18340 14590
rect 20300 14644 20356 16044
rect 21420 15988 21476 16270
rect 20636 15932 21476 15988
rect 21868 17108 21924 17118
rect 21868 16882 21924 17052
rect 22540 16996 22596 17006
rect 22652 16996 22708 17390
rect 22540 16994 22708 16996
rect 22540 16942 22542 16994
rect 22594 16942 22708 16994
rect 22540 16940 22708 16942
rect 22540 16930 22596 16940
rect 21868 16830 21870 16882
rect 21922 16830 21924 16882
rect 20636 15426 20692 15932
rect 21868 15540 21924 16830
rect 24668 16770 24724 17612
rect 25340 17668 25396 18398
rect 26012 18340 26068 18350
rect 26012 18246 26068 18284
rect 26236 17778 26292 18508
rect 28140 18338 28196 19068
rect 28140 18286 28142 18338
rect 28194 18286 28196 18338
rect 28140 18274 28196 18286
rect 26236 17726 26238 17778
rect 26290 17726 26292 17778
rect 26236 17714 26292 17726
rect 28364 17778 28420 19180
rect 28588 18452 28644 20188
rect 29148 20132 29540 20188
rect 29484 19906 29540 20132
rect 29484 19854 29486 19906
rect 29538 19854 29540 19906
rect 29484 19842 29540 19854
rect 37884 20018 37940 20030
rect 37884 19966 37886 20018
rect 37938 19966 37940 20018
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 37660 19236 37716 19246
rect 37660 19142 37716 19180
rect 37884 19124 37940 19966
rect 40012 19794 40068 19806
rect 40012 19742 40014 19794
rect 40066 19742 40068 19794
rect 40012 19572 40068 19742
rect 40012 19506 40068 19516
rect 37884 19058 37940 19068
rect 40012 19346 40068 19358
rect 40012 19294 40014 19346
rect 40066 19294 40068 19346
rect 37660 19012 37716 19022
rect 28588 18450 29316 18452
rect 28588 18398 28590 18450
rect 28642 18398 29316 18450
rect 28588 18396 29316 18398
rect 28588 18386 28644 18396
rect 28364 17726 28366 17778
rect 28418 17726 28420 17778
rect 28364 17714 28420 17726
rect 29260 17778 29316 18396
rect 37660 18450 37716 18956
rect 40012 18900 40068 19294
rect 40012 18834 40068 18844
rect 37660 18398 37662 18450
rect 37714 18398 37716 18450
rect 37660 18386 37716 18398
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 29260 17726 29262 17778
rect 29314 17726 29316 17778
rect 29260 17714 29316 17726
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 25452 17668 25508 17678
rect 25340 17666 25508 17668
rect 25340 17614 25454 17666
rect 25506 17614 25508 17666
rect 25340 17612 25508 17614
rect 25340 17108 25396 17612
rect 25452 17602 25508 17612
rect 37660 17668 37716 17678
rect 37660 17574 37716 17612
rect 40012 17556 40068 17726
rect 40012 17490 40068 17500
rect 25340 17014 25396 17052
rect 24668 16718 24670 16770
rect 24722 16718 24724 16770
rect 24668 16706 24724 16718
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 20636 15374 20638 15426
rect 20690 15374 20692 15426
rect 20636 15362 20692 15374
rect 21420 15538 21924 15540
rect 21420 15486 21870 15538
rect 21922 15486 21924 15538
rect 21420 15484 21924 15486
rect 21420 15314 21476 15484
rect 21868 15474 21924 15484
rect 21420 15262 21422 15314
rect 21474 15262 21476 15314
rect 21420 15250 21476 15262
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 20412 14644 20468 14654
rect 20300 14642 20468 14644
rect 20300 14590 20414 14642
rect 20466 14590 20468 14642
rect 20300 14588 20468 14590
rect 20412 14578 20468 14588
rect 17500 14478 17502 14530
rect 17554 14478 17556 14530
rect 17500 14466 17556 14478
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 17052 8372 17332 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 17052 3554 17108 8372
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 17052 3502 17054 3554
rect 17106 3502 17108 3554
rect 17052 3490 17108 3502
rect 16828 3444 16884 3454
rect 16828 800 16884 3388
rect 18060 3444 18116 3454
rect 18060 3330 18116 3388
rect 18060 3278 18062 3330
rect 18114 3278 18116 3330
rect 18060 3266 18116 3278
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 16800 0 16912 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4284 27074 4340 27076
rect 4284 27022 4286 27074
rect 4286 27022 4338 27074
rect 4338 27022 4340 27074
rect 4284 27020 4340 27022
rect 15372 27020 15428 27076
rect 16380 26348 16436 26404
rect 1932 26236 1988 26292
rect 4284 26290 4340 26292
rect 4284 26238 4286 26290
rect 4286 26238 4338 26290
rect 4338 26238 4340 26290
rect 4284 26236 4340 26238
rect 12124 26236 12180 26292
rect 14812 26236 14868 26292
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 1932 25564 1988 25620
rect 4284 25506 4340 25508
rect 4284 25454 4286 25506
rect 4286 25454 4338 25506
rect 4338 25454 4340 25506
rect 4284 25452 4340 25454
rect 9996 25452 10052 25508
rect 12796 25506 12852 25508
rect 12796 25454 12798 25506
rect 12798 25454 12850 25506
rect 12850 25454 12852 25506
rect 12796 25452 12852 25454
rect 2044 24892 2100 24948
rect 12572 24610 12628 24612
rect 12572 24558 12574 24610
rect 12574 24558 12626 24610
rect 12626 24558 12628 24610
rect 12572 24556 12628 24558
rect 4476 24330 4532 24332
rect 4284 24220 4340 24276
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 1932 21532 1988 21588
rect 13468 25340 13524 25396
rect 14252 24780 14308 24836
rect 13916 24722 13972 24724
rect 13916 24670 13918 24722
rect 13918 24670 13970 24722
rect 13970 24670 13972 24722
rect 13916 24668 13972 24670
rect 13804 24610 13860 24612
rect 13804 24558 13806 24610
rect 13806 24558 13858 24610
rect 13858 24558 13860 24610
rect 13804 24556 13860 24558
rect 13916 24444 13972 24500
rect 15596 26290 15652 26292
rect 15596 26238 15598 26290
rect 15598 26238 15650 26290
rect 15650 26238 15652 26290
rect 15596 26236 15652 26238
rect 17388 26402 17444 26404
rect 17388 26350 17390 26402
rect 17390 26350 17442 26402
rect 17442 26350 17444 26402
rect 17388 26348 17444 26350
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 24892 38220 24948 38276
rect 26124 38274 26180 38276
rect 26124 38222 26126 38274
rect 26126 38222 26178 38274
rect 26178 38222 26180 38274
rect 26124 38220 26180 38222
rect 20860 37436 20916 37492
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 17612 25676 17668 25732
rect 14924 25452 14980 25508
rect 15596 25506 15652 25508
rect 15596 25454 15598 25506
rect 15598 25454 15650 25506
rect 15650 25454 15652 25506
rect 15596 25452 15652 25454
rect 15484 24834 15540 24836
rect 15484 24782 15486 24834
rect 15486 24782 15538 24834
rect 15538 24782 15540 24834
rect 15484 24780 15540 24782
rect 15708 24780 15764 24836
rect 14700 24444 14756 24500
rect 14140 24332 14196 24388
rect 14028 23884 14084 23940
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4284 22092 4340 22148
rect 4172 21420 4228 21476
rect 9548 21474 9604 21476
rect 9548 21422 9550 21474
rect 9550 21422 9602 21474
rect 9602 21422 9604 21474
rect 9548 21420 9604 21422
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 11788 21532 11844 21588
rect 13020 22540 13076 22596
rect 13692 22540 13748 22596
rect 15596 24668 15652 24724
rect 17724 24668 17780 24724
rect 15148 23042 15204 23044
rect 15148 22990 15150 23042
rect 15150 22990 15202 23042
rect 15202 22990 15204 23042
rect 15148 22988 15204 22990
rect 15820 24332 15876 24388
rect 15820 23548 15876 23604
rect 16604 23436 16660 23492
rect 16044 23212 16100 23268
rect 12460 21586 12516 21588
rect 12460 21534 12462 21586
rect 12462 21534 12514 21586
rect 12514 21534 12516 21586
rect 12460 21532 12516 21534
rect 11564 21308 11620 21364
rect 11116 20802 11172 20804
rect 11116 20750 11118 20802
rect 11118 20750 11170 20802
rect 11170 20750 11172 20802
rect 11116 20748 11172 20750
rect 11452 20524 11508 20580
rect 4284 20018 4340 20020
rect 4284 19966 4286 20018
rect 4286 19966 4338 20018
rect 4338 19966 4340 20018
rect 4284 19964 4340 19966
rect 8876 19964 8932 20020
rect 1932 19794 1988 19796
rect 1932 19742 1934 19794
rect 1934 19742 1986 19794
rect 1986 19742 1988 19794
rect 1932 19740 1988 19742
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 8876 18620 8932 18676
rect 11228 20018 11284 20020
rect 11228 19966 11230 20018
rect 11230 19966 11282 20018
rect 11282 19966 11284 20018
rect 11228 19964 11284 19966
rect 12796 21420 12852 21476
rect 12908 21362 12964 21364
rect 12908 21310 12910 21362
rect 12910 21310 12962 21362
rect 12962 21310 12964 21362
rect 12908 21308 12964 21310
rect 12572 19906 12628 19908
rect 12572 19854 12574 19906
rect 12574 19854 12626 19906
rect 12626 19854 12628 19906
rect 12572 19852 12628 19854
rect 11116 18674 11172 18676
rect 11116 18622 11118 18674
rect 11118 18622 11170 18674
rect 11170 18622 11172 18674
rect 11116 18620 11172 18622
rect 11228 18562 11284 18564
rect 11228 18510 11230 18562
rect 11230 18510 11282 18562
rect 11282 18510 11284 18562
rect 11228 18508 11284 18510
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 1932 17778 1988 17780
rect 1932 17726 1934 17778
rect 1934 17726 1986 17778
rect 1986 17726 1988 17778
rect 1932 17724 1988 17726
rect 4284 17666 4340 17668
rect 4284 17614 4286 17666
rect 4286 17614 4338 17666
rect 4338 17614 4340 17666
rect 4284 17612 4340 17614
rect 9324 17612 9380 17668
rect 13468 20578 13524 20580
rect 13468 20526 13470 20578
rect 13470 20526 13522 20578
rect 13522 20526 13524 20578
rect 13468 20524 13524 20526
rect 13692 19964 13748 20020
rect 13580 19852 13636 19908
rect 13916 20524 13972 20580
rect 14252 20578 14308 20580
rect 14252 20526 14254 20578
rect 14254 20526 14306 20578
rect 14306 20526 14308 20578
rect 14252 20524 14308 20526
rect 16492 23266 16548 23268
rect 16492 23214 16494 23266
rect 16494 23214 16546 23266
rect 16546 23214 16548 23266
rect 16492 23212 16548 23214
rect 16492 22988 16548 23044
rect 16716 22594 16772 22596
rect 16716 22542 16718 22594
rect 16718 22542 16770 22594
rect 16770 22542 16772 22594
rect 16716 22540 16772 22542
rect 17388 22594 17444 22596
rect 17388 22542 17390 22594
rect 17390 22542 17442 22594
rect 17442 22542 17444 22594
rect 17388 22540 17444 22542
rect 16156 21586 16212 21588
rect 16156 21534 16158 21586
rect 16158 21534 16210 21586
rect 16210 21534 16212 21586
rect 16156 21532 16212 21534
rect 15820 20524 15876 20580
rect 14924 20018 14980 20020
rect 14924 19966 14926 20018
rect 14926 19966 14978 20018
rect 14978 19966 14980 20018
rect 14924 19964 14980 19966
rect 14700 19906 14756 19908
rect 14700 19854 14702 19906
rect 14702 19854 14754 19906
rect 14754 19854 14756 19906
rect 14700 19852 14756 19854
rect 13804 19180 13860 19236
rect 14588 19234 14644 19236
rect 14588 19182 14590 19234
rect 14590 19182 14642 19234
rect 14642 19182 14644 19234
rect 14588 19180 14644 19182
rect 12908 18732 12964 18788
rect 12684 18562 12740 18564
rect 12684 18510 12686 18562
rect 12686 18510 12738 18562
rect 12738 18510 12740 18562
rect 12684 18508 12740 18510
rect 13132 18508 13188 18564
rect 11228 16994 11284 16996
rect 11228 16942 11230 16994
rect 11230 16942 11282 16994
rect 11282 16942 11284 16994
rect 11228 16940 11284 16942
rect 1932 16828 1988 16884
rect 4284 16882 4340 16884
rect 4284 16830 4286 16882
rect 4286 16830 4338 16882
rect 4338 16830 4340 16882
rect 4284 16828 4340 16830
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 15708 20076 15764 20132
rect 15148 19740 15204 19796
rect 14476 18396 14532 18452
rect 12460 17612 12516 17668
rect 14476 17666 14532 17668
rect 14476 17614 14478 17666
rect 14478 17614 14530 17666
rect 14530 17614 14532 17666
rect 14476 17612 14532 17614
rect 15596 19122 15652 19124
rect 15596 19070 15598 19122
rect 15598 19070 15650 19122
rect 15650 19070 15652 19122
rect 15596 19068 15652 19070
rect 16268 20636 16324 20692
rect 18620 26290 18676 26292
rect 18620 26238 18622 26290
rect 18622 26238 18674 26290
rect 18674 26238 18676 26290
rect 18620 26236 18676 26238
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19404 26236 19460 26292
rect 18172 25676 18228 25732
rect 18508 25676 18564 25732
rect 19740 25676 19796 25732
rect 22092 37490 22148 37492
rect 22092 37438 22094 37490
rect 22094 37438 22146 37490
rect 22146 37438 22148 37490
rect 22092 37436 22148 37438
rect 40236 36988 40292 37044
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 28476 27804 28532 27860
rect 37660 27858 37716 27860
rect 37660 27806 37662 27858
rect 37662 27806 37714 27858
rect 37714 27806 37716 27858
rect 37660 27804 37716 27806
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 23100 26460 23156 26516
rect 23772 26514 23828 26516
rect 23772 26462 23774 26514
rect 23774 26462 23826 26514
rect 23826 26462 23828 26514
rect 23772 26460 23828 26462
rect 21868 26290 21924 26292
rect 21868 26238 21870 26290
rect 21870 26238 21922 26290
rect 21922 26238 21924 26290
rect 21868 26236 21924 26238
rect 20300 25730 20356 25732
rect 20300 25678 20302 25730
rect 20302 25678 20354 25730
rect 20354 25678 20356 25730
rect 20300 25676 20356 25678
rect 18732 25340 18788 25396
rect 17948 23660 18004 23716
rect 18060 23324 18116 23380
rect 15932 19628 15988 19684
rect 16156 19516 16212 19572
rect 15596 18620 15652 18676
rect 14924 18508 14980 18564
rect 15820 18844 15876 18900
rect 15820 18562 15876 18564
rect 15820 18510 15822 18562
rect 15822 18510 15874 18562
rect 15874 18510 15876 18562
rect 15820 18508 15876 18510
rect 16604 21532 16660 21588
rect 16604 19964 16660 20020
rect 16828 21586 16884 21588
rect 16828 21534 16830 21586
rect 16830 21534 16882 21586
rect 16882 21534 16884 21586
rect 16828 21532 16884 21534
rect 18172 23436 18228 23492
rect 18620 23212 18676 23268
rect 18620 22764 18676 22820
rect 19292 24892 19348 24948
rect 18396 22204 18452 22260
rect 17948 21586 18004 21588
rect 17948 21534 17950 21586
rect 17950 21534 18002 21586
rect 18002 21534 18004 21586
rect 17948 21532 18004 21534
rect 17500 21362 17556 21364
rect 17500 21310 17502 21362
rect 17502 21310 17554 21362
rect 17554 21310 17556 21362
rect 17500 21308 17556 21310
rect 17500 20748 17556 20804
rect 16716 20076 16772 20132
rect 17276 19234 17332 19236
rect 17276 19182 17278 19234
rect 17278 19182 17330 19234
rect 17330 19182 17332 19234
rect 17276 19180 17332 19182
rect 16380 18562 16436 18564
rect 16380 18510 16382 18562
rect 16382 18510 16434 18562
rect 16434 18510 16436 18562
rect 16380 18508 16436 18510
rect 16156 18396 16212 18452
rect 12796 16940 12852 16996
rect 12236 16044 12292 16100
rect 12908 16828 12964 16884
rect 15596 17666 15652 17668
rect 15596 17614 15598 17666
rect 15598 17614 15650 17666
rect 15650 17614 15652 17666
rect 15596 17612 15652 17614
rect 16380 17666 16436 17668
rect 16380 17614 16382 17666
rect 16382 17614 16434 17666
rect 16434 17614 16436 17666
rect 16380 17612 16436 17614
rect 14588 16828 14644 16884
rect 14700 16210 14756 16212
rect 14700 16158 14702 16210
rect 14702 16158 14754 16210
rect 14754 16158 14756 16210
rect 14700 16156 14756 16158
rect 14028 16098 14084 16100
rect 14028 16046 14030 16098
rect 14030 16046 14082 16098
rect 14082 16046 14084 16098
rect 14028 16044 14084 16046
rect 15260 16156 15316 16212
rect 15820 15932 15876 15988
rect 17164 15986 17220 15988
rect 17164 15934 17166 15986
rect 17166 15934 17218 15986
rect 17218 15934 17220 15986
rect 17164 15932 17220 15934
rect 14028 15260 14084 15316
rect 15820 15314 15876 15316
rect 15820 15262 15822 15314
rect 15822 15262 15874 15314
rect 15874 15262 15876 15314
rect 15820 15260 15876 15262
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 17500 20130 17556 20132
rect 17500 20078 17502 20130
rect 17502 20078 17554 20130
rect 17554 20078 17556 20130
rect 17500 20076 17556 20078
rect 17500 19516 17556 19572
rect 17612 20018 17668 20020
rect 17612 19966 17614 20018
rect 17614 19966 17666 20018
rect 17666 19966 17668 20018
rect 17612 19964 17668 19966
rect 17836 19964 17892 20020
rect 17836 19628 17892 19684
rect 19404 23772 19460 23828
rect 18620 21532 18676 21588
rect 18396 21308 18452 21364
rect 17948 19740 18004 19796
rect 18620 20524 18676 20580
rect 18060 19516 18116 19572
rect 18060 18844 18116 18900
rect 18284 18732 18340 18788
rect 19068 23548 19124 23604
rect 18844 21698 18900 21700
rect 18844 21646 18846 21698
rect 18846 21646 18898 21698
rect 18898 21646 18900 21698
rect 18844 21644 18900 21646
rect 18956 21532 19012 21588
rect 18844 20636 18900 20692
rect 18844 19852 18900 19908
rect 19180 20188 19236 20244
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20524 25116 20580 25172
rect 20044 25060 20100 25062
rect 20412 24946 20468 24948
rect 20412 24894 20414 24946
rect 20414 24894 20466 24946
rect 20466 24894 20468 24946
rect 20412 24892 20468 24894
rect 21308 25394 21364 25396
rect 21308 25342 21310 25394
rect 21310 25342 21362 25394
rect 21362 25342 21364 25394
rect 21308 25340 21364 25342
rect 21644 25394 21700 25396
rect 21644 25342 21646 25394
rect 21646 25342 21698 25394
rect 21698 25342 21700 25394
rect 21644 25340 21700 25342
rect 20748 25228 20804 25284
rect 19628 23884 19684 23940
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19740 23378 19796 23380
rect 19740 23326 19742 23378
rect 19742 23326 19794 23378
rect 19794 23326 19796 23378
rect 19740 23324 19796 23326
rect 19964 23378 20020 23380
rect 19964 23326 19966 23378
rect 19966 23326 20018 23378
rect 20018 23326 20020 23378
rect 19964 23324 20020 23326
rect 19628 22764 19684 22820
rect 19404 22146 19460 22148
rect 19404 22094 19406 22146
rect 19406 22094 19458 22146
rect 19458 22094 19460 22146
rect 19404 22092 19460 22094
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20076 21644 20132 21700
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20076 20242 20132 20244
rect 20076 20190 20078 20242
rect 20078 20190 20130 20242
rect 20130 20190 20132 20242
rect 20076 20188 20132 20190
rect 19516 20076 19572 20132
rect 18956 19404 19012 19460
rect 19068 20018 19124 20020
rect 19068 19966 19070 20018
rect 19070 19966 19122 20018
rect 19122 19966 19124 20018
rect 19068 19964 19124 19966
rect 18956 19180 19012 19236
rect 18732 18508 18788 18564
rect 18620 17666 18676 17668
rect 18620 17614 18622 17666
rect 18622 17614 18674 17666
rect 18674 17614 18676 17666
rect 18620 17612 18676 17614
rect 19740 20130 19796 20132
rect 19740 20078 19742 20130
rect 19742 20078 19794 20130
rect 19794 20078 19796 20130
rect 19740 20076 19796 20078
rect 19628 19516 19684 19572
rect 20300 20188 20356 20244
rect 21644 24780 21700 24836
rect 20860 23378 20916 23380
rect 20860 23326 20862 23378
rect 20862 23326 20914 23378
rect 20914 23326 20916 23378
rect 20860 23324 20916 23326
rect 20748 20130 20804 20132
rect 20748 20078 20750 20130
rect 20750 20078 20802 20130
rect 20802 20078 20804 20130
rect 20748 20076 20804 20078
rect 20412 19964 20468 20020
rect 20636 19404 20692 19460
rect 19852 19068 19908 19124
rect 19180 18956 19236 19012
rect 18956 18674 19012 18676
rect 18956 18622 18958 18674
rect 18958 18622 19010 18674
rect 19010 18622 19012 18674
rect 18956 18620 19012 18622
rect 20076 18956 20132 19012
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20636 18844 20692 18900
rect 21532 23154 21588 23156
rect 21532 23102 21534 23154
rect 21534 23102 21586 23154
rect 21586 23102 21588 23154
rect 21532 23100 21588 23102
rect 21420 22764 21476 22820
rect 21308 22146 21364 22148
rect 21308 22094 21310 22146
rect 21310 22094 21362 22146
rect 21362 22094 21364 22146
rect 21308 22092 21364 22094
rect 22092 25676 22148 25732
rect 24444 25506 24500 25508
rect 24444 25454 24446 25506
rect 24446 25454 24498 25506
rect 24498 25454 24500 25506
rect 24444 25452 24500 25454
rect 25116 25452 25172 25508
rect 27020 27020 27076 27076
rect 25452 26908 25508 26964
rect 26236 26012 26292 26068
rect 23996 25394 24052 25396
rect 23996 25342 23998 25394
rect 23998 25342 24050 25394
rect 24050 25342 24052 25394
rect 23996 25340 24052 25342
rect 23772 25116 23828 25172
rect 23548 24722 23604 24724
rect 23548 24670 23550 24722
rect 23550 24670 23602 24722
rect 23602 24670 23604 24722
rect 23548 24668 23604 24670
rect 21756 23826 21812 23828
rect 21756 23774 21758 23826
rect 21758 23774 21810 23826
rect 21810 23774 21812 23826
rect 21756 23772 21812 23774
rect 22764 23884 22820 23940
rect 22092 23660 22148 23716
rect 21868 23436 21924 23492
rect 21532 21532 21588 21588
rect 21308 20188 21364 20244
rect 23660 23826 23716 23828
rect 23660 23774 23662 23826
rect 23662 23774 23714 23826
rect 23714 23774 23716 23826
rect 23660 23772 23716 23774
rect 23324 23714 23380 23716
rect 23324 23662 23326 23714
rect 23326 23662 23378 23714
rect 23378 23662 23380 23714
rect 23324 23660 23380 23662
rect 22764 22092 22820 22148
rect 24332 25116 24388 25172
rect 25676 24780 25732 24836
rect 24892 23436 24948 23492
rect 25452 23436 25508 23492
rect 24668 23100 24724 23156
rect 25564 23884 25620 23940
rect 28028 27020 28084 27076
rect 27020 26066 27076 26068
rect 27020 26014 27022 26066
rect 27022 26014 27074 26066
rect 27074 26014 27076 26066
rect 27020 26012 27076 26014
rect 29260 26962 29316 26964
rect 29260 26910 29262 26962
rect 29262 26910 29314 26962
rect 29314 26910 29316 26962
rect 29260 26908 29316 26910
rect 39900 26908 39956 26964
rect 37660 26460 37716 26516
rect 28252 26402 28308 26404
rect 28252 26350 28254 26402
rect 28254 26350 28306 26402
rect 28306 26350 28308 26402
rect 28252 26348 28308 26350
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 27244 25116 27300 25172
rect 27020 24834 27076 24836
rect 27020 24782 27022 24834
rect 27022 24782 27074 24834
rect 27074 24782 27076 24834
rect 27020 24780 27076 24782
rect 27692 25564 27748 25620
rect 28588 25618 28644 25620
rect 28588 25566 28590 25618
rect 28590 25566 28642 25618
rect 28642 25566 28644 25618
rect 28588 25564 28644 25566
rect 29260 25564 29316 25620
rect 37660 25506 37716 25508
rect 37660 25454 37662 25506
rect 37662 25454 37714 25506
rect 37714 25454 37716 25506
rect 37660 25452 37716 25454
rect 29484 25282 29540 25284
rect 29484 25230 29486 25282
rect 29486 25230 29538 25282
rect 29538 25230 29540 25282
rect 29484 25228 29540 25230
rect 40012 26236 40068 26292
rect 39900 25564 39956 25620
rect 37884 25228 37940 25284
rect 40012 24892 40068 24948
rect 26012 23884 26068 23940
rect 25676 23772 25732 23828
rect 22316 21698 22372 21700
rect 22316 21646 22318 21698
rect 22318 21646 22370 21698
rect 22370 21646 22372 21698
rect 22316 21644 22372 21646
rect 22540 21868 22596 21924
rect 21756 20748 21812 20804
rect 23324 21868 23380 21924
rect 22204 20690 22260 20692
rect 22204 20638 22206 20690
rect 22206 20638 22258 20690
rect 22258 20638 22260 20690
rect 22204 20636 22260 20638
rect 21868 20524 21924 20580
rect 22988 21756 23044 21812
rect 22988 20802 23044 20804
rect 22988 20750 22990 20802
rect 22990 20750 23042 20802
rect 23042 20750 23044 20802
rect 22988 20748 23044 20750
rect 23100 20524 23156 20580
rect 23212 19964 23268 20020
rect 21084 19180 21140 19236
rect 20972 19068 21028 19124
rect 20972 18732 21028 18788
rect 21644 18956 21700 19012
rect 21420 18732 21476 18788
rect 20300 17948 20356 18004
rect 21420 17948 21476 18004
rect 21308 17890 21364 17892
rect 21308 17838 21310 17890
rect 21310 17838 21362 17890
rect 21362 17838 21364 17890
rect 21308 17836 21364 17838
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19740 16882 19796 16884
rect 19740 16830 19742 16882
rect 19742 16830 19794 16882
rect 19794 16830 19796 16882
rect 19740 16828 19796 16830
rect 17388 15260 17444 15316
rect 20300 16882 20356 16884
rect 20300 16830 20302 16882
rect 20302 16830 20354 16882
rect 20354 16830 20356 16882
rect 20300 16828 20356 16830
rect 21308 16828 21364 16884
rect 21644 18620 21700 18676
rect 22876 18620 22932 18676
rect 21868 17948 21924 18004
rect 21644 17890 21700 17892
rect 21644 17838 21646 17890
rect 21646 17838 21698 17890
rect 21698 17838 21700 17890
rect 21644 17836 21700 17838
rect 22540 18172 22596 18228
rect 22764 17836 22820 17892
rect 23660 19122 23716 19124
rect 23660 19070 23662 19122
rect 23662 19070 23714 19122
rect 23714 19070 23716 19122
rect 23660 19068 23716 19070
rect 23772 19010 23828 19012
rect 23772 18958 23774 19010
rect 23774 18958 23826 19010
rect 23826 18958 23828 19010
rect 23772 18956 23828 18958
rect 23436 18620 23492 18676
rect 23548 18562 23604 18564
rect 23548 18510 23550 18562
rect 23550 18510 23602 18562
rect 23602 18510 23604 18562
rect 23548 18508 23604 18510
rect 23436 18226 23492 18228
rect 23436 18174 23438 18226
rect 23438 18174 23490 18226
rect 23490 18174 23492 18226
rect 23436 18172 23492 18174
rect 24444 20076 24500 20132
rect 25676 21756 25732 21812
rect 25788 23266 25844 23268
rect 25788 23214 25790 23266
rect 25790 23214 25842 23266
rect 25842 23214 25844 23266
rect 25788 23212 25844 23214
rect 27020 23266 27076 23268
rect 27020 23214 27022 23266
rect 27022 23214 27074 23266
rect 27074 23214 27076 23266
rect 27020 23212 27076 23214
rect 29148 24668 29204 24724
rect 27692 23714 27748 23716
rect 27692 23662 27694 23714
rect 27694 23662 27746 23714
rect 27746 23662 27748 23714
rect 27692 23660 27748 23662
rect 28252 23266 28308 23268
rect 28252 23214 28254 23266
rect 28254 23214 28306 23266
rect 28306 23214 28308 23266
rect 28252 23212 28308 23214
rect 25788 21868 25844 21924
rect 25452 21308 25508 21364
rect 25340 20690 25396 20692
rect 25340 20638 25342 20690
rect 25342 20638 25394 20690
rect 25394 20638 25396 20690
rect 25340 20636 25396 20638
rect 25788 21084 25844 21140
rect 26012 22204 26068 22260
rect 25564 20188 25620 20244
rect 25004 19346 25060 19348
rect 25004 19294 25006 19346
rect 25006 19294 25058 19346
rect 25058 19294 25060 19346
rect 25004 19292 25060 19294
rect 24892 19234 24948 19236
rect 24892 19182 24894 19234
rect 24894 19182 24946 19234
rect 24946 19182 24948 19234
rect 24892 19180 24948 19182
rect 25004 19010 25060 19012
rect 25004 18958 25006 19010
rect 25006 18958 25058 19010
rect 25058 18958 25060 19010
rect 25004 18956 25060 18958
rect 24556 18844 24612 18900
rect 24668 18732 24724 18788
rect 25788 20524 25844 20580
rect 25452 19292 25508 19348
rect 26236 20242 26292 20244
rect 26236 20190 26238 20242
rect 26238 20190 26290 20242
rect 26290 20190 26292 20242
rect 26236 20188 26292 20190
rect 26572 20188 26628 20244
rect 37660 24722 37716 24724
rect 37660 24670 37662 24722
rect 37662 24670 37714 24722
rect 37714 24670 37716 24722
rect 37660 24668 37716 24670
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 40012 24220 40068 24276
rect 29148 23660 29204 23716
rect 29372 23266 29428 23268
rect 29372 23214 29374 23266
rect 29374 23214 29426 23266
rect 29426 23214 29428 23266
rect 29372 23212 29428 23214
rect 28028 21308 28084 21364
rect 28476 21308 28532 21364
rect 28588 20188 28644 20244
rect 40012 23548 40068 23604
rect 37660 23154 37716 23156
rect 37660 23102 37662 23154
rect 37662 23102 37714 23154
rect 37714 23102 37716 23154
rect 37660 23100 37716 23102
rect 37436 22876 37492 22932
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 37660 22764 37716 22820
rect 40012 22204 40068 22260
rect 37660 21586 37716 21588
rect 37660 21534 37662 21586
rect 37662 21534 37714 21586
rect 37714 21534 37716 21586
rect 37660 21532 37716 21534
rect 40012 21532 40068 21588
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 28364 19180 28420 19236
rect 27244 19068 27300 19124
rect 28140 19068 28196 19124
rect 27468 19010 27524 19012
rect 27468 18958 27470 19010
rect 27470 18958 27522 19010
rect 27522 18958 27524 19010
rect 27468 18956 27524 18958
rect 26012 18732 26068 18788
rect 24220 18338 24276 18340
rect 24220 18286 24222 18338
rect 24222 18286 24274 18338
rect 24274 18286 24276 18338
rect 24220 18284 24276 18286
rect 23772 17612 23828 17668
rect 24668 17612 24724 17668
rect 18508 15202 18564 15204
rect 18508 15150 18510 15202
rect 18510 15150 18562 15202
rect 18562 15150 18564 15202
rect 18508 15148 18564 15150
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19628 15148 19684 15204
rect 21868 17052 21924 17108
rect 26012 18338 26068 18340
rect 26012 18286 26014 18338
rect 26014 18286 26066 18338
rect 26066 18286 26068 18338
rect 26012 18284 26068 18286
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 37660 19234 37716 19236
rect 37660 19182 37662 19234
rect 37662 19182 37714 19234
rect 37714 19182 37716 19234
rect 37660 19180 37716 19182
rect 40012 19516 40068 19572
rect 37884 19068 37940 19124
rect 37660 18956 37716 19012
rect 40012 18844 40068 18900
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 37660 17666 37716 17668
rect 37660 17614 37662 17666
rect 37662 17614 37714 17666
rect 37714 17614 37716 17666
rect 37660 17612 37716 17614
rect 40012 17500 40068 17556
rect 25340 17106 25396 17108
rect 25340 17054 25342 17106
rect 25342 17054 25394 17106
rect 25394 17054 25396 17106
rect 25340 17052 25396 17054
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 16828 3388 16884 3444
rect 18060 3388 18116 3444
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 24882 38220 24892 38276
rect 24948 38220 26124 38276
rect 26180 38220 26190 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 20850 37436 20860 37492
rect 20916 37436 22092 37492
rect 22148 37436 22158 37492
rect 41200 37044 42000 37072
rect 40226 36988 40236 37044
rect 40292 36988 42000 37044
rect 41200 36960 42000 36988
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 28466 27804 28476 27860
rect 28532 27804 37660 27860
rect 37716 27804 37726 27860
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 4274 27020 4284 27076
rect 4340 27020 15372 27076
rect 15428 27020 15438 27076
rect 27010 27020 27020 27076
rect 27076 27020 28028 27076
rect 28084 27020 28094 27076
rect 41200 26964 42000 26992
rect 25442 26908 25452 26964
rect 25508 26908 29260 26964
rect 29316 26908 29326 26964
rect 39890 26908 39900 26964
rect 39956 26908 42000 26964
rect 41200 26880 42000 26908
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 23090 26460 23100 26516
rect 23156 26460 23772 26516
rect 23828 26460 23838 26516
rect 31892 26460 37660 26516
rect 37716 26460 37726 26516
rect 31892 26404 31948 26460
rect 16370 26348 16380 26404
rect 16436 26348 17388 26404
rect 17444 26348 17454 26404
rect 28242 26348 28252 26404
rect 28308 26348 31948 26404
rect 0 26292 800 26320
rect 41200 26292 42000 26320
rect 0 26236 1932 26292
rect 1988 26236 1998 26292
rect 4274 26236 4284 26292
rect 4340 26236 12124 26292
rect 12180 26236 14812 26292
rect 14868 26236 15596 26292
rect 15652 26236 15662 26292
rect 18610 26236 18620 26292
rect 18676 26236 19404 26292
rect 19460 26236 21868 26292
rect 21924 26236 21934 26292
rect 40002 26236 40012 26292
rect 40068 26236 42000 26292
rect 0 26208 800 26236
rect 41200 26208 42000 26236
rect 26226 26012 26236 26068
rect 26292 26012 27020 26068
rect 27076 26012 27086 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 17602 25676 17612 25732
rect 17668 25676 18172 25732
rect 18228 25676 18508 25732
rect 18564 25676 18574 25732
rect 19730 25676 19740 25732
rect 19796 25676 20300 25732
rect 20356 25676 22092 25732
rect 22148 25676 22158 25732
rect 0 25620 800 25648
rect 41200 25620 42000 25648
rect 0 25564 1932 25620
rect 1988 25564 1998 25620
rect 27682 25564 27692 25620
rect 27748 25564 28588 25620
rect 28644 25564 29260 25620
rect 29316 25564 31948 25620
rect 39890 25564 39900 25620
rect 39956 25564 42000 25620
rect 0 25536 800 25564
rect 31892 25508 31948 25564
rect 41200 25536 42000 25564
rect 4274 25452 4284 25508
rect 4340 25452 9996 25508
rect 10052 25452 10062 25508
rect 12786 25452 12796 25508
rect 12852 25452 14924 25508
rect 14980 25452 15596 25508
rect 15652 25452 15662 25508
rect 24434 25452 24444 25508
rect 24500 25452 25116 25508
rect 25172 25452 25182 25508
rect 31892 25452 37660 25508
rect 37716 25452 37726 25508
rect 9996 25396 10052 25452
rect 9996 25340 13468 25396
rect 13524 25340 13534 25396
rect 18722 25340 18732 25396
rect 18788 25340 21308 25396
rect 21364 25340 21374 25396
rect 21634 25340 21644 25396
rect 21700 25340 23996 25396
rect 24052 25340 24062 25396
rect 21644 25284 21700 25340
rect 20738 25228 20748 25284
rect 20804 25228 21700 25284
rect 29474 25228 29484 25284
rect 29540 25228 37884 25284
rect 37940 25228 37950 25284
rect 20514 25116 20524 25172
rect 20580 25116 20692 25172
rect 23762 25116 23772 25172
rect 23828 25116 24332 25172
rect 24388 25116 27244 25172
rect 27300 25116 27310 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 0 24948 800 24976
rect 0 24892 2044 24948
rect 2100 24892 2110 24948
rect 19282 24892 19292 24948
rect 19348 24892 20412 24948
rect 20468 24892 20478 24948
rect 0 24864 800 24892
rect 20636 24836 20692 25116
rect 41200 24948 42000 24976
rect 40002 24892 40012 24948
rect 40068 24892 42000 24948
rect 41200 24864 42000 24892
rect 14242 24780 14252 24836
rect 14308 24780 15484 24836
rect 15540 24780 15550 24836
rect 15698 24780 15708 24836
rect 15764 24780 21644 24836
rect 21700 24780 21710 24836
rect 25666 24780 25676 24836
rect 25732 24780 27020 24836
rect 27076 24780 27086 24836
rect 13906 24668 13916 24724
rect 13972 24668 15596 24724
rect 15652 24668 15662 24724
rect 17714 24668 17724 24724
rect 17780 24668 23548 24724
rect 23604 24668 23614 24724
rect 29138 24668 29148 24724
rect 29204 24668 37660 24724
rect 37716 24668 37726 24724
rect 17724 24612 17780 24668
rect 12562 24556 12572 24612
rect 12628 24556 13804 24612
rect 13860 24556 13870 24612
rect 15092 24556 17780 24612
rect 15092 24500 15148 24556
rect 13906 24444 13916 24500
rect 13972 24444 14700 24500
rect 14756 24444 15148 24500
rect 14130 24332 14140 24388
rect 14196 24332 15820 24388
rect 15876 24332 15886 24388
rect 0 24276 800 24304
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 41200 24276 42000 24304
rect 0 24220 4284 24276
rect 4340 24220 4350 24276
rect 40002 24220 40012 24276
rect 40068 24220 42000 24276
rect 0 24192 800 24220
rect 41200 24192 42000 24220
rect 14018 23884 14028 23940
rect 14084 23884 19628 23940
rect 19684 23884 22764 23940
rect 22820 23884 25564 23940
rect 25620 23884 26012 23940
rect 26068 23884 26078 23940
rect 19394 23772 19404 23828
rect 19460 23772 21756 23828
rect 21812 23772 21822 23828
rect 23650 23772 23660 23828
rect 23716 23772 25676 23828
rect 25732 23772 25742 23828
rect 17938 23660 17948 23716
rect 18004 23660 22092 23716
rect 22148 23660 23324 23716
rect 23380 23660 23390 23716
rect 27682 23660 27692 23716
rect 27748 23660 29148 23716
rect 29204 23660 29214 23716
rect 41200 23604 42000 23632
rect 15810 23548 15820 23604
rect 15876 23548 19068 23604
rect 19124 23548 19134 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 41200 23520 42000 23548
rect 16594 23436 16604 23492
rect 16660 23436 18172 23492
rect 18228 23436 18238 23492
rect 21858 23436 21868 23492
rect 21924 23436 24892 23492
rect 24948 23436 25452 23492
rect 25508 23436 25518 23492
rect 18050 23324 18060 23380
rect 18116 23324 19740 23380
rect 19796 23324 19806 23380
rect 19954 23324 19964 23380
rect 20020 23324 20860 23380
rect 20916 23324 20926 23380
rect 16034 23212 16044 23268
rect 16100 23212 16492 23268
rect 16548 23212 18620 23268
rect 18676 23212 18686 23268
rect 25778 23212 25788 23268
rect 25844 23212 27020 23268
rect 27076 23212 27086 23268
rect 28242 23212 28252 23268
rect 28308 23212 28318 23268
rect 29362 23212 29372 23268
rect 29428 23212 37716 23268
rect 28252 23156 28308 23212
rect 37660 23156 37716 23212
rect 21522 23100 21532 23156
rect 21588 23100 24668 23156
rect 24724 23100 26908 23156
rect 28252 23100 32564 23156
rect 37650 23100 37660 23156
rect 37716 23100 37726 23156
rect 26852 23044 26908 23100
rect 32508 23044 32564 23100
rect 15138 22988 15148 23044
rect 15204 22988 16492 23044
rect 16548 22988 16558 23044
rect 26852 22988 31948 23044
rect 32508 22988 37716 23044
rect 31892 22932 31948 22988
rect 31892 22876 37436 22932
rect 37492 22876 37502 22932
rect 37660 22820 37716 22988
rect 41200 22932 42000 22960
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 41200 22848 42000 22876
rect 18610 22764 18620 22820
rect 18676 22764 19628 22820
rect 19684 22764 21420 22820
rect 21476 22764 21486 22820
rect 37650 22764 37660 22820
rect 37716 22764 37726 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 13010 22540 13020 22596
rect 13076 22540 13692 22596
rect 13748 22540 13758 22596
rect 16706 22540 16716 22596
rect 16772 22540 17388 22596
rect 17444 22540 17454 22596
rect 41200 22260 42000 22288
rect 18386 22204 18396 22260
rect 18452 22204 26012 22260
rect 26068 22204 26078 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 41200 22176 42000 22204
rect 4274 22092 4284 22148
rect 4340 22092 19404 22148
rect 19460 22092 19470 22148
rect 21298 22092 21308 22148
rect 21364 22092 22764 22148
rect 22820 22092 22830 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 22530 21868 22540 21924
rect 22596 21868 23324 21924
rect 23380 21868 25788 21924
rect 25844 21868 25854 21924
rect 22978 21756 22988 21812
rect 23044 21756 25676 21812
rect 25732 21756 25742 21812
rect 16604 21644 18844 21700
rect 18900 21644 18910 21700
rect 20066 21644 20076 21700
rect 20132 21644 22316 21700
rect 22372 21644 22382 21700
rect 0 21588 800 21616
rect 16604 21588 16660 21644
rect 41200 21588 42000 21616
rect 0 21532 1932 21588
rect 1988 21532 1998 21588
rect 11778 21532 11788 21588
rect 11844 21532 12460 21588
rect 12516 21532 12526 21588
rect 16146 21532 16156 21588
rect 16212 21532 16604 21588
rect 16660 21532 16670 21588
rect 16818 21532 16828 21588
rect 16884 21532 17948 21588
rect 18004 21532 18620 21588
rect 18676 21532 18686 21588
rect 18946 21532 18956 21588
rect 19012 21532 21532 21588
rect 21588 21532 21598 21588
rect 31892 21532 37660 21588
rect 37716 21532 37726 21588
rect 40002 21532 40012 21588
rect 40068 21532 42000 21588
rect 0 21504 800 21532
rect 4162 21420 4172 21476
rect 4228 21420 9548 21476
rect 9604 21420 12796 21476
rect 12852 21420 12862 21476
rect 31892 21364 31948 21532
rect 41200 21504 42000 21532
rect 11554 21308 11564 21364
rect 11620 21308 12908 21364
rect 12964 21308 12974 21364
rect 17490 21308 17500 21364
rect 17556 21308 18396 21364
rect 18452 21308 18462 21364
rect 25442 21308 25452 21364
rect 25508 21308 28028 21364
rect 28084 21308 28476 21364
rect 28532 21308 31948 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 25778 21084 25788 21140
rect 25844 21084 25854 21140
rect 11106 20748 11116 20804
rect 11172 20748 17500 20804
rect 17556 20748 17566 20804
rect 21746 20748 21756 20804
rect 21812 20748 22988 20804
rect 23044 20748 23054 20804
rect 16258 20636 16268 20692
rect 16324 20636 18844 20692
rect 18900 20636 22204 20692
rect 22260 20636 25340 20692
rect 25396 20636 25406 20692
rect 25788 20580 25844 21084
rect 11442 20524 11452 20580
rect 11508 20524 13468 20580
rect 13524 20524 13916 20580
rect 13972 20524 13982 20580
rect 14242 20524 14252 20580
rect 14308 20524 15820 20580
rect 15876 20524 15886 20580
rect 18610 20524 18620 20580
rect 18676 20524 21868 20580
rect 21924 20524 23100 20580
rect 23156 20524 23166 20580
rect 25778 20524 25788 20580
rect 25844 20524 25854 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 19170 20188 19180 20244
rect 19236 20188 20076 20244
rect 20132 20188 20300 20244
rect 20356 20188 21308 20244
rect 21364 20188 21374 20244
rect 25554 20188 25564 20244
rect 25620 20188 26236 20244
rect 26292 20188 26572 20244
rect 26628 20188 28588 20244
rect 28644 20188 28654 20244
rect 15092 20076 15708 20132
rect 15764 20076 16716 20132
rect 16772 20076 16782 20132
rect 17490 20076 17500 20132
rect 17556 20076 19516 20132
rect 19572 20076 19582 20132
rect 19730 20076 19740 20132
rect 19796 20076 20748 20132
rect 20804 20076 24444 20132
rect 24500 20076 24510 20132
rect 4274 19964 4284 20020
rect 4340 19964 8876 20020
rect 8932 19964 8942 20020
rect 11218 19964 11228 20020
rect 11284 19964 13692 20020
rect 13748 19964 14924 20020
rect 14980 19964 14990 20020
rect 15092 19908 15148 20076
rect 16594 19964 16604 20020
rect 16660 19964 17612 20020
rect 17668 19964 17678 20020
rect 17826 19964 17836 20020
rect 17892 19964 19068 20020
rect 19124 19964 19134 20020
rect 20402 19964 20412 20020
rect 20468 19964 23212 20020
rect 23268 19964 23278 20020
rect 20412 19908 20468 19964
rect 12562 19852 12572 19908
rect 12628 19852 13580 19908
rect 13636 19852 13646 19908
rect 14690 19852 14700 19908
rect 14756 19852 15148 19908
rect 18834 19852 18844 19908
rect 18900 19852 20468 19908
rect 1922 19740 1932 19796
rect 1988 19740 1998 19796
rect 15138 19740 15148 19796
rect 15204 19740 17948 19796
rect 18004 19740 18014 19796
rect 0 19572 800 19600
rect 1932 19572 1988 19740
rect 15922 19628 15932 19684
rect 15988 19628 17836 19684
rect 17892 19628 17902 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 0 19516 1988 19572
rect 16146 19516 16156 19572
rect 16212 19516 17500 19572
rect 17556 19516 17566 19572
rect 18050 19516 18060 19572
rect 18116 19516 19628 19572
rect 19684 19516 21308 19572
rect 21364 19516 21374 19572
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 0 19488 800 19516
rect 41200 19488 42000 19516
rect 18946 19404 18956 19460
rect 19012 19404 20636 19460
rect 20692 19404 20702 19460
rect 24994 19292 25004 19348
rect 25060 19292 25452 19348
rect 25508 19292 25518 19348
rect 13794 19180 13804 19236
rect 13860 19180 14588 19236
rect 14644 19180 15148 19236
rect 17266 19180 17276 19236
rect 17332 19180 18956 19236
rect 19012 19180 21084 19236
rect 21140 19180 21150 19236
rect 24882 19180 24892 19236
rect 24948 19180 28364 19236
rect 28420 19180 37660 19236
rect 37716 19180 37726 19236
rect 15092 19124 15148 19180
rect 15092 19068 15596 19124
rect 15652 19068 15662 19124
rect 19842 19068 19852 19124
rect 19908 19068 20972 19124
rect 21028 19068 21038 19124
rect 23650 19068 23660 19124
rect 23716 19068 27244 19124
rect 27300 19068 28140 19124
rect 28196 19068 37884 19124
rect 37940 19068 37950 19124
rect 19170 18956 19180 19012
rect 19236 18956 20076 19012
rect 20132 18956 21644 19012
rect 21700 18956 21710 19012
rect 23762 18956 23772 19012
rect 23828 18956 25004 19012
rect 25060 18956 25070 19012
rect 27458 18956 27468 19012
rect 27524 18956 37660 19012
rect 37716 18956 37726 19012
rect 41200 18900 42000 18928
rect 15810 18844 15820 18900
rect 15876 18844 18060 18900
rect 18116 18844 18126 18900
rect 20626 18844 20636 18900
rect 20692 18844 24556 18900
rect 24612 18844 24622 18900
rect 40002 18844 40012 18900
rect 40068 18844 42000 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 41200 18816 42000 18844
rect 12898 18732 12908 18788
rect 12964 18732 18284 18788
rect 18340 18732 19684 18788
rect 20962 18732 20972 18788
rect 21028 18732 21420 18788
rect 21476 18732 21486 18788
rect 24658 18732 24668 18788
rect 24724 18732 26012 18788
rect 26068 18732 26078 18788
rect 19628 18676 19684 18732
rect 8866 18620 8876 18676
rect 8932 18620 11116 18676
rect 11172 18620 11182 18676
rect 15586 18620 15596 18676
rect 15652 18620 18956 18676
rect 19012 18620 19022 18676
rect 19628 18620 21644 18676
rect 21700 18620 22876 18676
rect 22932 18620 23436 18676
rect 23492 18620 23502 18676
rect 11218 18508 11228 18564
rect 11284 18508 12684 18564
rect 12740 18508 12750 18564
rect 13122 18508 13132 18564
rect 13188 18508 14924 18564
rect 14980 18508 15820 18564
rect 15876 18508 15886 18564
rect 16370 18508 16380 18564
rect 16436 18508 18732 18564
rect 18788 18508 23548 18564
rect 23604 18508 23614 18564
rect 14466 18396 14476 18452
rect 14532 18396 16156 18452
rect 16212 18396 16222 18452
rect 24210 18284 24220 18340
rect 24276 18284 26012 18340
rect 26068 18284 26078 18340
rect 41200 18228 42000 18256
rect 22530 18172 22540 18228
rect 22596 18172 23436 18228
rect 23492 18172 23502 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 41200 18144 42000 18172
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 20290 17948 20300 18004
rect 20356 17948 21420 18004
rect 21476 17948 21868 18004
rect 21924 17948 21934 18004
rect 21270 17836 21308 17892
rect 21364 17836 21374 17892
rect 21634 17836 21644 17892
rect 21700 17836 22764 17892
rect 22820 17836 22830 17892
rect 1922 17724 1932 17780
rect 1988 17724 1998 17780
rect 0 17556 800 17584
rect 1932 17556 1988 17724
rect 4274 17612 4284 17668
rect 4340 17612 9324 17668
rect 9380 17612 12460 17668
rect 12516 17612 12526 17668
rect 14466 17612 14476 17668
rect 14532 17612 15596 17668
rect 15652 17612 15662 17668
rect 16370 17612 16380 17668
rect 16436 17612 18620 17668
rect 18676 17612 18686 17668
rect 23762 17612 23772 17668
rect 23828 17612 24668 17668
rect 24724 17612 37660 17668
rect 37716 17612 37726 17668
rect 41200 17556 42000 17584
rect 0 17500 1988 17556
rect 40002 17500 40012 17556
rect 40068 17500 42000 17556
rect 0 17472 800 17500
rect 41200 17472 42000 17500
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 21858 17052 21868 17108
rect 21924 17052 25340 17108
rect 25396 17052 25406 17108
rect 11218 16940 11228 16996
rect 11284 16940 12796 16996
rect 12852 16940 12862 16996
rect 0 16884 800 16912
rect 0 16828 1932 16884
rect 1988 16828 1998 16884
rect 4274 16828 4284 16884
rect 4340 16828 12908 16884
rect 12964 16828 14588 16884
rect 14644 16828 14654 16884
rect 19730 16828 19740 16884
rect 19796 16828 20300 16884
rect 20356 16828 21308 16884
rect 21364 16828 21374 16884
rect 0 16800 800 16828
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 14690 16156 14700 16212
rect 14756 16156 15260 16212
rect 15316 16156 15326 16212
rect 12226 16044 12236 16100
rect 12292 16044 14028 16100
rect 14084 16044 14094 16100
rect 15810 15932 15820 15988
rect 15876 15932 17164 15988
rect 17220 15932 17230 15988
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 14018 15260 14028 15316
rect 14084 15260 15820 15316
rect 15876 15260 17388 15316
rect 17444 15260 17454 15316
rect 18498 15148 18508 15204
rect 18564 15148 19628 15204
rect 19684 15148 19694 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 16818 3388 16828 3444
rect 16884 3388 18060 3444
rect 18116 3388 18126 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 21308 19516 21364 19572
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 21308 17836 21364 17892
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 21308 19572 21364 19582
rect 21308 17892 21364 19516
rect 21308 17826 21364 17836
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _094_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16128 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _095_
timestamp 1698175906
transform -1 0 16352 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _096_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19936 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _097_
timestamp 1698175906
transform 1 0 19600 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _098_
timestamp 1698175906
transform 1 0 20944 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _099_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19488 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _101_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18704 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15456 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _103_
timestamp 1698175906
transform 1 0 15456 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_
timestamp 1698175906
transform -1 0 19376 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1698175906
transform -1 0 16464 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _107_
timestamp 1698175906
transform -1 0 17024 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16352 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _109_
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22064 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15232 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _112_
timestamp 1698175906
transform 1 0 14672 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _113_
timestamp 1698175906
transform -1 0 20608 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19264 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform -1 0 14000 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _116_
timestamp 1698175906
transform 1 0 14000 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16352 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22624 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform -1 0 23296 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _120_
timestamp 1698175906
transform -1 0 14224 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform 1 0 17808 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _122_
timestamp 1698175906
transform -1 0 15456 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _123_
timestamp 1698175906
transform -1 0 14784 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform -1 0 21280 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _126_
timestamp 1698175906
transform -1 0 19936 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _127_
timestamp 1698175906
transform 1 0 19488 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _128_
timestamp 1698175906
transform 1 0 20720 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _130_
timestamp 1698175906
transform -1 0 20384 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _131_
timestamp 1698175906
transform 1 0 19936 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _132_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19264 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _133_
timestamp 1698175906
transform 1 0 21280 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _134_
timestamp 1698175906
transform -1 0 23856 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21392 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _136_
timestamp 1698175906
transform 1 0 17248 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1698175906
transform -1 0 14112 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform -1 0 11424 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _139_
timestamp 1698175906
transform -1 0 11648 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _140_
timestamp 1698175906
transform -1 0 20944 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _141_
timestamp 1698175906
transform 1 0 23296 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _142_
timestamp 1698175906
transform -1 0 24752 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _143_
timestamp 1698175906
transform -1 0 24080 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _144_
timestamp 1698175906
transform -1 0 19152 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _145_
timestamp 1698175906
transform -1 0 21952 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _146_
timestamp 1698175906
transform 1 0 19936 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _147_
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _148_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _149_
timestamp 1698175906
transform 1 0 15456 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _150_
timestamp 1698175906
transform 1 0 14560 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _151_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15008 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _152_
timestamp 1698175906
transform -1 0 17472 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _153_
timestamp 1698175906
transform -1 0 19264 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _154_
timestamp 1698175906
transform 1 0 15680 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _155_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16464 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _156_
timestamp 1698175906
transform 1 0 27440 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _157_
timestamp 1698175906
transform -1 0 27328 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _158_
timestamp 1698175906
transform 1 0 20160 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _159_
timestamp 1698175906
transform 1 0 19152 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform -1 0 27328 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _161_
timestamp 1698175906
transform -1 0 26432 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _162_
timestamp 1698175906
transform -1 0 18592 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _163_
timestamp 1698175906
transform 1 0 12320 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _164_
timestamp 1698175906
transform -1 0 11424 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _165_
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _166_
timestamp 1698175906
transform -1 0 13216 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _167_
timestamp 1698175906
transform 1 0 10752 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _168_
timestamp 1698175906
transform -1 0 22624 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _169_
timestamp 1698175906
transform 1 0 27440 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _170_
timestamp 1698175906
transform -1 0 27328 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _171_
timestamp 1698175906
transform 1 0 24304 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _172_
timestamp 1698175906
transform 1 0 18032 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _173_
timestamp 1698175906
transform 1 0 25424 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _174_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22624 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _175_
timestamp 1698175906
transform 1 0 23072 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _176_
timestamp 1698175906
transform 1 0 23968 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform 1 0 25200 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _178_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25312 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _179_
timestamp 1698175906
transform -1 0 26432 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _180_
timestamp 1698175906
transform -1 0 18928 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _181_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18816 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _182_
timestamp 1698175906
transform -1 0 17920 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _183_
timestamp 1698175906
transform 1 0 13328 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _184_
timestamp 1698175906
transform -1 0 12768 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _185_
timestamp 1698175906
transform 1 0 23184 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _186_
timestamp 1698175906
transform 1 0 21616 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _187_
timestamp 1698175906
transform 1 0 22176 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _188_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16016 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _189_
timestamp 1698175906
transform -1 0 21616 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _190_
timestamp 1698175906
transform 1 0 17360 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _191_
timestamp 1698175906
transform 1 0 12096 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _192_
timestamp 1698175906
transform 1 0 11648 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _193_
timestamp 1698175906
transform 1 0 21616 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_
timestamp 1698175906
transform -1 0 11984 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1698175906
transform 1 0 22176 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _196_
timestamp 1698175906
transform 1 0 19152 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _197_
timestamp 1698175906
transform -1 0 15232 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _198_
timestamp 1698175906
transform 1 0 13776 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _199_
timestamp 1698175906
transform 1 0 25536 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _200_
timestamp 1698175906
transform 1 0 18368 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1698175906
transform 1 0 25424 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_
timestamp 1698175906
transform -1 0 12432 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform -1 0 12656 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform 1 0 26432 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform 1 0 25312 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform 1 0 25424 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform 1 0 15456 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform -1 0 13104 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 21616 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _212_
timestamp 1698175906
transform -1 0 15904 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _213_
timestamp 1698175906
transform 1 0 26992 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _214_
timestamp 1698175906
transform 1 0 27776 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _215_
timestamp 1698175906
transform 1 0 27776 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _216_
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _217_
timestamp 1698175906
transform 1 0 28896 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21840 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__CLK
timestamp 1698175906
transform 1 0 24864 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1698175906
transform 1 0 25424 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__CLK
timestamp 1698175906
transform -1 0 22848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__CLK
timestamp 1698175906
transform 1 0 28784 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__CLK
timestamp 1698175906
transform 1 0 21840 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__CLK
timestamp 1698175906
transform 1 0 29232 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform 1 0 26208 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 29232 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 28560 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 28896 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 19376 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 20944 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 22176 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_165 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698175906
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698175906
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_139
timestamp 1698175906
transform 1 0 16912 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698175906
transform 1 0 20608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_88 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11200 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_96
timestamp 1698175906
transform 1 0 12096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_100
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_131
timestamp 1698175906
transform 1 0 16016 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698175906
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_150
timestamp 1698175906
transform 1 0 18144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_181
timestamp 1698175906
transform 1 0 21616 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_185
timestamp 1698175906
transform 1 0 22064 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_201
timestamp 1698175906
transform 1 0 23856 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_144
timestamp 1698175906
transform 1 0 17472 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_152
timestamp 1698175906
transform 1 0 18368 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698175906
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_181
timestamp 1698175906
transform 1 0 21616 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 4480 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_80
timestamp 1698175906
transform 1 0 10304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_84
timestamp 1698175906
transform 1 0 10752 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_90
timestamp 1698175906
transform 1 0 11424 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_106
timestamp 1698175906
transform 1 0 13216 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_114
timestamp 1698175906
transform 1 0 14112 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_118
timestamp 1698175906
transform 1 0 14560 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_125
timestamp 1698175906
transform 1 0 15344 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_133
timestamp 1698175906
transform 1 0 16240 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698175906
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_176
timestamp 1698175906
transform 1 0 21056 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_180
timestamp 1698175906
transform 1 0 21504 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_216
timestamp 1698175906
transform 1 0 25536 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_69
timestamp 1698175906
transform 1 0 9072 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_99
timestamp 1698175906
transform 1 0 12432 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_103
timestamp 1698175906
transform 1 0 12880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_135
timestamp 1698175906
transform 1 0 16464 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_151
timestamp 1698175906
transform 1 0 18256 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_153
timestamp 1698175906
transform 1 0 18480 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_159
timestamp 1698175906
transform 1 0 19152 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698175906
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_185
timestamp 1698175906
transform 1 0 22064 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_195
timestamp 1698175906
transform 1 0 23184 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_211
timestamp 1698175906
transform 1 0 24976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_213
timestamp 1698175906
transform 1 0 25200 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698175906
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_251
timestamp 1698175906
transform 1 0 29456 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_80
timestamp 1698175906
transform 1 0 10304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_84
timestamp 1698175906
transform 1 0 10752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_90
timestamp 1698175906
transform 1 0 11424 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_107
timestamp 1698175906
transform 1 0 13328 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_123
timestamp 1698175906
transform 1 0 15120 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_127
timestamp 1698175906
transform 1 0 15568 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698175906
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_150
timestamp 1698175906
transform 1 0 18144 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_154
timestamp 1698175906
transform 1 0 18592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_156
timestamp 1698175906
transform 1 0 18816 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_162
timestamp 1698175906
transform 1 0 19488 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_164
timestamp 1698175906
transform 1 0 19712 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_186
timestamp 1698175906
transform 1 0 22176 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_194
timestamp 1698175906
transform 1 0 23072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_241
timestamp 1698175906
transform 1 0 28336 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_245
timestamp 1698175906
transform 1 0 28784 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698175906
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_53
timestamp 1698175906
transform 1 0 7280 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_61
timestamp 1698175906
transform 1 0 8176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_65
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_95
timestamp 1698175906
transform 1 0 11984 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_103
timestamp 1698175906
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_120
timestamp 1698175906
transform 1 0 14784 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_124
timestamp 1698175906
transform 1 0 15232 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_160
timestamp 1698175906
transform 1 0 19264 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_190
timestamp 1698175906
transform 1 0 22624 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_203
timestamp 1698175906
transform 1 0 24080 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_214
timestamp 1698175906
transform 1 0 25312 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_223
timestamp 1698175906
transform 1 0 26320 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_227
timestamp 1698175906
transform 1 0 26768 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_235
timestamp 1698175906
transform 1 0 27664 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698175906
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 4480 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 8064 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_80
timestamp 1698175906
transform 1 0 10304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_138
timestamp 1698175906
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_184
timestamp 1698175906
transform 1 0 21952 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_200
timestamp 1698175906
transform 1 0 23744 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_208
timestamp 1698175906
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_220
timestamp 1698175906
transform 1 0 25984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_253
timestamp 1698175906
transform 1 0 29680 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_269
timestamp 1698175906
transform 1 0 31472 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698175906
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_69
timestamp 1698175906
transform 1 0 9072 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_77
timestamp 1698175906
transform 1 0 9968 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_81
timestamp 1698175906
transform 1 0 10416 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_83
timestamp 1698175906
transform 1 0 10640 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_92
timestamp 1698175906
transform 1 0 11648 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_100
timestamp 1698175906
transform 1 0 12544 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698175906
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_118
timestamp 1698175906
transform 1 0 14560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_122
timestamp 1698175906
transform 1 0 15008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_124
timestamp 1698175906
transform 1 0 15232 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_200
timestamp 1698175906
transform 1 0 23744 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_208
timestamp 1698175906
transform 1 0 24640 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_212
timestamp 1698175906
transform 1 0 25088 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_224
timestamp 1698175906
transform 1 0 26432 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_240
timestamp 1698175906
transform 1 0 28224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_106
timestamp 1698175906
transform 1 0 13216 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_122
timestamp 1698175906
transform 1 0 15008 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_126
timestamp 1698175906
transform 1 0 15456 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_134
timestamp 1698175906
transform 1 0 16352 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_214
timestamp 1698175906
transform 1 0 25312 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_244
timestamp 1698175906
transform 1 0 28672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_248
timestamp 1698175906
transform 1 0 29120 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 4480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_109
timestamp 1698175906
transform 1 0 13552 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_115
timestamp 1698175906
transform 1 0 14224 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_123
timestamp 1698175906
transform 1 0 15120 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_127
timestamp 1698175906
transform 1 0 15568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_139
timestamp 1698175906
transform 1 0 16912 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_141
timestamp 1698175906
transform 1 0 17136 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_148
timestamp 1698175906
transform 1 0 17920 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_159
timestamp 1698175906
transform 1 0 19152 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_163
timestamp 1698175906
transform 1 0 19600 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_170
timestamp 1698175906
transform 1 0 20384 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_184
timestamp 1698175906
transform 1 0 21952 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_236
timestamp 1698175906
transform 1 0 27776 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_88
timestamp 1698175906
transform 1 0 11200 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_125
timestamp 1698175906
transform 1 0 15344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_127
timestamp 1698175906
transform 1 0 15568 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_156
timestamp 1698175906
transform 1 0 18816 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_160
timestamp 1698175906
transform 1 0 19264 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_167
timestamp 1698175906
transform 1 0 20048 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_171
timestamp 1698175906
transform 1 0 20496 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_225
timestamp 1698175906
transform 1 0 26544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_232
timestamp 1698175906
transform 1 0 27328 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_242
timestamp 1698175906
transform 1 0 28448 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_252
timestamp 1698175906
transform 1 0 29568 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_268
timestamp 1698175906
transform 1 0 31360 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698175906
transform 1 0 32256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_114
timestamp 1698175906
transform 1 0 14112 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_122
timestamp 1698175906
transform 1 0 15008 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_134
timestamp 1698175906
transform 1 0 16352 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_142
timestamp 1698175906
transform 1 0 17248 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_146
timestamp 1698175906
transform 1 0 17696 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_157
timestamp 1698175906
transform 1 0 18928 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_173
timestamp 1698175906
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_189
timestamp 1698175906
transform 1 0 22512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_201
timestamp 1698175906
transform 1 0 23856 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_209
timestamp 1698175906
transform 1 0 24752 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_212
timestamp 1698175906
transform 1 0 25088 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_228
timestamp 1698175906
transform 1 0 26880 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_232
timestamp 1698175906
transform 1 0 27328 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_238
timestamp 1698175906
transform 1 0 28000 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698175906
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_88
timestamp 1698175906
transform 1 0 11200 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_96
timestamp 1698175906
transform 1 0 12096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_102
timestamp 1698175906
transform 1 0 12768 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_106
timestamp 1698175906
transform 1 0 13216 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_116
timestamp 1698175906
transform 1 0 14336 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_120
timestamp 1698175906
transform 1 0 14784 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_133
timestamp 1698175906
transform 1 0 16240 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_137
timestamp 1698175906
transform 1 0 16688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_158
timestamp 1698175906
transform 1 0 19040 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_166
timestamp 1698175906
transform 1 0 19936 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_176
timestamp 1698175906
transform 1 0 21056 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_192
timestamp 1698175906
transform 1 0 22848 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_202
timestamp 1698175906
transform 1 0 23968 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_216
timestamp 1698175906
transform 1 0 25536 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_218
timestamp 1698175906
transform 1 0 25760 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_224
timestamp 1698175906
transform 1 0 26432 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_226
timestamp 1698175906
transform 1 0 26656 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_232
timestamp 1698175906
transform 1 0 27328 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_238
timestamp 1698175906
transform 1 0 28000 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_242
timestamp 1698175906
transform 1 0 28448 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_244
timestamp 1698175906
transform 1 0 28672 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_247
timestamp 1698175906
transform 1 0 29008 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 36512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 37408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_69
timestamp 1698175906
transform 1 0 9072 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_73
timestamp 1698175906
transform 1 0 9520 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_75
timestamp 1698175906
transform 1 0 9744 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_115
timestamp 1698175906
transform 1 0 14224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_117
timestamp 1698175906
transform 1 0 14448 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_123
timestamp 1698175906
transform 1 0 15120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_125
timestamp 1698175906
transform 1 0 15344 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_155
timestamp 1698175906
transform 1 0 18704 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_185
timestamp 1698175906
transform 1 0 22064 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_193
timestamp 1698175906
transform 1 0 22960 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_197
timestamp 1698175906
transform 1 0 23408 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_199
timestamp 1698175906
transform 1 0 23632 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_209
timestamp 1698175906
transform 1 0 24752 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_213
timestamp 1698175906
transform 1 0 25200 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_215
timestamp 1698175906
transform 1 0 25424 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_253
timestamp 1698175906
transform 1 0 29680 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_285
timestamp 1698175906
transform 1 0 33264 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_301
timestamp 1698175906
transform 1 0 35056 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_309
timestamp 1698175906
transform 1 0 35952 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_313
timestamp 1698175906
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 4480 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_88
timestamp 1698175906
transform 1 0 11200 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_92
timestamp 1698175906
transform 1 0 11648 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_94
timestamp 1698175906
transform 1 0 11872 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_130
timestamp 1698175906
transform 1 0 15904 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698175906
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_148
timestamp 1698175906
transform 1 0 17920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_181
timestamp 1698175906
transform 1 0 21616 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_185
timestamp 1698175906
transform 1 0 22064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_193
timestamp 1698175906
transform 1 0 22960 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_197
timestamp 1698175906
transform 1 0 23408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_203
timestamp 1698175906
transform 1 0 24080 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698175906
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_214
timestamp 1698175906
transform 1 0 25312 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_217
timestamp 1698175906
transform 1 0 25648 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_225
timestamp 1698175906
transform 1 0 26544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_232
timestamp 1698175906
transform 1 0 27328 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_242
timestamp 1698175906
transform 1 0 28448 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_274
timestamp 1698175906
transform 1 0 32032 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698175906
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 36512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 37408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698175906
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_185
timestamp 1698175906
transform 1 0 22064 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_251
timestamp 1698175906
transform 1 0 29456 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_158
timestamp 1698175906
transform 1 0 19040 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_188
timestamp 1698175906
transform 1 0 22400 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_192
timestamp 1698175906
transform 1 0 22848 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698175906
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_314
timestamp 1698175906
transform 1 0 36512 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_322
timestamp 1698175906
transform 1 0 37408 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_174
timestamp 1698175906
transform 1 0 20832 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_201
timestamp 1698175906
transform 1 0 23856 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_314
timestamp 1698175906
transform 1 0 36512 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_330
timestamp 1698175906
transform 1 0 38304 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_338
timestamp 1698175906
transform 1 0 39200 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_342
timestamp 1698175906
transform 1 0 39648 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_344
timestamp 1698175906
transform 1 0 39872 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_206
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_210
timestamp 1698175906
transform 1 0 24864 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_237
timestamp 1698175906
transform 1 0 27888 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita54_26 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 39984 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16912 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 37520 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 37520 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 4480 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 20944 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 37520 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 37520 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 21280 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform -1 0 4480 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 4480 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 24976 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 37520 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 37520 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 4480 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 4480 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 41200 36960 42000 37072 0 FreeSans 448 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 41200 21504 42000 21616 0 FreeSans 448 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 18816 41200 18928 42000 0 FreeSans 448 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 41200 26880 42000 26992 0 FreeSans 448 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 41200 24864 42000 24976 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 20832 41200 20944 42000 0 FreeSans 448 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 41200 24192 42000 24304 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 41200 18816 42000 18928 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 24864 41200 24976 42000 0 FreeSans 448 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 41200 26208 42000 26320 0 FreeSans 448 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 41200 25536 42000 25648 0 FreeSans 448 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 41200 17472 42000 17584 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 26264 24472 26264 24472 0 _000_
rlabel metal2 11144 17304 11144 17304 0 _001_
rlabel metal2 11032 21224 11032 21224 0 _002_
rlabel metal2 27048 21532 27048 21532 0 _003_
rlabel metal2 26264 18144 26264 18144 0 _004_
rlabel metal3 25144 18312 25144 18312 0 _005_
rlabel metal2 26152 21168 26152 21168 0 _006_
rlabel metal2 16408 25984 16408 25984 0 _007_
rlabel metal2 12488 25144 12488 25144 0 _008_
rlabel metal2 22624 16968 22624 16968 0 _009_
rlabel metal2 15064 16072 15064 16072 0 _010_
rlabel metal2 21896 17864 21896 17864 0 _011_
rlabel metal2 18816 15960 18816 15960 0 _012_
rlabel metal2 13720 22456 13720 22456 0 _013_
rlabel metal2 13608 19600 13608 19600 0 _014_
rlabel metal2 22568 23464 22568 23464 0 _015_
rlabel metal2 11200 19320 11200 19320 0 _016_
rlabel metal3 23464 26488 23464 26488 0 _017_
rlabel metal2 20104 27300 20104 27300 0 _018_
rlabel metal2 14280 25480 14280 25480 0 _019_
rlabel metal3 15008 16184 15008 16184 0 _020_
rlabel metal2 26824 25144 26824 25144 0 _021_
rlabel metal2 19376 25592 19376 25592 0 _022_
rlabel metal2 21336 25592 21336 25592 0 _023_
rlabel metal2 16352 23688 16352 23688 0 _024_
rlabel metal2 15064 25032 15064 25032 0 _025_
rlabel metal3 16520 15960 16520 15960 0 _026_
rlabel metal2 18760 18760 18760 18760 0 _027_
rlabel metal2 15960 17976 15960 17976 0 _028_
rlabel metal2 27160 24584 27160 24584 0 _029_
rlabel metal3 19880 24920 19880 24920 0 _030_
rlabel metal2 26264 25424 26264 25424 0 _031_
rlabel metal2 18312 18872 18312 18872 0 _032_
rlabel metal3 12040 16968 12040 16968 0 _033_
rlabel metal2 17528 21056 17528 21056 0 _034_
rlabel metal2 11592 21056 11592 21056 0 _035_
rlabel metal2 25816 19880 25816 19880 0 _036_
rlabel metal2 27160 23688 27160 23688 0 _037_
rlabel metal2 25480 19264 25480 19264 0 _038_
rlabel metal2 18368 22120 18368 22120 0 _039_
rlabel metal2 24360 19488 24360 19488 0 _040_
rlabel metal2 24024 18872 24024 18872 0 _041_
rlabel metal2 25816 20776 25816 20776 0 _042_
rlabel metal2 26376 21000 26376 21000 0 _043_
rlabel metal2 18480 23128 18480 23128 0 _044_
rlabel metal2 17808 26264 17808 26264 0 _045_
rlabel metal3 13216 24584 13216 24584 0 _046_
rlabel metal2 22568 17920 22568 17920 0 _047_
rlabel metal2 22344 18032 22344 18032 0 _048_
rlabel metal2 16632 20888 16632 20888 0 _049_
rlabel metal2 16016 19096 16016 19096 0 _050_
rlabel metal2 19208 17696 19208 17696 0 _051_
rlabel metal2 21112 18760 21112 18760 0 _052_
rlabel metal2 21448 18704 21448 18704 0 _053_
rlabel metal2 15624 18872 15624 18872 0 _054_
rlabel metal2 17976 20776 17976 20776 0 _055_
rlabel metal3 18536 20104 18536 20104 0 _056_
rlabel metal2 15792 17864 15792 17864 0 _057_
rlabel metal2 19376 19208 19376 19208 0 _058_
rlabel metal3 23800 20664 23800 20664 0 _059_
rlabel metal2 15960 21728 15960 21728 0 _060_
rlabel metal2 16744 22848 16744 22848 0 _061_
rlabel metal2 19656 22960 19656 22960 0 _062_
rlabel metal2 15792 22904 15792 22904 0 _063_
rlabel metal2 19656 19824 19656 19824 0 _064_
rlabel metal2 14784 16968 14784 16968 0 _065_
rlabel metal2 19264 15960 19264 15960 0 _066_
rlabel metal2 11480 20384 11480 20384 0 _067_
rlabel metal2 14280 21560 14280 21560 0 _068_
rlabel metal2 21112 19600 21112 19600 0 _069_
rlabel metal2 22792 20048 22792 20048 0 _070_
rlabel metal2 19656 24640 19656 24640 0 _071_
rlabel metal2 17976 19488 17976 19488 0 _072_
rlabel metal2 13720 19600 13720 19600 0 _073_
rlabel metal2 14168 19208 14168 19208 0 _074_
rlabel metal3 22848 25368 22848 25368 0 _075_
rlabel metal2 19376 20104 19376 20104 0 _076_
rlabel metal2 20888 24024 20888 24024 0 _077_
rlabel metal2 21000 23576 21000 23576 0 _078_
rlabel metal2 20216 20832 20216 20832 0 _079_
rlabel metal2 19768 25536 19768 25536 0 _080_
rlabel metal3 20216 20216 20216 20216 0 _081_
rlabel metal2 21560 21840 21560 21840 0 _082_
rlabel metal2 25704 24024 25704 24024 0 _083_
rlabel metal2 22120 23800 22120 23800 0 _084_
rlabel metal2 17752 23632 17752 23632 0 _085_
rlabel metal3 11984 18536 11984 18536 0 _086_
rlabel metal2 10920 19320 10920 19320 0 _087_
rlabel metal2 20664 18760 20664 18760 0 _088_
rlabel metal2 27720 24696 27720 24696 0 _089_
rlabel metal2 23968 25592 23968 25592 0 _090_
rlabel metal3 17528 17640 17528 17640 0 _091_
rlabel metal2 20552 25312 20552 25312 0 _092_
rlabel metal2 20440 20048 20440 20048 0 _093_
rlabel metal2 19432 21840 19432 21840 0 clk
rlabel metal2 22344 22008 22344 22008 0 clknet_0_clk
rlabel metal2 17528 14812 17528 14812 0 clknet_1_0__leaf_clk
rlabel metal2 22792 27384 22792 27384 0 clknet_1_1__leaf_clk
rlabel metal2 19880 16016 19880 16016 0 dut54.count\[0\]
rlabel metal2 20384 14616 20384 14616 0 dut54.count\[1\]
rlabel metal2 16632 22736 16632 22736 0 dut54.count\[2\]
rlabel metal2 16744 20384 16744 20384 0 dut54.count\[3\]
rlabel metal2 17080 5964 17080 5964 0 net1
rlabel metal2 29176 23912 29176 23912 0 net10
rlabel metal2 28392 18480 28392 18480 0 net11
rlabel metal2 37688 18704 37688 18704 0 net12
rlabel metal2 28168 18704 28168 18704 0 net13
rlabel metal2 22176 27720 22176 27720 0 net14
rlabel metal2 9352 17696 9352 17696 0 net15
rlabel metal3 6888 21448 6888 21448 0 net16
rlabel metal2 25200 27048 25200 27048 0 net17
rlabel metal3 31920 22960 31920 22960 0 net18
rlabel metal3 30100 26376 30100 26376 0 net19
rlabel metal3 28280 23184 28280 23184 0 net2
rlabel metal2 37912 25760 37912 25760 0 net20
rlabel metal2 10024 25536 10024 25536 0 net21
rlabel metal2 12936 16016 12936 16016 0 net22
rlabel metal2 8904 19656 8904 19656 0 net23
rlabel metal3 37688 23184 37688 23184 0 net24
rlabel metal2 24696 17192 24696 17192 0 net25
rlabel metal2 40264 37184 40264 37184 0 net26
rlabel metal2 28504 21392 28504 21392 0 net3
rlabel metal2 18536 25648 18536 25648 0 net4
rlabel metal3 9856 27048 9856 27048 0 net5
rlabel metal2 28504 27496 28504 27496 0 net6
rlabel metal2 29288 25536 29288 25536 0 net7
rlabel metal2 12152 26208 12152 26208 0 net8
rlabel metal2 21448 26040 21448 26040 0 net9
rlabel metal2 16856 2086 16856 2086 0 segm[10]
rlabel metal2 40040 22344 40040 22344 0 segm[11]
rlabel metal2 40040 21504 40040 21504 0 segm[12]
rlabel metal2 18872 39690 18872 39690 0 segm[13]
rlabel metal3 1358 26264 1358 26264 0 segm[1]
rlabel metal2 39928 27328 39928 27328 0 segm[2]
rlabel metal2 40040 25256 40040 25256 0 segm[3]
rlabel metal3 1358 25592 1358 25592 0 segm[4]
rlabel metal2 20888 39354 20888 39354 0 segm[5]
rlabel metal2 40040 24360 40040 24360 0 segm[6]
rlabel metal2 40040 19096 40040 19096 0 segm[7]
rlabel metal3 40642 18200 40642 18200 0 segm[8]
rlabel metal2 40040 19656 40040 19656 0 segm[9]
rlabel metal2 22232 39746 22232 39746 0 sel[0]
rlabel metal3 1358 17528 1358 17528 0 sel[10]
rlabel metal3 1358 21560 1358 21560 0 sel[11]
rlabel metal2 24920 39746 24920 39746 0 sel[1]
rlabel metal2 40040 23800 40040 23800 0 sel[2]
rlabel metal2 40040 26712 40040 26712 0 sel[3]
rlabel metal2 39928 25872 39928 25872 0 sel[4]
rlabel metal3 1414 24920 1414 24920 0 sel[5]
rlabel metal3 1358 16856 1358 16856 0 sel[6]
rlabel metal3 1358 19544 1358 19544 0 sel[7]
rlabel metal3 40642 22904 40642 22904 0 sel[8]
rlabel metal2 40040 17640 40040 17640 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
