magic
tech gf180mcuD
magscale 1 10
timestamp 1699642721
<< metal1 >>
rect 26898 38558 26910 38610
rect 26962 38607 26974 38610
rect 28354 38607 28366 38610
rect 26962 38561 28366 38607
rect 26962 38558 26974 38561
rect 28354 38558 28366 38561
rect 28418 38558 28430 38610
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 22430 38274 22482 38286
rect 19506 38222 19518 38274
rect 19570 38222 19582 38274
rect 22430 38210 22482 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 17826 37998 17838 38050
rect 17890 37998 17902 38050
rect 21746 37998 21758 38050
rect 21810 37998 21822 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 27470 37938 27522 37950
rect 27470 37874 27522 37886
rect 28366 37938 28418 37950
rect 28366 37874 28418 37886
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 19070 37490 19122 37502
rect 19070 37426 19122 37438
rect 21422 37490 21474 37502
rect 21422 37426 21474 37438
rect 26798 37490 26850 37502
rect 26798 37426 26850 37438
rect 19618 37214 19630 37266
rect 19682 37214 19694 37266
rect 20626 37214 20638 37266
rect 20690 37214 20702 37266
rect 25778 37214 25790 37266
rect 25842 37214 25854 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 17390 36706 17442 36718
rect 17390 36642 17442 36654
rect 16594 36430 16606 36482
rect 16658 36430 16670 36482
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 22318 29426 22370 29438
rect 18946 29374 18958 29426
rect 19010 29374 19022 29426
rect 22318 29362 22370 29374
rect 19618 29262 19630 29314
rect 19682 29262 19694 29314
rect 21746 29262 21758 29314
rect 21810 29262 21822 29314
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 19170 28702 19182 28754
rect 19234 28702 19246 28754
rect 16370 28590 16382 28642
rect 16434 28590 16446 28642
rect 19630 28530 19682 28542
rect 17042 28478 17054 28530
rect 17106 28478 17118 28530
rect 19630 28466 19682 28478
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 17390 28082 17442 28094
rect 17390 28018 17442 28030
rect 19070 28082 19122 28094
rect 19070 28018 19122 28030
rect 19854 28082 19906 28094
rect 19854 28018 19906 28030
rect 20750 28082 20802 28094
rect 20750 28018 20802 28030
rect 17614 27970 17666 27982
rect 17614 27906 17666 27918
rect 20078 27970 20130 27982
rect 20078 27906 20130 27918
rect 17726 27858 17778 27870
rect 14802 27806 14814 27858
rect 14866 27806 14878 27858
rect 17726 27794 17778 27806
rect 18846 27858 18898 27870
rect 18846 27794 18898 27806
rect 19182 27858 19234 27870
rect 19182 27794 19234 27806
rect 20190 27858 20242 27870
rect 20190 27794 20242 27806
rect 20526 27858 20578 27870
rect 20526 27794 20578 27806
rect 20862 27858 20914 27870
rect 21746 27806 21758 27858
rect 21810 27806 21822 27858
rect 20862 27794 20914 27806
rect 15374 27746 15426 27758
rect 25342 27746 25394 27758
rect 12002 27694 12014 27746
rect 12066 27694 12078 27746
rect 14130 27694 14142 27746
rect 14194 27694 14206 27746
rect 22418 27694 22430 27746
rect 22482 27694 22494 27746
rect 24546 27694 24558 27746
rect 24610 27694 24622 27746
rect 15374 27682 15426 27694
rect 25342 27682 25394 27694
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 22542 27298 22594 27310
rect 22542 27234 22594 27246
rect 22430 27074 22482 27086
rect 22430 27010 22482 27022
rect 23326 27074 23378 27086
rect 23326 27010 23378 27022
rect 18846 26962 18898 26974
rect 18846 26898 18898 26910
rect 18958 26962 19010 26974
rect 18958 26898 19010 26910
rect 22542 26962 22594 26974
rect 22542 26898 22594 26910
rect 22990 26962 23042 26974
rect 22990 26898 23042 26910
rect 23214 26962 23266 26974
rect 23214 26898 23266 26910
rect 19182 26850 19234 26862
rect 19182 26786 19234 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 25342 26402 25394 26414
rect 25342 26338 25394 26350
rect 4274 26238 4286 26290
rect 4338 26238 4350 26290
rect 13570 26238 13582 26290
rect 13634 26238 13646 26290
rect 20290 26238 20302 26290
rect 20354 26238 20366 26290
rect 16830 26178 16882 26190
rect 20750 26178 20802 26190
rect 14242 26126 14254 26178
rect 14306 26126 14318 26178
rect 16370 26126 16382 26178
rect 16434 26126 16446 26178
rect 17378 26126 17390 26178
rect 17442 26126 17454 26178
rect 19506 26126 19518 26178
rect 19570 26126 19582 26178
rect 16830 26114 16882 26126
rect 20750 26114 20802 26126
rect 1934 26066 1986 26078
rect 1934 26002 1986 26014
rect 25230 26066 25282 26078
rect 25230 26002 25282 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 15822 25730 15874 25742
rect 15822 25666 15874 25678
rect 21646 25730 21698 25742
rect 21646 25666 21698 25678
rect 14478 25618 14530 25630
rect 40014 25618 40066 25630
rect 19506 25566 19518 25618
rect 19570 25566 19582 25618
rect 25666 25566 25678 25618
rect 25730 25566 25742 25618
rect 14478 25554 14530 25566
rect 40014 25554 40066 25566
rect 15150 25506 15202 25518
rect 14914 25454 14926 25506
rect 14978 25454 14990 25506
rect 15150 25442 15202 25454
rect 19182 25506 19234 25518
rect 22866 25454 22878 25506
rect 22930 25454 22942 25506
rect 37650 25454 37662 25506
rect 37714 25454 37726 25506
rect 19182 25442 19234 25454
rect 14366 25394 14418 25406
rect 14366 25330 14418 25342
rect 15374 25394 15426 25406
rect 15374 25330 15426 25342
rect 15486 25394 15538 25406
rect 15486 25330 15538 25342
rect 15934 25394 15986 25406
rect 15934 25330 15986 25342
rect 19742 25394 19794 25406
rect 19742 25330 19794 25342
rect 21534 25394 21586 25406
rect 21534 25330 21586 25342
rect 22094 25394 22146 25406
rect 26126 25394 26178 25406
rect 22418 25342 22430 25394
rect 22482 25342 22494 25394
rect 23538 25342 23550 25394
rect 23602 25342 23614 25394
rect 22094 25330 22146 25342
rect 26126 25330 26178 25342
rect 26238 25394 26290 25406
rect 26238 25330 26290 25342
rect 14590 25282 14642 25294
rect 14590 25218 14642 25230
rect 19518 25282 19570 25294
rect 19518 25218 19570 25230
rect 21646 25282 21698 25294
rect 21646 25218 21698 25230
rect 26462 25282 26514 25294
rect 26462 25218 26514 25230
rect 26798 25282 26850 25294
rect 26798 25218 26850 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 16046 24946 16098 24958
rect 16046 24882 16098 24894
rect 16158 24946 16210 24958
rect 20190 24946 20242 24958
rect 17714 24894 17726 24946
rect 17778 24894 17790 24946
rect 16158 24882 16210 24894
rect 20190 24882 20242 24894
rect 21758 24946 21810 24958
rect 21758 24882 21810 24894
rect 23326 24946 23378 24958
rect 23326 24882 23378 24894
rect 28590 24946 28642 24958
rect 28590 24882 28642 24894
rect 20526 24834 20578 24846
rect 20526 24770 20578 24782
rect 21534 24834 21586 24846
rect 21534 24770 21586 24782
rect 23438 24834 23490 24846
rect 23438 24770 23490 24782
rect 13918 24722 13970 24734
rect 4274 24670 4286 24722
rect 4338 24670 4350 24722
rect 13458 24670 13470 24722
rect 13522 24670 13534 24722
rect 13918 24658 13970 24670
rect 16382 24722 16434 24734
rect 17390 24722 17442 24734
rect 16594 24670 16606 24722
rect 16658 24670 16670 24722
rect 16382 24658 16434 24670
rect 17390 24658 17442 24670
rect 20078 24722 20130 24734
rect 20078 24658 20130 24670
rect 20302 24722 20354 24734
rect 22430 24722 22482 24734
rect 21186 24670 21198 24722
rect 21250 24670 21262 24722
rect 22754 24670 22766 24722
rect 22818 24670 22830 24722
rect 25330 24670 25342 24722
rect 25394 24670 25406 24722
rect 20302 24658 20354 24670
rect 22430 24658 22482 24670
rect 21646 24610 21698 24622
rect 10546 24558 10558 24610
rect 10610 24558 10622 24610
rect 12674 24558 12686 24610
rect 12738 24558 12750 24610
rect 16034 24558 16046 24610
rect 16098 24558 16110 24610
rect 21646 24546 21698 24558
rect 22990 24610 23042 24622
rect 22990 24546 23042 24558
rect 23214 24610 23266 24622
rect 26002 24558 26014 24610
rect 26066 24558 26078 24610
rect 28130 24558 28142 24610
rect 28194 24558 28206 24610
rect 23214 24546 23266 24558
rect 1934 24498 1986 24510
rect 1934 24434 1986 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 12462 24162 12514 24174
rect 12462 24098 12514 24110
rect 25566 24050 25618 24062
rect 13794 23998 13806 24050
rect 13858 23998 13870 24050
rect 20178 23998 20190 24050
rect 20242 23998 20254 24050
rect 25566 23986 25618 23998
rect 12350 23938 12402 23950
rect 13918 23938 13970 23950
rect 25678 23938 25730 23950
rect 13682 23886 13694 23938
rect 13746 23886 13758 23938
rect 17266 23886 17278 23938
rect 17330 23886 17342 23938
rect 12350 23874 12402 23886
rect 13918 23874 13970 23886
rect 25678 23874 25730 23886
rect 26126 23938 26178 23950
rect 26126 23874 26178 23886
rect 14366 23826 14418 23838
rect 18050 23774 18062 23826
rect 18114 23774 18126 23826
rect 14366 23762 14418 23774
rect 14142 23714 14194 23726
rect 14142 23650 14194 23662
rect 16942 23714 16994 23726
rect 16942 23650 16994 23662
rect 25454 23714 25506 23726
rect 25454 23650 25506 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 19406 23378 19458 23390
rect 19406 23314 19458 23326
rect 19518 23378 19570 23390
rect 19518 23314 19570 23326
rect 19630 23378 19682 23390
rect 19630 23314 19682 23326
rect 19966 23378 20018 23390
rect 19966 23314 20018 23326
rect 13694 23266 13746 23278
rect 13694 23202 13746 23214
rect 18174 23266 18226 23278
rect 18174 23202 18226 23214
rect 20190 23266 20242 23278
rect 20190 23202 20242 23214
rect 26574 23266 26626 23278
rect 26574 23202 26626 23214
rect 26686 23266 26738 23278
rect 26786 23214 26798 23266
rect 26850 23214 26862 23266
rect 26686 23202 26738 23214
rect 13358 23154 13410 23166
rect 13358 23090 13410 23102
rect 16270 23154 16322 23166
rect 16270 23090 16322 23102
rect 16494 23154 16546 23166
rect 18510 23154 18562 23166
rect 19294 23154 19346 23166
rect 16818 23102 16830 23154
rect 16882 23102 16894 23154
rect 19058 23102 19070 23154
rect 19122 23102 19134 23154
rect 16494 23090 16546 23102
rect 18510 23090 18562 23102
rect 19294 23090 19346 23102
rect 20302 23154 20354 23166
rect 20302 23090 20354 23102
rect 20862 23154 20914 23166
rect 20862 23090 20914 23102
rect 21198 23154 21250 23166
rect 21198 23090 21250 23102
rect 21310 23154 21362 23166
rect 26350 23154 26402 23166
rect 24658 23102 24670 23154
rect 24722 23102 24734 23154
rect 21310 23090 21362 23102
rect 26350 23090 26402 23102
rect 16382 23042 16434 23054
rect 16382 22978 16434 22990
rect 20974 23042 21026 23054
rect 25342 23042 25394 23054
rect 21746 22990 21758 23042
rect 21810 22990 21822 23042
rect 23874 22990 23886 23042
rect 23938 22990 23950 23042
rect 26674 22990 26686 23042
rect 26738 22990 26750 23042
rect 20974 22978 21026 22990
rect 25342 22978 25394 22990
rect 18286 22930 18338 22942
rect 18286 22866 18338 22878
rect 18622 22930 18674 22942
rect 18622 22866 18674 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 17502 22594 17554 22606
rect 17502 22530 17554 22542
rect 19182 22594 19234 22606
rect 19182 22530 19234 22542
rect 19294 22594 19346 22606
rect 19294 22530 19346 22542
rect 28142 22594 28194 22606
rect 28142 22530 28194 22542
rect 40014 22482 40066 22494
rect 10658 22430 10670 22482
rect 10722 22430 10734 22482
rect 12786 22430 12798 22482
rect 12850 22430 12862 22482
rect 40014 22418 40066 22430
rect 14030 22370 14082 22382
rect 9986 22318 9998 22370
rect 10050 22318 10062 22370
rect 14030 22306 14082 22318
rect 17614 22370 17666 22382
rect 18958 22370 19010 22382
rect 18722 22318 18734 22370
rect 18786 22318 18798 22370
rect 19618 22318 19630 22370
rect 19682 22318 19694 22370
rect 21858 22318 21870 22370
rect 21922 22318 21934 22370
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 17614 22306 17666 22318
rect 18958 22306 19010 22318
rect 15262 22258 15314 22270
rect 14354 22206 14366 22258
rect 14418 22206 14430 22258
rect 15262 22194 15314 22206
rect 18174 22258 18226 22270
rect 28254 22258 28306 22270
rect 19730 22206 19742 22258
rect 19794 22206 19806 22258
rect 20402 22206 20414 22258
rect 20466 22206 20478 22258
rect 26226 22206 26238 22258
rect 26290 22206 26302 22258
rect 18174 22194 18226 22206
rect 28254 22194 28306 22206
rect 13582 22146 13634 22158
rect 13582 22082 13634 22094
rect 15598 22146 15650 22158
rect 15598 22082 15650 22094
rect 17054 22146 17106 22158
rect 17054 22082 17106 22094
rect 17502 22146 17554 22158
rect 17502 22082 17554 22094
rect 18286 22146 18338 22158
rect 18286 22082 18338 22094
rect 18510 22146 18562 22158
rect 20626 22094 20638 22146
rect 20690 22094 20702 22146
rect 18510 22082 18562 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 12910 21810 12962 21822
rect 12910 21746 12962 21758
rect 15262 21810 15314 21822
rect 15262 21746 15314 21758
rect 15822 21810 15874 21822
rect 15822 21746 15874 21758
rect 16606 21810 16658 21822
rect 16606 21746 16658 21758
rect 14814 21698 14866 21710
rect 14814 21634 14866 21646
rect 15710 21698 15762 21710
rect 15710 21634 15762 21646
rect 15934 21698 15986 21710
rect 15934 21634 15986 21646
rect 16494 21698 16546 21710
rect 23886 21698 23938 21710
rect 17714 21646 17726 21698
rect 17778 21646 17790 21698
rect 21746 21646 21758 21698
rect 21810 21646 21822 21698
rect 27010 21646 27022 21698
rect 27074 21646 27086 21698
rect 16494 21634 16546 21646
rect 23886 21634 23938 21646
rect 24334 21586 24386 21598
rect 14354 21534 14366 21586
rect 14418 21534 14430 21586
rect 16818 21534 16830 21586
rect 16882 21534 16894 21586
rect 17490 21534 17502 21586
rect 17554 21534 17566 21586
rect 18274 21534 18286 21586
rect 18338 21534 18350 21586
rect 26226 21534 26238 21586
rect 26290 21534 26302 21586
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 24334 21522 24386 21534
rect 13470 21474 13522 21486
rect 15150 21474 15202 21486
rect 14018 21422 14030 21474
rect 14082 21422 14094 21474
rect 13470 21410 13522 21422
rect 15150 21410 15202 21422
rect 25342 21474 25394 21486
rect 25342 21410 25394 21422
rect 25902 21474 25954 21486
rect 40014 21474 40066 21486
rect 29138 21422 29150 21474
rect 29202 21422 29214 21474
rect 25902 21410 25954 21422
rect 40014 21410 40066 21422
rect 23998 21362 24050 21374
rect 23998 21298 24050 21310
rect 24222 21362 24274 21374
rect 25330 21310 25342 21362
rect 25394 21359 25406 21362
rect 25890 21359 25902 21362
rect 25394 21313 25902 21359
rect 25394 21310 25406 21313
rect 25890 21310 25902 21313
rect 25954 21310 25966 21362
rect 24222 21298 24274 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 22542 20914 22594 20926
rect 40014 20914 40066 20926
rect 28578 20862 28590 20914
rect 28642 20862 28654 20914
rect 22542 20850 22594 20862
rect 40014 20850 40066 20862
rect 14142 20802 14194 20814
rect 14142 20738 14194 20750
rect 14702 20802 14754 20814
rect 24446 20802 24498 20814
rect 20290 20750 20302 20802
rect 20354 20750 20366 20802
rect 21298 20750 21310 20802
rect 21362 20750 21374 20802
rect 23202 20750 23214 20802
rect 23266 20750 23278 20802
rect 14702 20738 14754 20750
rect 24446 20738 24498 20750
rect 25006 20802 25058 20814
rect 25778 20750 25790 20802
rect 25842 20750 25854 20802
rect 37650 20750 37662 20802
rect 37714 20750 37726 20802
rect 25006 20738 25058 20750
rect 22430 20690 22482 20702
rect 16818 20638 16830 20690
rect 16882 20638 16894 20690
rect 22430 20626 22482 20638
rect 22654 20690 22706 20702
rect 22654 20626 22706 20638
rect 22766 20690 22818 20702
rect 24110 20690 24162 20702
rect 23874 20638 23886 20690
rect 23938 20638 23950 20690
rect 25330 20638 25342 20690
rect 25394 20638 25406 20690
rect 26450 20638 26462 20690
rect 26514 20638 26526 20690
rect 22766 20626 22818 20638
rect 24110 20626 24162 20638
rect 21646 20578 21698 20590
rect 21646 20514 21698 20526
rect 21758 20578 21810 20590
rect 21758 20514 21810 20526
rect 21870 20578 21922 20590
rect 21870 20514 21922 20526
rect 23550 20578 23602 20590
rect 23550 20514 23602 20526
rect 24334 20578 24386 20590
rect 24334 20514 24386 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 14702 20242 14754 20254
rect 14702 20178 14754 20190
rect 18958 20242 19010 20254
rect 18958 20178 19010 20190
rect 26350 20242 26402 20254
rect 26350 20178 26402 20190
rect 14142 20130 14194 20142
rect 18846 20130 18898 20142
rect 15026 20078 15038 20130
rect 15090 20078 15102 20130
rect 15698 20078 15710 20130
rect 15762 20078 15774 20130
rect 14142 20066 14194 20078
rect 18846 20066 18898 20078
rect 19070 20130 19122 20142
rect 19070 20066 19122 20078
rect 21086 20130 21138 20142
rect 21086 20066 21138 20078
rect 22654 20130 22706 20142
rect 22654 20066 22706 20078
rect 24222 20130 24274 20142
rect 25902 20130 25954 20142
rect 27918 20130 27970 20142
rect 24546 20078 24558 20130
rect 24610 20078 24622 20130
rect 26226 20078 26238 20130
rect 26290 20078 26302 20130
rect 24222 20066 24274 20078
rect 25902 20066 25954 20078
rect 27918 20066 27970 20078
rect 13246 20018 13298 20030
rect 9986 19966 9998 20018
rect 10050 19966 10062 20018
rect 13246 19954 13298 19966
rect 13694 20018 13746 20030
rect 13694 19954 13746 19966
rect 13918 20018 13970 20030
rect 17390 20018 17442 20030
rect 15474 19966 15486 20018
rect 15538 19966 15550 20018
rect 16258 19966 16270 20018
rect 16322 19966 16334 20018
rect 16706 19966 16718 20018
rect 16770 19966 16782 20018
rect 13918 19954 13970 19966
rect 17390 19954 17442 19966
rect 17950 20018 18002 20030
rect 21198 20018 21250 20030
rect 25566 20018 25618 20030
rect 19842 19966 19854 20018
rect 19906 19966 19918 20018
rect 20066 19966 20078 20018
rect 20130 19966 20142 20018
rect 22082 19966 22094 20018
rect 22146 19966 22158 20018
rect 22866 19966 22878 20018
rect 22930 19966 22942 20018
rect 17950 19954 18002 19966
rect 21198 19954 21250 19966
rect 25566 19954 25618 19966
rect 26462 20018 26514 20030
rect 26462 19954 26514 19966
rect 27806 20018 27858 20030
rect 27806 19954 27858 19966
rect 14030 19906 14082 19918
rect 25678 19906 25730 19918
rect 10658 19854 10670 19906
rect 10722 19854 10734 19906
rect 12786 19854 12798 19906
rect 12850 19854 12862 19906
rect 19954 19854 19966 19906
rect 20018 19854 20030 19906
rect 21970 19854 21982 19906
rect 22034 19854 22046 19906
rect 23090 19854 23102 19906
rect 23154 19854 23166 19906
rect 14030 19842 14082 19854
rect 25678 19842 25730 19854
rect 16706 19742 16718 19794
rect 16770 19742 16782 19794
rect 20626 19742 20638 19794
rect 20690 19742 20702 19794
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 16382 19458 16434 19470
rect 16382 19394 16434 19406
rect 16718 19458 16770 19470
rect 21310 19458 21362 19470
rect 18610 19406 18622 19458
rect 18674 19406 18686 19458
rect 16718 19394 16770 19406
rect 21310 19394 21362 19406
rect 21870 19458 21922 19470
rect 21870 19394 21922 19406
rect 22094 19458 22146 19470
rect 22094 19394 22146 19406
rect 14030 19346 14082 19358
rect 14030 19282 14082 19294
rect 19182 19346 19234 19358
rect 19618 19294 19630 19346
rect 19682 19294 19694 19346
rect 19182 19282 19234 19294
rect 14142 19234 14194 19246
rect 14142 19170 14194 19182
rect 14478 19234 14530 19246
rect 15710 19234 15762 19246
rect 15362 19182 15374 19234
rect 15426 19182 15438 19234
rect 14478 19170 14530 19182
rect 15710 19170 15762 19182
rect 16046 19234 16098 19246
rect 16046 19170 16098 19182
rect 18958 19234 19010 19246
rect 20862 19234 20914 19246
rect 19842 19182 19854 19234
rect 19906 19182 19918 19234
rect 20178 19182 20190 19234
rect 20242 19182 20254 19234
rect 18958 19170 19010 19182
rect 20862 19170 20914 19182
rect 21422 19234 21474 19246
rect 21422 19170 21474 19182
rect 26126 19234 26178 19246
rect 26126 19170 26178 19182
rect 16494 19122 16546 19134
rect 14802 19070 14814 19122
rect 14866 19070 14878 19122
rect 16494 19058 16546 19070
rect 26462 19122 26514 19134
rect 26562 19070 26574 19122
rect 26626 19070 26638 19122
rect 26462 19058 26514 19070
rect 15934 19010 15986 19022
rect 15138 18958 15150 19010
rect 15202 18958 15214 19010
rect 15934 18946 15986 18958
rect 22206 19010 22258 19022
rect 22206 18946 22258 18958
rect 22542 19010 22594 19022
rect 26238 19010 26290 19022
rect 22866 18958 22878 19010
rect 22930 18958 22942 19010
rect 22542 18946 22594 18958
rect 26238 18946 26290 18958
rect 26350 19010 26402 19022
rect 26350 18946 26402 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 13470 18674 13522 18686
rect 12562 18622 12574 18674
rect 12626 18622 12638 18674
rect 13470 18610 13522 18622
rect 19182 18674 19234 18686
rect 19182 18610 19234 18622
rect 19406 18674 19458 18686
rect 22642 18622 22654 18674
rect 22706 18622 22718 18674
rect 19406 18610 19458 18622
rect 20290 18510 20302 18562
rect 20354 18510 20366 18562
rect 22194 18510 22206 18562
rect 22258 18510 22270 18562
rect 26562 18510 26574 18562
rect 26626 18510 26638 18562
rect 11678 18450 11730 18462
rect 4274 18398 4286 18450
rect 4338 18398 4350 18450
rect 11678 18386 11730 18398
rect 13134 18450 13186 18462
rect 13134 18386 13186 18398
rect 13694 18450 13746 18462
rect 13694 18386 13746 18398
rect 14142 18450 14194 18462
rect 14142 18386 14194 18398
rect 18846 18450 18898 18462
rect 22990 18450 23042 18462
rect 21186 18398 21198 18450
rect 21250 18398 21262 18450
rect 21410 18398 21422 18450
rect 21474 18398 21486 18450
rect 25778 18398 25790 18450
rect 25842 18398 25854 18450
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 18846 18386 18898 18398
rect 22990 18386 23042 18398
rect 12910 18338 12962 18350
rect 12910 18274 12962 18286
rect 13582 18338 13634 18350
rect 13582 18274 13634 18286
rect 24670 18338 24722 18350
rect 24670 18274 24722 18286
rect 25230 18338 25282 18350
rect 28690 18286 28702 18338
rect 28754 18286 28766 18338
rect 25230 18274 25282 18286
rect 1934 18226 1986 18238
rect 1934 18162 1986 18174
rect 11790 18226 11842 18238
rect 11790 18162 11842 18174
rect 19070 18226 19122 18238
rect 19070 18162 19122 18174
rect 25342 18226 25394 18238
rect 25342 18162 25394 18174
rect 40014 18226 40066 18238
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 27694 17890 27746 17902
rect 21858 17838 21870 17890
rect 21922 17838 21934 17890
rect 27694 17826 27746 17838
rect 1934 17778 1986 17790
rect 27806 17778 27858 17790
rect 9874 17726 9886 17778
rect 9938 17726 9950 17778
rect 12002 17726 12014 17778
rect 12066 17726 12078 17778
rect 26114 17726 26126 17778
rect 26178 17726 26190 17778
rect 1934 17714 1986 17726
rect 27806 17714 27858 17726
rect 40014 17778 40066 17790
rect 40014 17714 40066 17726
rect 15262 17666 15314 17678
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 12674 17614 12686 17666
rect 12738 17614 12750 17666
rect 13682 17614 13694 17666
rect 13746 17614 13758 17666
rect 15262 17602 15314 17614
rect 16158 17666 16210 17678
rect 16158 17602 16210 17614
rect 16494 17666 16546 17678
rect 16494 17602 16546 17614
rect 17726 17666 17778 17678
rect 21310 17666 21362 17678
rect 26462 17666 26514 17678
rect 20066 17614 20078 17666
rect 20130 17614 20142 17666
rect 20402 17614 20414 17666
rect 20466 17614 20478 17666
rect 21522 17614 21534 17666
rect 21586 17614 21598 17666
rect 21858 17614 21870 17666
rect 21922 17614 21934 17666
rect 25666 17614 25678 17666
rect 25730 17614 25742 17666
rect 17726 17602 17778 17614
rect 21310 17602 21362 17614
rect 26462 17602 26514 17614
rect 27134 17666 27186 17678
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 27134 17602 27186 17614
rect 15150 17554 15202 17566
rect 26126 17554 26178 17566
rect 13458 17502 13470 17554
rect 13522 17502 13534 17554
rect 16818 17502 16830 17554
rect 16882 17502 16894 17554
rect 18050 17502 18062 17554
rect 18114 17502 18126 17554
rect 15150 17490 15202 17502
rect 26126 17490 26178 17502
rect 26238 17554 26290 17566
rect 26238 17490 26290 17502
rect 14926 17442 14978 17454
rect 14926 17378 14978 17390
rect 15822 17442 15874 17454
rect 15822 17378 15874 17390
rect 16046 17442 16098 17454
rect 16046 17378 16098 17390
rect 19854 17442 19906 17454
rect 27022 17442 27074 17454
rect 21746 17390 21758 17442
rect 21810 17390 21822 17442
rect 19854 17378 19906 17390
rect 27022 17378 27074 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 13022 17106 13074 17118
rect 13022 17042 13074 17054
rect 14702 17106 14754 17118
rect 21646 17106 21698 17118
rect 20402 17054 20414 17106
rect 20466 17054 20478 17106
rect 14702 17042 14754 17054
rect 21646 17042 21698 17054
rect 14926 16994 14978 17006
rect 14926 16930 14978 16942
rect 15038 16994 15090 17006
rect 26002 16942 26014 16994
rect 26066 16942 26078 16994
rect 15038 16930 15090 16942
rect 20750 16882 20802 16894
rect 4274 16830 4286 16882
rect 4338 16830 4350 16882
rect 15474 16830 15486 16882
rect 15538 16830 15550 16882
rect 15810 16830 15822 16882
rect 15874 16830 15886 16882
rect 20750 16818 20802 16830
rect 21086 16882 21138 16894
rect 28590 16882 28642 16894
rect 22754 16830 22766 16882
rect 22818 16830 22830 16882
rect 22978 16830 22990 16882
rect 23042 16830 23054 16882
rect 25218 16830 25230 16882
rect 25282 16830 25294 16882
rect 21086 16818 21138 16830
rect 28590 16818 28642 16830
rect 14814 16770 14866 16782
rect 14814 16706 14866 16718
rect 16158 16770 16210 16782
rect 16158 16706 16210 16718
rect 23214 16770 23266 16782
rect 28130 16718 28142 16770
rect 28194 16718 28206 16770
rect 23214 16706 23266 16718
rect 1934 16658 1986 16670
rect 1934 16594 1986 16606
rect 15822 16658 15874 16670
rect 15822 16594 15874 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 20750 16210 20802 16222
rect 20514 16158 20526 16210
rect 20578 16158 20590 16210
rect 21858 16158 21870 16210
rect 21922 16158 21934 16210
rect 23986 16158 23998 16210
rect 24050 16158 24062 16210
rect 20750 16146 20802 16158
rect 14814 16098 14866 16110
rect 14814 16034 14866 16046
rect 15038 16098 15090 16110
rect 15038 16034 15090 16046
rect 15374 16098 15426 16110
rect 15374 16034 15426 16046
rect 17614 16098 17666 16110
rect 25230 16098 25282 16110
rect 24770 16046 24782 16098
rect 24834 16046 24846 16098
rect 17614 16034 17666 16046
rect 25230 16034 25282 16046
rect 14926 15874 14978 15886
rect 14926 15810 14978 15822
rect 17726 15874 17778 15886
rect 17726 15810 17778 15822
rect 17950 15874 18002 15886
rect 17950 15810 18002 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 23774 15538 23826 15550
rect 23774 15474 23826 15486
rect 16046 15426 16098 15438
rect 13682 15374 13694 15426
rect 13746 15374 13758 15426
rect 16046 15362 16098 15374
rect 16158 15426 16210 15438
rect 16158 15362 16210 15374
rect 17390 15426 17442 15438
rect 17390 15362 17442 15374
rect 17614 15426 17666 15438
rect 17614 15362 17666 15374
rect 17950 15426 18002 15438
rect 17950 15362 18002 15374
rect 18398 15426 18450 15438
rect 23438 15426 23490 15438
rect 20962 15374 20974 15426
rect 21026 15374 21038 15426
rect 18398 15362 18450 15374
rect 23438 15362 23490 15374
rect 15150 15314 15202 15326
rect 14354 15262 14366 15314
rect 14418 15262 14430 15314
rect 15150 15250 15202 15262
rect 15374 15314 15426 15326
rect 15374 15250 15426 15262
rect 15598 15314 15650 15326
rect 15598 15250 15650 15262
rect 15822 15314 15874 15326
rect 15822 15250 15874 15262
rect 18734 15314 18786 15326
rect 18734 15250 18786 15262
rect 19070 15314 19122 15326
rect 24222 15314 24274 15326
rect 20290 15262 20302 15314
rect 20354 15262 20366 15314
rect 19070 15250 19122 15262
rect 24222 15250 24274 15262
rect 15486 15202 15538 15214
rect 11554 15150 11566 15202
rect 11618 15150 11630 15202
rect 15486 15138 15538 15150
rect 17838 15202 17890 15214
rect 17838 15138 17890 15150
rect 18846 15202 18898 15214
rect 23090 15150 23102 15202
rect 23154 15150 23166 15202
rect 18846 15138 18898 15150
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 19070 14754 19122 14766
rect 19070 14690 19122 14702
rect 14702 14642 14754 14654
rect 16370 14590 16382 14642
rect 16434 14590 16446 14642
rect 18498 14590 18510 14642
rect 18562 14590 18574 14642
rect 14702 14578 14754 14590
rect 19182 14530 19234 14542
rect 15586 14478 15598 14530
rect 15650 14478 15662 14530
rect 19182 14466 19234 14478
rect 19070 14306 19122 14318
rect 19070 14242 19122 14254
rect 19630 14306 19682 14318
rect 19630 14242 19682 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 16382 13970 16434 13982
rect 16382 13906 16434 13918
rect 16830 13970 16882 13982
rect 16830 13906 16882 13918
rect 13794 13806 13806 13858
rect 13858 13806 13870 13858
rect 18274 13806 18286 13858
rect 18338 13806 18350 13858
rect 20738 13806 20750 13858
rect 20802 13806 20814 13858
rect 13010 13694 13022 13746
rect 13074 13694 13086 13746
rect 17490 13694 17502 13746
rect 17554 13694 17566 13746
rect 20962 13694 20974 13746
rect 21026 13694 21038 13746
rect 15922 13582 15934 13634
rect 15986 13582 15998 13634
rect 20402 13582 20414 13634
rect 20466 13582 20478 13634
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 19854 12738 19906 12750
rect 20178 12686 20190 12738
rect 20242 12686 20254 12738
rect 19854 12674 19906 12686
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 40238 11170 40290 11182
rect 40238 11106 40290 11118
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 17390 5234 17442 5246
rect 17390 5170 17442 5182
rect 16370 5070 16382 5122
rect 16434 5070 16446 5122
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 17602 4286 17614 4338
rect 17666 4286 17678 4338
rect 20402 4286 20414 4338
rect 20466 4286 20478 4338
rect 18510 4114 18562 4126
rect 18510 4050 18562 4062
rect 21422 4114 21474 4126
rect 21422 4050 21474 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 22094 3666 22146 3678
rect 22094 3602 22146 3614
rect 19730 3502 19742 3554
rect 19794 3502 19806 3554
rect 21074 3502 21086 3554
rect 21138 3502 21150 3554
rect 19182 3330 19234 3342
rect 19182 3266 19234 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 26910 38558 26962 38610
rect 28366 38558 28418 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 19518 38222 19570 38274
rect 22430 38222 22482 38274
rect 25566 38222 25618 38274
rect 17838 37998 17890 38050
rect 21758 37998 21810 38050
rect 24558 37998 24610 38050
rect 27470 37886 27522 37938
rect 28366 37886 28418 37938
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 19070 37438 19122 37490
rect 21422 37438 21474 37490
rect 26798 37438 26850 37490
rect 19630 37214 19682 37266
rect 20638 37214 20690 37266
rect 25790 37214 25842 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 17390 36654 17442 36706
rect 16606 36430 16658 36482
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 18958 29374 19010 29426
rect 22318 29374 22370 29426
rect 19630 29262 19682 29314
rect 21758 29262 21810 29314
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19182 28702 19234 28754
rect 16382 28590 16434 28642
rect 17054 28478 17106 28530
rect 19630 28478 19682 28530
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 17390 28030 17442 28082
rect 19070 28030 19122 28082
rect 19854 28030 19906 28082
rect 20750 28030 20802 28082
rect 17614 27918 17666 27970
rect 20078 27918 20130 27970
rect 14814 27806 14866 27858
rect 17726 27806 17778 27858
rect 18846 27806 18898 27858
rect 19182 27806 19234 27858
rect 20190 27806 20242 27858
rect 20526 27806 20578 27858
rect 20862 27806 20914 27858
rect 21758 27806 21810 27858
rect 12014 27694 12066 27746
rect 14142 27694 14194 27746
rect 15374 27694 15426 27746
rect 22430 27694 22482 27746
rect 24558 27694 24610 27746
rect 25342 27694 25394 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 22542 27246 22594 27298
rect 22430 27022 22482 27074
rect 23326 27022 23378 27074
rect 18846 26910 18898 26962
rect 18958 26910 19010 26962
rect 22542 26910 22594 26962
rect 22990 26910 23042 26962
rect 23214 26910 23266 26962
rect 19182 26798 19234 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 25342 26350 25394 26402
rect 4286 26238 4338 26290
rect 13582 26238 13634 26290
rect 20302 26238 20354 26290
rect 14254 26126 14306 26178
rect 16382 26126 16434 26178
rect 16830 26126 16882 26178
rect 17390 26126 17442 26178
rect 19518 26126 19570 26178
rect 20750 26126 20802 26178
rect 1934 26014 1986 26066
rect 25230 26014 25282 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 15822 25678 15874 25730
rect 21646 25678 21698 25730
rect 14478 25566 14530 25618
rect 19518 25566 19570 25618
rect 25678 25566 25730 25618
rect 40014 25566 40066 25618
rect 14926 25454 14978 25506
rect 15150 25454 15202 25506
rect 19182 25454 19234 25506
rect 22878 25454 22930 25506
rect 37662 25454 37714 25506
rect 14366 25342 14418 25394
rect 15374 25342 15426 25394
rect 15486 25342 15538 25394
rect 15934 25342 15986 25394
rect 19742 25342 19794 25394
rect 21534 25342 21586 25394
rect 22094 25342 22146 25394
rect 22430 25342 22482 25394
rect 23550 25342 23602 25394
rect 26126 25342 26178 25394
rect 26238 25342 26290 25394
rect 14590 25230 14642 25282
rect 19518 25230 19570 25282
rect 21646 25230 21698 25282
rect 26462 25230 26514 25282
rect 26798 25230 26850 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 16046 24894 16098 24946
rect 16158 24894 16210 24946
rect 17726 24894 17778 24946
rect 20190 24894 20242 24946
rect 21758 24894 21810 24946
rect 23326 24894 23378 24946
rect 28590 24894 28642 24946
rect 20526 24782 20578 24834
rect 21534 24782 21586 24834
rect 23438 24782 23490 24834
rect 4286 24670 4338 24722
rect 13470 24670 13522 24722
rect 13918 24670 13970 24722
rect 16382 24670 16434 24722
rect 16606 24670 16658 24722
rect 17390 24670 17442 24722
rect 20078 24670 20130 24722
rect 20302 24670 20354 24722
rect 21198 24670 21250 24722
rect 22430 24670 22482 24722
rect 22766 24670 22818 24722
rect 25342 24670 25394 24722
rect 10558 24558 10610 24610
rect 12686 24558 12738 24610
rect 16046 24558 16098 24610
rect 21646 24558 21698 24610
rect 22990 24558 23042 24610
rect 23214 24558 23266 24610
rect 26014 24558 26066 24610
rect 28142 24558 28194 24610
rect 1934 24446 1986 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 12462 24110 12514 24162
rect 13806 23998 13858 24050
rect 20190 23998 20242 24050
rect 25566 23998 25618 24050
rect 12350 23886 12402 23938
rect 13694 23886 13746 23938
rect 13918 23886 13970 23938
rect 17278 23886 17330 23938
rect 25678 23886 25730 23938
rect 26126 23886 26178 23938
rect 14366 23774 14418 23826
rect 18062 23774 18114 23826
rect 14142 23662 14194 23714
rect 16942 23662 16994 23714
rect 25454 23662 25506 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 19406 23326 19458 23378
rect 19518 23326 19570 23378
rect 19630 23326 19682 23378
rect 19966 23326 20018 23378
rect 13694 23214 13746 23266
rect 18174 23214 18226 23266
rect 20190 23214 20242 23266
rect 26574 23214 26626 23266
rect 26686 23214 26738 23266
rect 26798 23214 26850 23266
rect 13358 23102 13410 23154
rect 16270 23102 16322 23154
rect 16494 23102 16546 23154
rect 16830 23102 16882 23154
rect 18510 23102 18562 23154
rect 19070 23102 19122 23154
rect 19294 23102 19346 23154
rect 20302 23102 20354 23154
rect 20862 23102 20914 23154
rect 21198 23102 21250 23154
rect 21310 23102 21362 23154
rect 24670 23102 24722 23154
rect 26350 23102 26402 23154
rect 16382 22990 16434 23042
rect 20974 22990 21026 23042
rect 21758 22990 21810 23042
rect 23886 22990 23938 23042
rect 25342 22990 25394 23042
rect 26686 22990 26738 23042
rect 18286 22878 18338 22930
rect 18622 22878 18674 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 17502 22542 17554 22594
rect 19182 22542 19234 22594
rect 19294 22542 19346 22594
rect 28142 22542 28194 22594
rect 10670 22430 10722 22482
rect 12798 22430 12850 22482
rect 40014 22430 40066 22482
rect 9998 22318 10050 22370
rect 14030 22318 14082 22370
rect 17614 22318 17666 22370
rect 18734 22318 18786 22370
rect 18958 22318 19010 22370
rect 19630 22318 19682 22370
rect 21870 22318 21922 22370
rect 37662 22318 37714 22370
rect 14366 22206 14418 22258
rect 15262 22206 15314 22258
rect 18174 22206 18226 22258
rect 19742 22206 19794 22258
rect 20414 22206 20466 22258
rect 26238 22206 26290 22258
rect 28254 22206 28306 22258
rect 13582 22094 13634 22146
rect 15598 22094 15650 22146
rect 17054 22094 17106 22146
rect 17502 22094 17554 22146
rect 18286 22094 18338 22146
rect 18510 22094 18562 22146
rect 20638 22094 20690 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 12910 21758 12962 21810
rect 15262 21758 15314 21810
rect 15822 21758 15874 21810
rect 16606 21758 16658 21810
rect 14814 21646 14866 21698
rect 15710 21646 15762 21698
rect 15934 21646 15986 21698
rect 16494 21646 16546 21698
rect 17726 21646 17778 21698
rect 21758 21646 21810 21698
rect 23886 21646 23938 21698
rect 27022 21646 27074 21698
rect 14366 21534 14418 21586
rect 16830 21534 16882 21586
rect 17502 21534 17554 21586
rect 18286 21534 18338 21586
rect 24334 21534 24386 21586
rect 26238 21534 26290 21586
rect 37662 21534 37714 21586
rect 13470 21422 13522 21474
rect 14030 21422 14082 21474
rect 15150 21422 15202 21474
rect 25342 21422 25394 21474
rect 25902 21422 25954 21474
rect 29150 21422 29202 21474
rect 40014 21422 40066 21474
rect 23998 21310 24050 21362
rect 24222 21310 24274 21362
rect 25342 21310 25394 21362
rect 25902 21310 25954 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 22542 20862 22594 20914
rect 28590 20862 28642 20914
rect 40014 20862 40066 20914
rect 14142 20750 14194 20802
rect 14702 20750 14754 20802
rect 20302 20750 20354 20802
rect 21310 20750 21362 20802
rect 23214 20750 23266 20802
rect 24446 20750 24498 20802
rect 25006 20750 25058 20802
rect 25790 20750 25842 20802
rect 37662 20750 37714 20802
rect 16830 20638 16882 20690
rect 22430 20638 22482 20690
rect 22654 20638 22706 20690
rect 22766 20638 22818 20690
rect 23886 20638 23938 20690
rect 24110 20638 24162 20690
rect 25342 20638 25394 20690
rect 26462 20638 26514 20690
rect 21646 20526 21698 20578
rect 21758 20526 21810 20578
rect 21870 20526 21922 20578
rect 23550 20526 23602 20578
rect 24334 20526 24386 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 14702 20190 14754 20242
rect 18958 20190 19010 20242
rect 26350 20190 26402 20242
rect 14142 20078 14194 20130
rect 15038 20078 15090 20130
rect 15710 20078 15762 20130
rect 18846 20078 18898 20130
rect 19070 20078 19122 20130
rect 21086 20078 21138 20130
rect 22654 20078 22706 20130
rect 24222 20078 24274 20130
rect 24558 20078 24610 20130
rect 25902 20078 25954 20130
rect 26238 20078 26290 20130
rect 27918 20078 27970 20130
rect 9998 19966 10050 20018
rect 13246 19966 13298 20018
rect 13694 19966 13746 20018
rect 13918 19966 13970 20018
rect 15486 19966 15538 20018
rect 16270 19966 16322 20018
rect 16718 19966 16770 20018
rect 17390 19966 17442 20018
rect 17950 19966 18002 20018
rect 19854 19966 19906 20018
rect 20078 19966 20130 20018
rect 21198 19966 21250 20018
rect 22094 19966 22146 20018
rect 22878 19966 22930 20018
rect 25566 19966 25618 20018
rect 26462 19966 26514 20018
rect 27806 19966 27858 20018
rect 10670 19854 10722 19906
rect 12798 19854 12850 19906
rect 14030 19854 14082 19906
rect 19966 19854 20018 19906
rect 21982 19854 22034 19906
rect 23102 19854 23154 19906
rect 25678 19854 25730 19906
rect 16718 19742 16770 19794
rect 20638 19742 20690 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 16382 19406 16434 19458
rect 16718 19406 16770 19458
rect 18622 19406 18674 19458
rect 21310 19406 21362 19458
rect 21870 19406 21922 19458
rect 22094 19406 22146 19458
rect 14030 19294 14082 19346
rect 19182 19294 19234 19346
rect 19630 19294 19682 19346
rect 14142 19182 14194 19234
rect 14478 19182 14530 19234
rect 15374 19182 15426 19234
rect 15710 19182 15762 19234
rect 16046 19182 16098 19234
rect 18958 19182 19010 19234
rect 19854 19182 19906 19234
rect 20190 19182 20242 19234
rect 20862 19182 20914 19234
rect 21422 19182 21474 19234
rect 26126 19182 26178 19234
rect 14814 19070 14866 19122
rect 16494 19070 16546 19122
rect 26462 19070 26514 19122
rect 26574 19070 26626 19122
rect 15150 18958 15202 19010
rect 15934 18958 15986 19010
rect 22206 18958 22258 19010
rect 22542 18958 22594 19010
rect 22878 18958 22930 19010
rect 26238 18958 26290 19010
rect 26350 18958 26402 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 12574 18622 12626 18674
rect 13470 18622 13522 18674
rect 19182 18622 19234 18674
rect 19406 18622 19458 18674
rect 22654 18622 22706 18674
rect 20302 18510 20354 18562
rect 22206 18510 22258 18562
rect 26574 18510 26626 18562
rect 4286 18398 4338 18450
rect 11678 18398 11730 18450
rect 13134 18398 13186 18450
rect 13694 18398 13746 18450
rect 14142 18398 14194 18450
rect 18846 18398 18898 18450
rect 21198 18398 21250 18450
rect 21422 18398 21474 18450
rect 22990 18398 23042 18450
rect 25790 18398 25842 18450
rect 37662 18398 37714 18450
rect 12910 18286 12962 18338
rect 13582 18286 13634 18338
rect 24670 18286 24722 18338
rect 25230 18286 25282 18338
rect 28702 18286 28754 18338
rect 1934 18174 1986 18226
rect 11790 18174 11842 18226
rect 19070 18174 19122 18226
rect 25342 18174 25394 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 21870 17838 21922 17890
rect 27694 17838 27746 17890
rect 1934 17726 1986 17778
rect 9886 17726 9938 17778
rect 12014 17726 12066 17778
rect 26126 17726 26178 17778
rect 27806 17726 27858 17778
rect 40014 17726 40066 17778
rect 4286 17614 4338 17666
rect 12686 17614 12738 17666
rect 13694 17614 13746 17666
rect 15262 17614 15314 17666
rect 16158 17614 16210 17666
rect 16494 17614 16546 17666
rect 17726 17614 17778 17666
rect 20078 17614 20130 17666
rect 20414 17614 20466 17666
rect 21310 17614 21362 17666
rect 21534 17614 21586 17666
rect 21870 17614 21922 17666
rect 25678 17614 25730 17666
rect 26462 17614 26514 17666
rect 27134 17614 27186 17666
rect 37662 17614 37714 17666
rect 13470 17502 13522 17554
rect 15150 17502 15202 17554
rect 16830 17502 16882 17554
rect 18062 17502 18114 17554
rect 26126 17502 26178 17554
rect 26238 17502 26290 17554
rect 14926 17390 14978 17442
rect 15822 17390 15874 17442
rect 16046 17390 16098 17442
rect 19854 17390 19906 17442
rect 21758 17390 21810 17442
rect 27022 17390 27074 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 13022 17054 13074 17106
rect 14702 17054 14754 17106
rect 20414 17054 20466 17106
rect 21646 17054 21698 17106
rect 14926 16942 14978 16994
rect 15038 16942 15090 16994
rect 26014 16942 26066 16994
rect 4286 16830 4338 16882
rect 15486 16830 15538 16882
rect 15822 16830 15874 16882
rect 20750 16830 20802 16882
rect 21086 16830 21138 16882
rect 22766 16830 22818 16882
rect 22990 16830 23042 16882
rect 25230 16830 25282 16882
rect 28590 16830 28642 16882
rect 14814 16718 14866 16770
rect 16158 16718 16210 16770
rect 23214 16718 23266 16770
rect 28142 16718 28194 16770
rect 1934 16606 1986 16658
rect 15822 16606 15874 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 20526 16158 20578 16210
rect 20750 16158 20802 16210
rect 21870 16158 21922 16210
rect 23998 16158 24050 16210
rect 14814 16046 14866 16098
rect 15038 16046 15090 16098
rect 15374 16046 15426 16098
rect 17614 16046 17666 16098
rect 24782 16046 24834 16098
rect 25230 16046 25282 16098
rect 14926 15822 14978 15874
rect 17726 15822 17778 15874
rect 17950 15822 18002 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 23774 15486 23826 15538
rect 13694 15374 13746 15426
rect 16046 15374 16098 15426
rect 16158 15374 16210 15426
rect 17390 15374 17442 15426
rect 17614 15374 17666 15426
rect 17950 15374 18002 15426
rect 18398 15374 18450 15426
rect 20974 15374 21026 15426
rect 23438 15374 23490 15426
rect 14366 15262 14418 15314
rect 15150 15262 15202 15314
rect 15374 15262 15426 15314
rect 15598 15262 15650 15314
rect 15822 15262 15874 15314
rect 18734 15262 18786 15314
rect 19070 15262 19122 15314
rect 20302 15262 20354 15314
rect 24222 15262 24274 15314
rect 11566 15150 11618 15202
rect 15486 15150 15538 15202
rect 17838 15150 17890 15202
rect 18846 15150 18898 15202
rect 23102 15150 23154 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 19070 14702 19122 14754
rect 14702 14590 14754 14642
rect 16382 14590 16434 14642
rect 18510 14590 18562 14642
rect 15598 14478 15650 14530
rect 19182 14478 19234 14530
rect 19070 14254 19122 14306
rect 19630 14254 19682 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 16382 13918 16434 13970
rect 16830 13918 16882 13970
rect 13806 13806 13858 13858
rect 18286 13806 18338 13858
rect 20750 13806 20802 13858
rect 13022 13694 13074 13746
rect 17502 13694 17554 13746
rect 20974 13694 21026 13746
rect 15934 13582 15986 13634
rect 20414 13582 20466 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 19854 12686 19906 12738
rect 20190 12686 20242 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 40238 11118 40290 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 17390 5182 17442 5234
rect 16382 5070 16434 5122
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 17614 4286 17666 4338
rect 20414 4286 20466 4338
rect 18510 4062 18562 4114
rect 21422 4062 21474 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 22094 3614 22146 3666
rect 19742 3502 19794 3554
rect 21086 3502 21138 3554
rect 19182 3278 19234 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 16128 41200 16240 42000
rect 18816 41200 18928 42000
rect 19488 41200 19600 42000
rect 20160 41200 20272 42000
rect 21504 41200 21616 42000
rect 24192 41200 24304 42000
rect 25536 41200 25648 42000
rect 26208 41200 26320 42000
rect 26880 41200 26992 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 16156 36708 16212 41200
rect 18844 38668 18900 41200
rect 18844 38612 19124 38668
rect 17836 38050 17892 38062
rect 17836 37998 17838 38050
rect 17890 37998 17892 38050
rect 16156 36642 16212 36652
rect 17388 36708 17444 36718
rect 17388 36614 17444 36652
rect 16604 36482 16660 36494
rect 16604 36430 16606 36482
rect 16658 36430 16660 36482
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 16380 28642 16436 28654
rect 16380 28590 16382 28642
rect 16434 28590 16436 28642
rect 16380 28532 16436 28590
rect 16380 28466 16436 28476
rect 4172 28308 4228 28318
rect 1932 26066 1988 26078
rect 1932 26014 1934 26066
rect 1986 26014 1988 26066
rect 1932 25620 1988 26014
rect 1932 25554 1988 25564
rect 1932 24500 1988 24510
rect 1932 24406 1988 24444
rect 4172 22148 4228 28252
rect 14812 27858 14868 27870
rect 14812 27806 14814 27858
rect 14866 27806 14868 27858
rect 12012 27746 12068 27758
rect 12012 27694 12014 27746
rect 12066 27694 12068 27746
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4284 26292 4340 26302
rect 4284 26198 4340 26236
rect 12012 26292 12068 27694
rect 14140 27748 14196 27758
rect 14812 27748 14868 27806
rect 15372 27748 15428 27758
rect 14140 27746 14532 27748
rect 14140 27694 14142 27746
rect 14194 27694 14532 27746
rect 14140 27692 14532 27694
rect 14140 27682 14196 27692
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 12012 25396 12068 26236
rect 12012 25330 12068 25340
rect 13580 26964 13636 26974
rect 13580 26290 13636 26908
rect 13580 26238 13582 26290
rect 13634 26238 13636 26290
rect 4284 24724 4340 24734
rect 4284 24630 4340 24668
rect 13468 24724 13524 24734
rect 13580 24724 13636 26238
rect 14252 26180 14308 26190
rect 14252 26086 14308 26124
rect 14476 25618 14532 27692
rect 14812 27746 15428 27748
rect 14812 27694 15374 27746
rect 15426 27694 15428 27746
rect 14812 27692 15428 27694
rect 14812 26964 14868 27692
rect 15372 27682 15428 27692
rect 16604 26908 16660 36430
rect 14812 26898 14868 26908
rect 16380 26852 16660 26908
rect 16828 28532 16884 28542
rect 15820 26180 15876 26190
rect 15820 25730 15876 26124
rect 15820 25678 15822 25730
rect 15874 25678 15876 25730
rect 15820 25666 15876 25678
rect 16380 26178 16436 26852
rect 16380 26126 16382 26178
rect 16434 26126 16436 26178
rect 14476 25566 14478 25618
rect 14530 25566 14532 25618
rect 14476 25554 14532 25566
rect 14924 25508 14980 25518
rect 15148 25508 15204 25518
rect 14924 25506 15204 25508
rect 14924 25454 14926 25506
rect 14978 25454 15150 25506
rect 15202 25454 15204 25506
rect 14924 25452 15204 25454
rect 14924 25442 14980 25452
rect 15148 25442 15204 25452
rect 14364 25394 14420 25406
rect 14364 25342 14366 25394
rect 14418 25342 14420 25394
rect 14364 25284 14420 25342
rect 15372 25396 15428 25406
rect 15372 25302 15428 25340
rect 15484 25394 15540 25406
rect 15484 25342 15486 25394
rect 15538 25342 15540 25394
rect 14364 25218 14420 25228
rect 14588 25282 14644 25294
rect 14588 25230 14590 25282
rect 14642 25230 14644 25282
rect 14588 24836 14644 25230
rect 14476 24780 14588 24836
rect 13916 24724 13972 24734
rect 13468 24722 13972 24724
rect 13468 24670 13470 24722
rect 13522 24670 13918 24722
rect 13970 24670 13972 24722
rect 13468 24668 13972 24670
rect 10556 24610 10612 24622
rect 12684 24612 12740 24622
rect 10556 24558 10558 24610
rect 10610 24558 10612 24610
rect 10556 24388 10612 24558
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 10556 24322 10612 24332
rect 12460 24610 12740 24612
rect 12460 24558 12686 24610
rect 12738 24558 12740 24610
rect 12460 24556 12740 24558
rect 4476 24266 4740 24276
rect 12460 24162 12516 24556
rect 12684 24546 12740 24556
rect 12460 24110 12462 24162
rect 12514 24110 12516 24162
rect 12460 24098 12516 24110
rect 12348 23940 12404 23950
rect 12348 23846 12404 23884
rect 13356 23156 13412 23166
rect 12796 23154 13412 23156
rect 12796 23102 13358 23154
rect 13410 23102 13412 23154
rect 12796 23100 13412 23102
rect 10668 23044 10724 23054
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 10668 22482 10724 22988
rect 10668 22430 10670 22482
rect 10722 22430 10724 22482
rect 10668 22418 10724 22430
rect 12796 22484 12852 23100
rect 13356 23090 13412 23100
rect 12796 22482 12964 22484
rect 12796 22430 12798 22482
rect 12850 22430 12964 22482
rect 12796 22428 12964 22430
rect 12796 22418 12852 22428
rect 4172 22082 4228 22092
rect 9996 22370 10052 22382
rect 9996 22318 9998 22370
rect 10050 22318 10052 22370
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 9996 20020 10052 22318
rect 12908 21810 12964 22428
rect 13468 21924 13524 24668
rect 13916 24658 13972 24668
rect 13804 24500 13860 24510
rect 13692 24444 13804 24500
rect 13692 23938 13748 24444
rect 13804 24434 13860 24444
rect 13916 24388 13972 24398
rect 13692 23886 13694 23938
rect 13746 23886 13748 23938
rect 13692 23874 13748 23886
rect 13804 24050 13860 24062
rect 13804 23998 13806 24050
rect 13858 23998 13860 24050
rect 13804 23940 13860 23998
rect 13804 23874 13860 23884
rect 13916 23938 13972 24332
rect 13916 23886 13918 23938
rect 13970 23886 13972 23938
rect 13916 23874 13972 23886
rect 14364 23828 14420 23838
rect 14364 23734 14420 23772
rect 14140 23714 14196 23726
rect 14140 23662 14142 23714
rect 14194 23662 14196 23714
rect 13692 23268 13748 23278
rect 13692 23266 14084 23268
rect 13692 23214 13694 23266
rect 13746 23214 14084 23266
rect 13692 23212 14084 23214
rect 13692 23202 13748 23212
rect 14028 22370 14084 23212
rect 14140 22596 14196 23662
rect 14140 22530 14196 22540
rect 14028 22318 14030 22370
rect 14082 22318 14084 22370
rect 13580 22146 13636 22158
rect 13580 22094 13582 22146
rect 13634 22094 13636 22146
rect 13580 21924 13636 22094
rect 12908 21758 12910 21810
rect 12962 21758 12964 21810
rect 12908 21746 12964 21758
rect 13356 21868 13636 21924
rect 9996 19926 10052 19964
rect 12684 20020 12740 20030
rect 10668 19908 10724 19918
rect 10668 19814 10724 19852
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 11676 18676 11732 18686
rect 4284 18452 4340 18462
rect 4284 18358 4340 18396
rect 9884 18452 9940 18462
rect 1932 18228 1988 18238
rect 1932 18134 1988 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1932 17780 1988 17790
rect 1932 17686 1988 17724
rect 9884 17778 9940 18396
rect 11676 18450 11732 18620
rect 12572 18676 12628 18686
rect 12572 18582 12628 18620
rect 11676 18398 11678 18450
rect 11730 18398 11732 18450
rect 11676 18386 11732 18398
rect 11788 18228 11844 18238
rect 11788 18226 12068 18228
rect 11788 18174 11790 18226
rect 11842 18174 12068 18226
rect 11788 18172 12068 18174
rect 11788 18162 11844 18172
rect 9884 17726 9886 17778
rect 9938 17726 9940 17778
rect 9884 17714 9940 17726
rect 12012 17778 12068 18172
rect 12012 17726 12014 17778
rect 12066 17726 12068 17778
rect 12012 17714 12068 17726
rect 4284 17668 4340 17678
rect 4284 17574 4340 17612
rect 12684 17668 12740 19964
rect 13244 20020 13300 20030
rect 13356 20020 13412 21868
rect 13300 19964 13412 20020
rect 13468 21474 13524 21486
rect 13468 21422 13470 21474
rect 13522 21422 13524 21474
rect 13244 19926 13300 19964
rect 12796 19906 12852 19918
rect 12796 19854 12798 19906
rect 12850 19854 12852 19906
rect 12796 19348 12852 19854
rect 13468 19796 13524 21422
rect 14028 21476 14084 22318
rect 14364 22260 14420 22270
rect 14476 22260 14532 24780
rect 14588 24770 14644 24780
rect 15484 24948 15540 25342
rect 15484 24500 15540 24892
rect 15932 25394 15988 25406
rect 15932 25342 15934 25394
rect 15986 25342 15988 25394
rect 15932 24612 15988 25342
rect 16044 24948 16100 24958
rect 16044 24854 16100 24892
rect 16156 24948 16212 24958
rect 16380 24948 16436 26126
rect 16828 26180 16884 28476
rect 17052 28532 17108 28542
rect 17052 28530 17444 28532
rect 17052 28478 17054 28530
rect 17106 28478 17444 28530
rect 17052 28476 17444 28478
rect 17052 28466 17108 28476
rect 17388 28082 17444 28476
rect 17388 28030 17390 28082
rect 17442 28030 17444 28082
rect 17388 28018 17444 28030
rect 17612 27972 17668 27982
rect 17500 27970 17668 27972
rect 17500 27918 17614 27970
rect 17666 27918 17668 27970
rect 17500 27916 17668 27918
rect 17388 27748 17444 27758
rect 16828 26178 16996 26180
rect 16828 26126 16830 26178
rect 16882 26126 16996 26178
rect 16828 26124 16996 26126
rect 16828 26114 16884 26124
rect 16156 24946 16436 24948
rect 16156 24894 16158 24946
rect 16210 24894 16436 24946
rect 16156 24892 16436 24894
rect 16156 24882 16212 24892
rect 16380 24724 16436 24734
rect 16156 24722 16436 24724
rect 16156 24670 16382 24722
rect 16434 24670 16436 24722
rect 16156 24668 16436 24670
rect 16044 24612 16100 24622
rect 15932 24610 16100 24612
rect 15932 24558 16046 24610
rect 16098 24558 16100 24610
rect 15932 24556 16100 24558
rect 16044 24546 16100 24556
rect 15484 24434 15540 24444
rect 16156 22932 16212 24668
rect 16380 24658 16436 24668
rect 16604 24724 16660 24734
rect 16156 22866 16212 22876
rect 16268 23828 16324 23838
rect 16268 23154 16324 23772
rect 16268 23102 16270 23154
rect 16322 23102 16324 23154
rect 14812 22596 14868 22606
rect 14364 22258 14756 22260
rect 14364 22206 14366 22258
rect 14418 22206 14756 22258
rect 14364 22204 14756 22206
rect 14364 22194 14420 22204
rect 14364 21586 14420 21598
rect 14364 21534 14366 21586
rect 14418 21534 14420 21586
rect 14140 21476 14196 21486
rect 14028 21474 14140 21476
rect 14028 21422 14030 21474
rect 14082 21422 14140 21474
rect 14028 21420 14140 21422
rect 14028 21410 14084 21420
rect 14140 20802 14196 21420
rect 14140 20750 14142 20802
rect 14194 20750 14196 20802
rect 14140 20738 14196 20750
rect 14364 20188 14420 21534
rect 14700 21476 14756 22204
rect 14812 21698 14868 22540
rect 16268 22484 16324 23102
rect 16492 23156 16548 23166
rect 16492 23062 16548 23100
rect 16380 23044 16436 23054
rect 16380 22950 16436 22988
rect 16268 22418 16324 22428
rect 15260 22258 15316 22270
rect 15260 22206 15262 22258
rect 15314 22206 15316 22258
rect 15260 21812 15316 22206
rect 15596 22148 15652 22158
rect 15596 22146 16548 22148
rect 15596 22094 15598 22146
rect 15650 22094 16548 22146
rect 15596 22092 16548 22094
rect 15596 22082 15652 22092
rect 15820 21924 15876 21934
rect 15260 21810 15764 21812
rect 15260 21758 15262 21810
rect 15314 21758 15764 21810
rect 15260 21756 15764 21758
rect 15260 21746 15316 21756
rect 14812 21646 14814 21698
rect 14866 21646 14868 21698
rect 14812 21634 14868 21646
rect 15708 21698 15764 21756
rect 15820 21810 15876 21868
rect 15820 21758 15822 21810
rect 15874 21758 15876 21810
rect 15820 21746 15876 21758
rect 15708 21646 15710 21698
rect 15762 21646 15764 21698
rect 15708 21634 15764 21646
rect 15932 21698 15988 21710
rect 15932 21646 15934 21698
rect 15986 21646 15988 21698
rect 15820 21588 15876 21598
rect 15148 21476 15204 21486
rect 14700 21420 14980 21476
rect 14700 20804 14756 20814
rect 14700 20802 14868 20804
rect 14700 20750 14702 20802
rect 14754 20750 14868 20802
rect 14700 20748 14868 20750
rect 14700 20738 14756 20748
rect 14700 20242 14756 20254
rect 14700 20190 14702 20242
rect 14754 20190 14756 20242
rect 14700 20188 14756 20190
rect 14140 20132 14196 20142
rect 14364 20132 14756 20188
rect 14140 20038 14196 20076
rect 13468 19730 13524 19740
rect 13692 20018 13748 20030
rect 13692 19966 13694 20018
rect 13746 19966 13748 20018
rect 12796 19282 12852 19292
rect 13132 19460 13188 19470
rect 13132 18450 13188 19404
rect 13692 19460 13748 19966
rect 13916 20018 13972 20030
rect 13916 19966 13918 20018
rect 13970 19966 13972 20018
rect 13916 19684 13972 19966
rect 14028 19908 14084 19918
rect 14028 19814 14084 19852
rect 14700 19908 14756 20132
rect 13916 19618 13972 19628
rect 13692 19394 13748 19404
rect 14028 19348 14084 19358
rect 14028 19254 14084 19292
rect 14476 19348 14532 19358
rect 14140 19236 14196 19246
rect 14140 19142 14196 19180
rect 14476 19234 14532 19292
rect 14476 19182 14478 19234
rect 14530 19182 14532 19234
rect 14476 19170 14532 19182
rect 14700 19124 14756 19852
rect 14812 19572 14868 20748
rect 14812 19506 14868 19516
rect 14812 19124 14868 19134
rect 14700 19122 14868 19124
rect 14700 19070 14814 19122
rect 14866 19070 14868 19122
rect 14700 19068 14868 19070
rect 14812 19058 14868 19068
rect 13468 19012 13524 19022
rect 13468 18674 13524 18956
rect 13468 18622 13470 18674
rect 13522 18622 13524 18674
rect 13468 18610 13524 18622
rect 13132 18398 13134 18450
rect 13186 18398 13188 18450
rect 13132 18386 13188 18398
rect 13692 18452 13748 18462
rect 12908 18340 12964 18350
rect 12908 18246 12964 18284
rect 13580 18340 13636 18350
rect 13580 18246 13636 18284
rect 13468 17668 13524 17678
rect 12684 17666 13076 17668
rect 12684 17614 12686 17666
rect 12738 17614 13076 17666
rect 12684 17612 13076 17614
rect 12684 17602 12740 17612
rect 13020 17108 13076 17612
rect 13468 17554 13524 17612
rect 13692 17666 13748 18396
rect 14140 18450 14196 18462
rect 14140 18398 14142 18450
rect 14194 18398 14196 18450
rect 14140 18340 14196 18398
rect 14140 18274 14196 18284
rect 14924 18340 14980 21420
rect 15148 21382 15204 21420
rect 15708 20692 15764 20702
rect 15596 20636 15708 20692
rect 15596 20244 15652 20636
rect 15708 20626 15764 20636
rect 14924 18274 14980 18284
rect 15036 20130 15092 20142
rect 15036 20078 15038 20130
rect 15090 20078 15092 20130
rect 15036 17892 15092 20078
rect 15484 20132 15540 20142
rect 15484 20018 15540 20076
rect 15484 19966 15486 20018
rect 15538 19966 15540 20018
rect 15484 19908 15540 19966
rect 15484 19842 15540 19852
rect 15372 19236 15428 19246
rect 15596 19236 15652 20188
rect 15820 20244 15876 21532
rect 15708 20132 15764 20142
rect 15820 20132 15876 20188
rect 15708 20130 15876 20132
rect 15708 20078 15710 20130
rect 15762 20078 15876 20130
rect 15708 20076 15876 20078
rect 15708 20066 15764 20076
rect 15708 19236 15764 19246
rect 15596 19234 15764 19236
rect 15596 19182 15710 19234
rect 15762 19182 15764 19234
rect 15596 19180 15764 19182
rect 15372 19142 15428 19180
rect 15708 19170 15764 19180
rect 15932 19236 15988 21646
rect 15932 19170 15988 19180
rect 16044 19572 16100 19582
rect 16044 19234 16100 19516
rect 16044 19182 16046 19234
rect 16098 19182 16100 19234
rect 16044 19170 16100 19182
rect 15036 17826 15092 17836
rect 15148 19012 15204 19022
rect 15148 17668 15204 18956
rect 15932 19012 15988 19022
rect 15932 18918 15988 18956
rect 13692 17614 13694 17666
rect 13746 17614 13748 17666
rect 13692 17602 13748 17614
rect 14700 17612 15204 17668
rect 13468 17502 13470 17554
rect 13522 17502 13524 17554
rect 13468 17490 13524 17502
rect 13020 17106 13412 17108
rect 13020 17054 13022 17106
rect 13074 17054 13412 17106
rect 13020 17052 13412 17054
rect 13020 17042 13076 17052
rect 4284 16884 4340 16894
rect 4284 16790 4340 16828
rect 11564 16884 11620 16894
rect 1932 16658 1988 16670
rect 1932 16606 1934 16658
rect 1986 16606 1988 16658
rect 1932 16212 1988 16606
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 1932 16146 1988 16156
rect 11564 15202 11620 16828
rect 13356 16772 13412 17052
rect 14700 17106 14756 17612
rect 15148 17554 15204 17612
rect 15260 17668 15316 17678
rect 16156 17668 16212 22092
rect 16492 21698 16548 22092
rect 16604 21810 16660 24668
rect 16940 23716 16996 26124
rect 17388 26178 17444 27692
rect 17500 26908 17556 27916
rect 17612 27906 17668 27916
rect 17724 27860 17780 27870
rect 17724 27766 17780 27804
rect 17836 27748 17892 37998
rect 19068 37490 19124 38612
rect 19516 38274 19572 41200
rect 19516 38222 19518 38274
rect 19570 38222 19572 38274
rect 19516 38210 19572 38222
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19068 37438 19070 37490
rect 19122 37438 19124 37490
rect 19068 37426 19124 37438
rect 20188 37492 20244 41200
rect 21532 38276 21588 41200
rect 21532 38210 21588 38220
rect 22428 38276 22484 38286
rect 22428 38182 22484 38220
rect 24220 38276 24276 41200
rect 25564 38500 25620 41200
rect 25564 38434 25620 38444
rect 24220 38210 24276 38220
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 21756 38050 21812 38062
rect 21756 37998 21758 38050
rect 21810 37998 21812 38050
rect 20188 37426 20244 37436
rect 21420 37492 21476 37502
rect 21420 37398 21476 37436
rect 19628 37268 19684 37278
rect 19180 37266 19684 37268
rect 19180 37214 19630 37266
rect 19682 37214 19684 37266
rect 19180 37212 19684 37214
rect 18956 29428 19012 29438
rect 18956 29334 19012 29372
rect 19180 28754 19236 37212
rect 19628 37202 19684 37212
rect 20636 37266 20692 37278
rect 20636 37214 20638 37266
rect 20690 37214 20692 37266
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19628 29316 19684 29326
rect 19180 28702 19182 28754
rect 19234 28702 19236 28754
rect 19068 28084 19124 28094
rect 19180 28084 19236 28702
rect 19516 29314 19684 29316
rect 19516 29262 19630 29314
rect 19682 29262 19684 29314
rect 19516 29260 19684 29262
rect 19516 28196 19572 29260
rect 19628 29250 19684 29260
rect 19628 28532 19684 28542
rect 19628 28438 19684 28476
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19516 28140 19684 28196
rect 19836 28186 20100 28196
rect 19068 28082 19236 28084
rect 19068 28030 19070 28082
rect 19122 28030 19236 28082
rect 19068 28028 19236 28030
rect 19628 28084 19684 28140
rect 19852 28084 19908 28094
rect 19628 28082 19908 28084
rect 19628 28030 19854 28082
rect 19906 28030 19908 28082
rect 19628 28028 19908 28030
rect 19068 28018 19124 28028
rect 19852 28018 19908 28028
rect 20076 27972 20132 27982
rect 19964 27970 20132 27972
rect 19964 27918 20078 27970
rect 20130 27918 20132 27970
rect 19964 27916 20132 27918
rect 18844 27860 18900 27870
rect 18844 27766 18900 27804
rect 19180 27860 19236 27870
rect 19180 27766 19236 27804
rect 17836 27682 17892 27692
rect 18956 27748 19012 27758
rect 18844 26962 18900 26974
rect 18844 26910 18846 26962
rect 18898 26910 18900 26962
rect 17500 26852 17668 26908
rect 17388 26126 17390 26178
rect 17442 26126 17444 26178
rect 17388 26114 17444 26126
rect 17388 25396 17444 25406
rect 17388 24722 17444 25340
rect 17388 24670 17390 24722
rect 17442 24670 17444 24722
rect 17276 23938 17332 23950
rect 17276 23886 17278 23938
rect 17330 23886 17332 23938
rect 17276 23716 17332 23886
rect 16940 23714 17332 23716
rect 16940 23662 16942 23714
rect 16994 23662 17332 23714
rect 16940 23660 17332 23662
rect 16828 23380 16884 23390
rect 16828 23154 16884 23324
rect 16828 23102 16830 23154
rect 16882 23102 16884 23154
rect 16828 23090 16884 23102
rect 16828 22260 16884 22270
rect 16604 21758 16606 21810
rect 16658 21758 16660 21810
rect 16604 21746 16660 21758
rect 16716 21924 16772 21934
rect 16492 21646 16494 21698
rect 16546 21646 16548 21698
rect 16492 21634 16548 21646
rect 16716 21476 16772 21868
rect 16828 21588 16884 22204
rect 16828 21522 16884 21532
rect 16604 21420 16772 21476
rect 16380 20244 16436 20254
rect 16436 20188 16548 20244
rect 16380 20178 16436 20188
rect 16268 20132 16324 20142
rect 16268 20018 16324 20076
rect 16268 19966 16270 20018
rect 16322 19966 16324 20018
rect 16268 19954 16324 19966
rect 16380 19460 16436 19470
rect 16380 19366 16436 19404
rect 16492 19122 16548 20188
rect 16604 19796 16660 21420
rect 16828 20692 16884 20702
rect 16940 20692 16996 23660
rect 17052 23156 17108 23166
rect 17052 22372 17108 23100
rect 17052 22316 17220 22372
rect 17052 22148 17108 22158
rect 17052 21588 17108 22092
rect 17052 21522 17108 21532
rect 16828 20690 16996 20692
rect 16828 20638 16830 20690
rect 16882 20638 16996 20690
rect 16828 20636 16996 20638
rect 16716 20132 16772 20142
rect 16716 20018 16772 20076
rect 16716 19966 16718 20018
rect 16770 19966 16772 20018
rect 16716 19954 16772 19966
rect 16828 20020 16884 20636
rect 16828 19954 16884 19964
rect 16716 19796 16772 19806
rect 16604 19794 16772 19796
rect 16604 19742 16718 19794
rect 16770 19742 16772 19794
rect 16604 19740 16772 19742
rect 16716 19730 16772 19740
rect 16716 19460 16772 19470
rect 16716 19366 16772 19404
rect 16492 19070 16494 19122
rect 16546 19070 16548 19122
rect 16492 19058 16548 19070
rect 17164 18900 17220 22316
rect 17388 22036 17444 24670
rect 17612 23380 17668 26852
rect 17724 24948 17780 24958
rect 17724 24854 17780 24892
rect 18844 24948 18900 26910
rect 18956 26962 19012 27692
rect 18956 26910 18958 26962
rect 19010 26910 19012 26962
rect 18956 26898 19012 26910
rect 19964 26908 20020 27916
rect 20076 27906 20132 27916
rect 20188 27860 20244 27870
rect 20524 27860 20580 27870
rect 20188 27858 20580 27860
rect 20188 27806 20190 27858
rect 20242 27806 20526 27858
rect 20578 27806 20580 27858
rect 20188 27804 20580 27806
rect 20188 27794 20244 27804
rect 20524 27794 20580 27804
rect 20636 26908 20692 37214
rect 21756 29316 21812 37998
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 20748 29314 21812 29316
rect 20748 29262 21758 29314
rect 21810 29262 21812 29314
rect 20748 29260 21812 29262
rect 20748 28082 20804 29260
rect 21756 29250 21812 29260
rect 21868 29428 21924 29438
rect 20748 28030 20750 28082
rect 20802 28030 20804 28082
rect 20748 28018 20804 28030
rect 20860 27860 20916 27870
rect 20860 27766 20916 27804
rect 21756 27860 21812 27870
rect 21868 27860 21924 29372
rect 22316 29428 22372 29438
rect 22316 29334 22372 29372
rect 21756 27858 21924 27860
rect 21756 27806 21758 27858
rect 21810 27806 21924 27858
rect 21756 27804 21924 27806
rect 23324 27860 23380 27870
rect 19180 26850 19236 26862
rect 19180 26798 19182 26850
rect 19234 26798 19236 26850
rect 19180 25506 19236 26798
rect 19628 26852 20020 26908
rect 20412 26852 20692 26908
rect 19516 26178 19572 26190
rect 19516 26126 19518 26178
rect 19570 26126 19572 26178
rect 19516 25618 19572 26126
rect 19516 25566 19518 25618
rect 19570 25566 19572 25618
rect 19516 25554 19572 25566
rect 19180 25454 19182 25506
rect 19234 25454 19236 25506
rect 19180 25442 19236 25454
rect 18844 24882 18900 24892
rect 19516 25282 19572 25294
rect 19516 25230 19518 25282
rect 19570 25230 19572 25282
rect 19516 24948 19572 25230
rect 19516 24882 19572 24892
rect 18060 23828 18116 23838
rect 18060 23826 18228 23828
rect 18060 23774 18062 23826
rect 18114 23774 18228 23826
rect 18060 23772 18228 23774
rect 18060 23762 18116 23772
rect 17500 22596 17556 22606
rect 17612 22596 17668 23324
rect 17836 23268 17892 23278
rect 17500 22594 17668 22596
rect 17500 22542 17502 22594
rect 17554 22542 17668 22594
rect 17500 22540 17668 22542
rect 17724 23212 17836 23268
rect 17500 22530 17556 22540
rect 17612 22372 17668 22382
rect 17724 22372 17780 23212
rect 17836 23202 17892 23212
rect 18172 23266 18228 23772
rect 19404 23380 19460 23390
rect 18172 23214 18174 23266
rect 18226 23214 18228 23266
rect 18172 23202 18228 23214
rect 18508 23378 19460 23380
rect 18508 23326 19406 23378
rect 19458 23326 19460 23378
rect 18508 23324 19460 23326
rect 18508 23154 18564 23324
rect 19404 23314 19460 23324
rect 19516 23380 19572 23390
rect 19516 23286 19572 23324
rect 19628 23380 19684 26852
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20300 26290 20356 26302
rect 20300 26238 20302 26290
rect 20354 26238 20356 26290
rect 20300 26180 20356 26238
rect 20300 26114 20356 26124
rect 19740 25508 19796 25518
rect 19740 25394 19796 25452
rect 19740 25342 19742 25394
rect 19794 25342 19796 25394
rect 19740 25330 19796 25342
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20188 24948 20244 24958
rect 20188 24854 20244 24892
rect 20076 24722 20132 24734
rect 20076 24670 20078 24722
rect 20130 24670 20132 24722
rect 20076 23716 20132 24670
rect 20300 24724 20356 24734
rect 20300 24630 20356 24668
rect 20188 24052 20244 24062
rect 20412 24052 20468 26852
rect 20748 26180 20804 26190
rect 20748 25284 20804 26124
rect 21644 25730 21700 25742
rect 21644 25678 21646 25730
rect 21698 25678 21700 25730
rect 21644 25508 21700 25678
rect 21644 25442 21700 25452
rect 20748 25218 20804 25228
rect 21532 25394 21588 25406
rect 21532 25342 21534 25394
rect 21586 25342 21588 25394
rect 21532 25060 21588 25342
rect 21532 24994 21588 25004
rect 21644 25282 21700 25294
rect 21644 25230 21646 25282
rect 21698 25230 21700 25282
rect 21644 24948 21700 25230
rect 21756 25284 21812 27804
rect 22428 27748 22484 27758
rect 23212 27748 23268 27758
rect 22428 27746 22596 27748
rect 22428 27694 22430 27746
rect 22482 27694 22596 27746
rect 22428 27692 22596 27694
rect 22428 27682 22484 27692
rect 22540 27298 22596 27692
rect 22540 27246 22542 27298
rect 22594 27246 22596 27298
rect 22540 27234 22596 27246
rect 22428 27074 22484 27086
rect 22428 27022 22430 27074
rect 22482 27022 22484 27074
rect 22428 26908 22484 27022
rect 21868 26852 22484 26908
rect 22540 26962 22596 26974
rect 22540 26910 22542 26962
rect 22594 26910 22596 26962
rect 22540 26908 22596 26910
rect 22988 26962 23044 26974
rect 22988 26910 22990 26962
rect 23042 26910 23044 26962
rect 22988 26908 23044 26910
rect 22540 26852 23044 26908
rect 23212 26962 23268 27692
rect 23212 26910 23214 26962
rect 23266 26910 23268 26962
rect 23212 26898 23268 26910
rect 23324 27074 23380 27804
rect 24556 27748 24612 37998
rect 26236 37940 26292 41200
rect 26908 38610 26964 41200
rect 26908 38558 26910 38610
rect 26962 38558 26964 38610
rect 26908 38546 26964 38558
rect 28364 38610 28420 38622
rect 28364 38558 28366 38610
rect 28418 38558 28420 38610
rect 26236 37874 26292 37884
rect 26796 38500 26852 38510
rect 26796 37490 26852 38444
rect 27468 37940 27524 37950
rect 27468 37846 27524 37884
rect 28364 37938 28420 38558
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 28364 37886 28366 37938
rect 28418 37886 28420 37938
rect 28364 37874 28420 37886
rect 26796 37438 26798 37490
rect 26850 37438 26852 37490
rect 26796 37426 26852 37438
rect 25788 37266 25844 37278
rect 25788 37214 25790 37266
rect 25842 37214 25844 37266
rect 24556 27654 24612 27692
rect 25340 27746 25396 27758
rect 25340 27694 25342 27746
rect 25394 27694 25396 27746
rect 23324 27022 23326 27074
rect 23378 27022 23380 27074
rect 21868 25508 21924 26852
rect 21868 25442 21924 25452
rect 22428 25676 23156 25732
rect 22092 25396 22148 25406
rect 22092 25302 22148 25340
rect 22428 25394 22484 25676
rect 23100 25620 23156 25676
rect 23324 25620 23380 27022
rect 25340 26628 25396 27694
rect 23100 25564 23380 25620
rect 25116 26572 25396 26628
rect 22428 25342 22430 25394
rect 22482 25342 22484 25394
rect 22428 25330 22484 25342
rect 22876 25506 22932 25518
rect 22876 25454 22878 25506
rect 22930 25454 22932 25506
rect 21756 25218 21812 25228
rect 22876 25284 22932 25454
rect 22876 25218 22932 25228
rect 21868 25172 21924 25182
rect 21868 25060 21924 25116
rect 21644 24882 21700 24892
rect 21756 25004 21924 25060
rect 22764 25060 22820 25070
rect 21756 24946 21812 25004
rect 21756 24894 21758 24946
rect 21810 24894 21812 24946
rect 20188 24050 20468 24052
rect 20188 23998 20190 24050
rect 20242 23998 20468 24050
rect 20188 23996 20468 23998
rect 20524 24834 20580 24846
rect 20524 24782 20526 24834
rect 20578 24782 20580 24834
rect 20188 23986 20244 23996
rect 20076 23660 20244 23716
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20188 23492 20244 23660
rect 20188 23426 20244 23436
rect 19964 23380 20020 23390
rect 19628 23378 20020 23380
rect 19628 23326 19630 23378
rect 19682 23326 19966 23378
rect 20018 23326 20020 23378
rect 19628 23324 20020 23326
rect 19628 23314 19684 23324
rect 19964 23314 20020 23324
rect 20300 23380 20356 23996
rect 20300 23314 20356 23324
rect 20188 23268 20244 23278
rect 20188 23174 20244 23212
rect 18508 23102 18510 23154
rect 18562 23102 18564 23154
rect 18508 23090 18564 23102
rect 19068 23156 19124 23166
rect 19068 23062 19124 23100
rect 19292 23154 19348 23166
rect 19292 23102 19294 23154
rect 19346 23102 19348 23154
rect 18284 22930 18340 22942
rect 18284 22878 18286 22930
rect 18338 22878 18340 22930
rect 17612 22370 17780 22372
rect 17612 22318 17614 22370
rect 17666 22318 17780 22370
rect 17612 22316 17780 22318
rect 17836 22484 17892 22494
rect 17388 21970 17444 21980
rect 17500 22146 17556 22158
rect 17500 22094 17502 22146
rect 17554 22094 17556 22146
rect 17500 21586 17556 22094
rect 17612 21924 17668 22316
rect 17612 21858 17668 21868
rect 17500 21534 17502 21586
rect 17554 21534 17556 21586
rect 17388 20018 17444 20030
rect 17388 19966 17390 20018
rect 17442 19966 17444 20018
rect 17388 19236 17444 19966
rect 17500 19460 17556 21534
rect 17724 21700 17780 21710
rect 17836 21700 17892 22428
rect 18284 22372 18340 22878
rect 18284 22306 18340 22316
rect 18620 22930 18676 22942
rect 18620 22878 18622 22930
rect 18674 22878 18676 22930
rect 18172 22258 18228 22270
rect 18172 22206 18174 22258
rect 18226 22206 18228 22258
rect 18172 21924 18228 22206
rect 18396 22260 18452 22270
rect 18284 22148 18340 22158
rect 18396 22148 18452 22204
rect 18284 22146 18452 22148
rect 18284 22094 18286 22146
rect 18338 22094 18452 22146
rect 18284 22092 18452 22094
rect 18508 22146 18564 22158
rect 18508 22094 18510 22146
rect 18562 22094 18564 22146
rect 18284 22082 18340 22092
rect 18172 21858 18228 21868
rect 18508 21812 18564 22094
rect 18620 21924 18676 22878
rect 19180 22596 19236 22606
rect 19180 22502 19236 22540
rect 19292 22594 19348 23102
rect 19292 22542 19294 22594
rect 19346 22542 19348 22594
rect 19292 22530 19348 22542
rect 20300 23154 20356 23166
rect 20300 23102 20302 23154
rect 20354 23102 20356 23154
rect 20300 22932 20356 23102
rect 18732 22370 18788 22382
rect 18732 22318 18734 22370
rect 18786 22318 18788 22370
rect 18732 22260 18788 22318
rect 18956 22372 19012 22382
rect 19628 22372 19684 22382
rect 18956 22370 19124 22372
rect 18956 22318 18958 22370
rect 19010 22318 19124 22370
rect 18956 22316 19124 22318
rect 18956 22306 19012 22316
rect 18732 22194 18788 22204
rect 18620 21858 18676 21868
rect 18956 21924 19012 21934
rect 18508 21746 18564 21756
rect 17724 21698 17892 21700
rect 17724 21646 17726 21698
rect 17778 21646 17892 21698
rect 17724 21644 17892 21646
rect 17724 19908 17780 21644
rect 18284 21588 18340 21598
rect 18284 21494 18340 21532
rect 18844 20244 18900 20254
rect 18844 20130 18900 20188
rect 18956 20242 19012 21868
rect 19068 20580 19124 22316
rect 19628 22278 19684 22316
rect 19740 22258 19796 22270
rect 19740 22206 19742 22258
rect 19794 22206 19796 22258
rect 19740 22148 19796 22206
rect 19068 20514 19124 20524
rect 19628 22092 19796 22148
rect 18956 20190 18958 20242
rect 19010 20190 19012 20242
rect 18956 20178 19012 20190
rect 18844 20078 18846 20130
rect 18898 20078 18900 20130
rect 18844 20066 18900 20078
rect 19068 20132 19124 20142
rect 19628 20132 19684 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20300 21924 20356 22876
rect 20524 22596 20580 24782
rect 21532 24836 21588 24846
rect 21532 24742 21588 24780
rect 21196 24722 21252 24734
rect 21196 24670 21198 24722
rect 21250 24670 21252 24722
rect 20300 21858 20356 21868
rect 20412 22258 20468 22270
rect 20412 22206 20414 22258
rect 20466 22206 20468 22258
rect 20300 21700 20356 21710
rect 20300 20802 20356 21644
rect 20300 20750 20302 20802
rect 20354 20750 20356 20802
rect 20300 20738 20356 20750
rect 20300 20580 20356 20590
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19964 20244 20020 20254
rect 19740 20132 19796 20142
rect 19628 20076 19740 20132
rect 17948 20020 18004 20030
rect 17948 19926 18004 19964
rect 18956 20020 19012 20030
rect 17724 19842 17780 19852
rect 17500 19394 17556 19404
rect 18620 19460 18676 19470
rect 18956 19460 19012 19964
rect 18620 19366 18676 19404
rect 18844 19404 19012 19460
rect 17388 19170 17444 19180
rect 16828 18844 17220 18900
rect 16492 17668 16548 17678
rect 15260 17666 16548 17668
rect 15260 17614 15262 17666
rect 15314 17614 16158 17666
rect 16210 17614 16494 17666
rect 16546 17614 16548 17666
rect 15260 17612 16548 17614
rect 15260 17602 15316 17612
rect 16156 17602 16212 17612
rect 16492 17602 16548 17612
rect 15148 17502 15150 17554
rect 15202 17502 15204 17554
rect 15148 17490 15204 17502
rect 16828 17556 16884 18844
rect 18844 18450 18900 19404
rect 18956 19234 19012 19246
rect 18956 19182 18958 19234
rect 19010 19182 19012 19234
rect 18956 18564 19012 19182
rect 19068 18676 19124 20076
rect 19740 20066 19796 20076
rect 19852 20020 19908 20030
rect 19628 19572 19684 19582
rect 19180 19460 19236 19470
rect 19180 19346 19236 19404
rect 19180 19294 19182 19346
rect 19234 19294 19236 19346
rect 19180 19282 19236 19294
rect 19628 19346 19684 19516
rect 19628 19294 19630 19346
rect 19682 19294 19684 19346
rect 19628 19282 19684 19294
rect 19852 19234 19908 19964
rect 19964 19906 20020 20188
rect 20076 20132 20132 20142
rect 20076 20018 20132 20076
rect 20076 19966 20078 20018
rect 20130 19966 20132 20018
rect 20076 19954 20132 19966
rect 19964 19854 19966 19906
rect 20018 19854 20020 19906
rect 19964 19842 20020 19854
rect 19852 19182 19854 19234
rect 19906 19182 19908 19234
rect 19852 19012 19908 19182
rect 20188 19236 20244 19246
rect 20300 19236 20356 20524
rect 20188 19234 20356 19236
rect 20188 19182 20190 19234
rect 20242 19182 20356 19234
rect 20188 19180 20356 19182
rect 20412 19460 20468 22206
rect 20188 19170 20244 19180
rect 19852 18956 20356 19012
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20188 18788 20244 18798
rect 19180 18676 19236 18686
rect 19068 18674 19236 18676
rect 19068 18622 19182 18674
rect 19234 18622 19236 18674
rect 19068 18620 19236 18622
rect 19180 18610 19236 18620
rect 19404 18676 19460 18686
rect 20188 18676 20244 18732
rect 19404 18582 19460 18620
rect 20076 18620 20244 18676
rect 18956 18498 19012 18508
rect 18844 18398 18846 18450
rect 18898 18398 18900 18450
rect 18844 18386 18900 18398
rect 17836 18228 17892 18238
rect 19068 18228 19124 18238
rect 17724 17668 17780 17678
rect 17836 17668 17892 18172
rect 18732 18226 19124 18228
rect 18732 18174 19070 18226
rect 19122 18174 19124 18226
rect 18732 18172 19124 18174
rect 17724 17666 17892 17668
rect 17724 17614 17726 17666
rect 17778 17614 17892 17666
rect 17724 17612 17892 17614
rect 18060 17668 18116 17678
rect 16828 17554 17444 17556
rect 16828 17502 16830 17554
rect 16882 17502 17444 17554
rect 16828 17500 17444 17502
rect 16828 17490 16884 17500
rect 14924 17444 14980 17454
rect 14924 17442 15092 17444
rect 14924 17390 14926 17442
rect 14978 17390 15092 17442
rect 14924 17388 15092 17390
rect 14924 17378 14980 17388
rect 14700 17054 14702 17106
rect 14754 17054 14756 17106
rect 14700 17042 14756 17054
rect 14924 16994 14980 17006
rect 14924 16942 14926 16994
rect 14978 16942 14980 16994
rect 14924 16884 14980 16942
rect 15036 16994 15092 17388
rect 15036 16942 15038 16994
rect 15090 16942 15092 16994
rect 15036 16930 15092 16942
rect 15820 17442 15876 17454
rect 15820 17390 15822 17442
rect 15874 17390 15876 17442
rect 14924 16818 14980 16828
rect 15484 16884 15540 16894
rect 15484 16790 15540 16828
rect 15820 16884 15876 17390
rect 16044 17444 16100 17454
rect 16044 17350 16100 17388
rect 16268 17332 16324 17342
rect 16156 17276 16268 17332
rect 15820 16882 15988 16884
rect 15820 16830 15822 16882
rect 15874 16830 15988 16882
rect 15820 16828 15988 16830
rect 15820 16818 15876 16828
rect 13356 16716 13524 16772
rect 11564 15150 11566 15202
rect 11618 15150 11620 15202
rect 11564 15138 11620 15150
rect 13020 15092 13076 15102
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 13020 13746 13076 15036
rect 13468 15092 13524 16716
rect 14812 16770 14868 16782
rect 14812 16718 14814 16770
rect 14866 16718 14868 16770
rect 14812 16098 14868 16718
rect 15820 16660 15876 16670
rect 15372 16658 15876 16660
rect 15372 16606 15822 16658
rect 15874 16606 15876 16658
rect 15372 16604 15876 16606
rect 14812 16046 14814 16098
rect 14866 16046 14868 16098
rect 14812 16034 14868 16046
rect 15036 16100 15092 16110
rect 15372 16100 15428 16604
rect 15820 16594 15876 16604
rect 15036 16006 15092 16044
rect 15148 16098 15428 16100
rect 15148 16046 15374 16098
rect 15426 16046 15428 16098
rect 15148 16044 15428 16046
rect 14924 15876 14980 15886
rect 13692 15874 14980 15876
rect 13692 15822 14926 15874
rect 14978 15822 14980 15874
rect 13692 15820 14980 15822
rect 13692 15426 13748 15820
rect 14924 15810 14980 15820
rect 13692 15374 13694 15426
rect 13746 15374 13748 15426
rect 13692 15362 13748 15374
rect 14364 15314 14420 15326
rect 14364 15262 14366 15314
rect 14418 15262 14420 15314
rect 13468 15026 13524 15036
rect 13804 15204 13860 15214
rect 13804 13858 13860 15148
rect 14364 15092 14420 15262
rect 15148 15314 15204 16044
rect 15372 16034 15428 16044
rect 15484 16100 15540 16110
rect 15484 15428 15540 16044
rect 15932 16100 15988 16828
rect 16156 16770 16212 17276
rect 16268 17266 16324 17276
rect 16156 16718 16158 16770
rect 16210 16718 16212 16770
rect 16156 16706 16212 16718
rect 15932 16034 15988 16044
rect 16156 16100 16212 16110
rect 15148 15262 15150 15314
rect 15202 15262 15204 15314
rect 15148 15250 15204 15262
rect 15372 15372 15540 15428
rect 16044 15426 16100 15438
rect 16044 15374 16046 15426
rect 16098 15374 16100 15426
rect 15372 15314 15428 15372
rect 15372 15262 15374 15314
rect 15426 15262 15428 15314
rect 15372 15250 15428 15262
rect 15596 15316 15652 15326
rect 15820 15316 15876 15326
rect 15596 15314 15876 15316
rect 15596 15262 15598 15314
rect 15650 15262 15822 15314
rect 15874 15262 15876 15314
rect 15596 15260 15876 15262
rect 15596 15250 15652 15260
rect 15820 15250 15876 15260
rect 15484 15204 15540 15242
rect 15484 15138 15540 15148
rect 14420 15036 14756 15092
rect 14364 15026 14420 15036
rect 14700 14644 14756 15036
rect 14700 14550 14756 14588
rect 15596 14644 15652 14654
rect 15596 14530 15652 14588
rect 15596 14478 15598 14530
rect 15650 14478 15652 14530
rect 15596 14466 15652 14478
rect 13804 13806 13806 13858
rect 13858 13806 13860 13858
rect 13804 13794 13860 13806
rect 13020 13694 13022 13746
rect 13074 13694 13076 13746
rect 13020 13682 13076 13694
rect 15932 13636 15988 13646
rect 16044 13636 16100 15374
rect 16156 15426 16212 16044
rect 16156 15374 16158 15426
rect 16210 15374 16212 15426
rect 16156 15362 16212 15374
rect 17388 15428 17444 17500
rect 17724 17444 17780 17612
rect 18060 17556 18116 17612
rect 17724 17378 17780 17388
rect 17836 17554 18116 17556
rect 17836 17502 18062 17554
rect 18114 17502 18116 17554
rect 17836 17500 18116 17502
rect 17612 16100 17668 16110
rect 17836 16100 17892 17500
rect 18060 17490 18116 17500
rect 17612 16098 17836 16100
rect 17612 16046 17614 16098
rect 17666 16046 17836 16098
rect 17612 16044 17836 16046
rect 17612 16034 17668 16044
rect 17836 16006 17892 16044
rect 18732 16884 18788 18172
rect 19068 18162 19124 18172
rect 20076 17666 20132 18620
rect 20300 18562 20356 18956
rect 20412 18788 20468 19404
rect 20412 18722 20468 18732
rect 20300 18510 20302 18562
rect 20354 18510 20356 18562
rect 20300 18498 20356 18510
rect 20412 18564 20468 18574
rect 20076 17614 20078 17666
rect 20130 17614 20132 17666
rect 19852 17444 19908 17482
rect 20076 17444 20132 17614
rect 20412 17666 20468 18508
rect 20412 17614 20414 17666
rect 20466 17614 20468 17666
rect 20412 17602 20468 17614
rect 20524 18452 20580 22540
rect 20860 23492 20916 23502
rect 20860 23154 20916 23436
rect 21196 23380 21252 24670
rect 21644 24612 21700 24622
rect 21644 24518 21700 24556
rect 20860 23102 20862 23154
rect 20914 23102 20916 23154
rect 20636 22146 20692 22158
rect 20636 22094 20638 22146
rect 20690 22094 20692 22146
rect 20636 21588 20692 22094
rect 20748 21588 20804 21598
rect 20636 21532 20748 21588
rect 20748 21522 20804 21532
rect 20636 19796 20692 19806
rect 20636 19702 20692 19740
rect 20860 19234 20916 23102
rect 21084 23324 21252 23380
rect 20972 23042 21028 23054
rect 20972 22990 20974 23042
rect 21026 22990 21028 23042
rect 20972 22148 21028 22990
rect 20972 22082 21028 22092
rect 20860 19182 20862 19234
rect 20914 19182 20916 19234
rect 20860 19170 20916 19182
rect 20972 21924 21028 21934
rect 20076 17388 20468 17444
rect 19852 17378 19908 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20412 17106 20468 17388
rect 20412 17054 20414 17106
rect 20466 17054 20468 17106
rect 20412 17042 20468 17054
rect 17388 15334 17444 15372
rect 17612 15876 17668 15886
rect 17612 15426 17668 15820
rect 17612 15374 17614 15426
rect 17666 15374 17668 15426
rect 17612 15362 17668 15374
rect 17724 15874 17780 15886
rect 17724 15822 17726 15874
rect 17778 15822 17780 15874
rect 16380 15204 16436 15214
rect 17724 15148 17780 15822
rect 17948 15874 18004 15886
rect 17948 15822 17950 15874
rect 18002 15822 18004 15874
rect 17948 15426 18004 15822
rect 17948 15374 17950 15426
rect 18002 15374 18004 15426
rect 17948 15362 18004 15374
rect 18060 15428 18116 15438
rect 18396 15428 18452 15438
rect 18116 15426 18452 15428
rect 18116 15374 18398 15426
rect 18450 15374 18452 15426
rect 18116 15372 18452 15374
rect 18060 15362 18116 15372
rect 18396 15362 18452 15372
rect 18732 15314 18788 16828
rect 20524 16212 20580 18396
rect 20860 18564 20916 18574
rect 20748 16882 20804 16894
rect 20748 16830 20750 16882
rect 20802 16830 20804 16882
rect 20748 16212 20804 16830
rect 20860 16884 20916 18508
rect 20972 18004 21028 21868
rect 21084 21588 21140 23324
rect 21756 23268 21812 24894
rect 22428 24948 22484 24958
rect 22428 24722 22484 24892
rect 22428 24670 22430 24722
rect 22482 24670 22484 24722
rect 22428 23940 22484 24670
rect 22764 24722 22820 25004
rect 22764 24670 22766 24722
rect 22818 24670 22820 24722
rect 22484 23884 22708 23940
rect 22428 23874 22484 23884
rect 21644 23212 21812 23268
rect 22540 23380 22596 23390
rect 21084 21522 21140 21532
rect 21196 23154 21252 23166
rect 21196 23102 21198 23154
rect 21250 23102 21252 23154
rect 21196 21028 21252 23102
rect 21308 23154 21364 23166
rect 21308 23102 21310 23154
rect 21362 23102 21364 23154
rect 21308 23044 21364 23102
rect 21308 22978 21364 22988
rect 21196 20972 21476 21028
rect 21308 20802 21364 20814
rect 21308 20750 21310 20802
rect 21362 20750 21364 20802
rect 21084 20132 21140 20142
rect 21084 20038 21140 20076
rect 21196 20018 21252 20030
rect 21196 19966 21198 20018
rect 21250 19966 21252 20018
rect 21196 18564 21252 19966
rect 21196 18450 21252 18508
rect 21196 18398 21198 18450
rect 21250 18398 21252 18450
rect 21196 18386 21252 18398
rect 21308 19458 21364 20750
rect 21308 19406 21310 19458
rect 21362 19406 21364 19458
rect 21308 18228 21364 19406
rect 21420 19234 21476 20972
rect 21644 20804 21700 23212
rect 21756 23044 21812 23054
rect 21756 22950 21812 22988
rect 21868 22370 21924 22382
rect 21868 22318 21870 22370
rect 21922 22318 21924 22370
rect 21756 21700 21812 21710
rect 21868 21700 21924 22318
rect 21812 21644 21924 21700
rect 21756 21606 21812 21644
rect 22540 20914 22596 23324
rect 22540 20862 22542 20914
rect 22594 20862 22596 20914
rect 22540 20850 22596 20862
rect 22652 20804 22708 23884
rect 22764 23604 22820 24670
rect 22988 24612 23044 24622
rect 23100 24612 23156 25564
rect 23660 25508 23716 25518
rect 23548 25396 23604 25406
rect 23324 25394 23604 25396
rect 23324 25342 23550 25394
rect 23602 25342 23604 25394
rect 23324 25340 23604 25342
rect 23324 24946 23380 25340
rect 23548 25330 23604 25340
rect 23660 25172 23716 25452
rect 23324 24894 23326 24946
rect 23378 24894 23380 24946
rect 23324 24882 23380 24894
rect 23436 25116 23716 25172
rect 23436 24834 23492 25116
rect 25116 24948 25172 26572
rect 25340 26404 25396 26414
rect 25788 26404 25844 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 25340 26402 25844 26404
rect 25340 26350 25342 26402
rect 25394 26350 25844 26402
rect 25340 26348 25844 26350
rect 25340 26338 25396 26348
rect 25228 26066 25284 26078
rect 25228 26014 25230 26066
rect 25282 26014 25284 26066
rect 25228 25508 25284 26014
rect 25676 25620 25732 25630
rect 25788 25620 25844 26348
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 25676 25618 25844 25620
rect 25676 25566 25678 25618
rect 25730 25566 25844 25618
rect 25676 25564 25844 25566
rect 40012 25618 40068 25630
rect 40012 25566 40014 25618
rect 40066 25566 40068 25618
rect 25676 25554 25732 25564
rect 25228 25442 25284 25452
rect 26236 25508 26292 25518
rect 26124 25396 26180 25406
rect 26124 25302 26180 25340
rect 26236 25394 26292 25452
rect 26236 25342 26238 25394
rect 26290 25342 26292 25394
rect 26236 25330 26292 25342
rect 28140 25508 28196 25518
rect 26460 25284 26516 25294
rect 26348 25282 26516 25284
rect 26348 25230 26462 25282
rect 26514 25230 26516 25282
rect 26348 25228 26516 25230
rect 25340 24948 25396 24958
rect 25116 24892 25340 24948
rect 23436 24782 23438 24834
rect 23490 24782 23492 24834
rect 23436 24770 23492 24782
rect 25340 24722 25396 24892
rect 25340 24670 25342 24722
rect 25394 24670 25396 24722
rect 23212 24612 23268 24622
rect 23100 24610 23268 24612
rect 23100 24558 23214 24610
rect 23266 24558 23268 24610
rect 23100 24556 23268 24558
rect 22988 24518 23044 24556
rect 23212 24546 23268 24556
rect 22764 23538 22820 23548
rect 23436 23604 23492 23614
rect 22876 21588 22932 21598
rect 21644 20748 22036 20804
rect 21644 20580 21700 20590
rect 21532 20524 21644 20580
rect 21532 19796 21588 20524
rect 21644 20486 21700 20524
rect 21756 20578 21812 20590
rect 21756 20526 21758 20578
rect 21810 20526 21812 20578
rect 21756 20132 21812 20526
rect 21868 20578 21924 20590
rect 21868 20526 21870 20578
rect 21922 20526 21924 20578
rect 21868 20244 21924 20526
rect 21868 20178 21924 20188
rect 21756 20066 21812 20076
rect 21980 19906 22036 20748
rect 22428 20692 22484 20702
rect 22428 20598 22484 20636
rect 22652 20690 22708 20748
rect 22652 20638 22654 20690
rect 22706 20638 22708 20690
rect 22652 20626 22708 20638
rect 22764 21364 22820 21374
rect 22764 20690 22820 21308
rect 22764 20638 22766 20690
rect 22818 20638 22820 20690
rect 22764 20356 22820 20638
rect 22428 20300 22820 20356
rect 21980 19854 21982 19906
rect 22034 19854 22036 19906
rect 21532 19740 21924 19796
rect 21868 19460 21924 19740
rect 21868 19366 21924 19404
rect 21420 19182 21422 19234
rect 21474 19182 21476 19234
rect 21420 18676 21476 19182
rect 21420 18610 21476 18620
rect 21980 18564 22036 19854
rect 22092 20018 22148 20030
rect 22092 19966 22094 20018
rect 22146 19966 22148 20018
rect 22092 19572 22148 19966
rect 22092 19458 22148 19516
rect 22092 19406 22094 19458
rect 22146 19406 22148 19458
rect 22092 19394 22148 19406
rect 22204 19012 22260 19022
rect 22428 19012 22484 20300
rect 22652 20132 22708 20142
rect 22652 20038 22708 20076
rect 22876 20018 22932 21532
rect 23436 21252 23492 23548
rect 24444 23268 24500 23278
rect 23884 23042 23940 23054
rect 23884 22990 23886 23042
rect 23938 22990 23940 23042
rect 23884 21698 23940 22990
rect 23884 21646 23886 21698
rect 23938 21646 23940 21698
rect 23884 21634 23940 21646
rect 24332 22148 24388 22158
rect 24332 21586 24388 22092
rect 24332 21534 24334 21586
rect 24386 21534 24388 21586
rect 24332 21522 24388 21534
rect 23996 21362 24052 21374
rect 23996 21310 23998 21362
rect 24050 21310 24052 21362
rect 23996 21252 24052 21310
rect 24220 21364 24276 21374
rect 24220 21270 24276 21308
rect 23436 21196 24052 21252
rect 23212 20802 23268 20814
rect 23212 20750 23214 20802
rect 23266 20750 23268 20802
rect 23212 20692 23268 20750
rect 23212 20626 23268 20636
rect 22876 19966 22878 20018
rect 22930 19966 22932 20018
rect 22876 19954 22932 19966
rect 23100 19908 23156 19918
rect 23100 19814 23156 19852
rect 23436 19796 23492 21196
rect 23884 20804 23940 20814
rect 23884 20690 23940 20748
rect 24444 20802 24500 23212
rect 24668 23156 24724 23166
rect 24668 23062 24724 23100
rect 25340 23156 25396 24670
rect 26012 24612 26068 24622
rect 25564 24610 26068 24612
rect 25564 24558 26014 24610
rect 26066 24558 26068 24610
rect 25564 24556 26068 24558
rect 25564 24050 25620 24556
rect 26012 24546 26068 24556
rect 25564 23998 25566 24050
rect 25618 23998 25620 24050
rect 25564 23986 25620 23998
rect 25676 23940 25732 23950
rect 25676 23846 25732 23884
rect 26124 23940 26180 23950
rect 26348 23940 26404 25228
rect 26460 25218 26516 25228
rect 26796 25282 26852 25294
rect 26796 25230 26798 25282
rect 26850 25230 26852 25282
rect 26796 24948 26852 25230
rect 26796 24882 26852 24892
rect 28140 24610 28196 25452
rect 37660 25508 37716 25518
rect 37660 25414 37716 25452
rect 28588 24948 28644 24958
rect 28588 24854 28644 24892
rect 40012 24948 40068 25566
rect 40012 24882 40068 24892
rect 28140 24558 28142 24610
rect 28194 24558 28196 24610
rect 28140 24546 28196 24558
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 26124 23938 26404 23940
rect 26124 23886 26126 23938
rect 26178 23886 26404 23938
rect 26124 23884 26404 23886
rect 26124 23874 26180 23884
rect 25340 23042 25396 23100
rect 25340 22990 25342 23042
rect 25394 22990 25396 23042
rect 24444 20750 24446 20802
rect 24498 20750 24500 20802
rect 24444 20738 24500 20750
rect 25004 21812 25060 21822
rect 25004 20802 25060 21756
rect 25340 21474 25396 22990
rect 25340 21422 25342 21474
rect 25394 21422 25396 21474
rect 25340 21362 25396 21422
rect 25340 21310 25342 21362
rect 25394 21310 25396 21362
rect 25340 21298 25396 21310
rect 25452 23714 25508 23726
rect 25452 23662 25454 23714
rect 25506 23662 25508 23714
rect 25452 23492 25508 23662
rect 25452 21924 25508 23436
rect 26796 23492 26852 23502
rect 26684 23380 26740 23390
rect 26572 23268 26628 23278
rect 26572 23174 26628 23212
rect 26684 23266 26740 23324
rect 26684 23214 26686 23266
rect 26738 23214 26740 23266
rect 26684 23202 26740 23214
rect 26796 23266 26852 23436
rect 26796 23214 26798 23266
rect 26850 23214 26852 23266
rect 26796 23202 26852 23214
rect 28140 23268 28196 23278
rect 26348 23154 26404 23166
rect 26348 23102 26350 23154
rect 26402 23102 26404 23154
rect 25004 20750 25006 20802
rect 25058 20750 25060 20802
rect 23884 20638 23886 20690
rect 23938 20638 23940 20690
rect 23884 20626 23940 20638
rect 24108 20692 24164 20702
rect 24108 20598 24164 20636
rect 23436 19730 23492 19740
rect 23548 20578 23604 20590
rect 23548 20526 23550 20578
rect 23602 20526 23604 20578
rect 22652 19460 22708 19470
rect 22204 19010 22484 19012
rect 22204 18958 22206 19010
rect 22258 18958 22484 19010
rect 22204 18956 22484 18958
rect 22540 19010 22596 19022
rect 22540 18958 22542 19010
rect 22594 18958 22596 19010
rect 22204 18946 22260 18956
rect 22540 18788 22596 18958
rect 22540 18722 22596 18732
rect 22652 18674 22708 19404
rect 22652 18622 22654 18674
rect 22706 18622 22708 18674
rect 22652 18610 22708 18622
rect 22876 19010 22932 19022
rect 22876 18958 22878 19010
rect 22930 18958 22932 19010
rect 22876 18676 22932 18958
rect 22876 18610 22932 18620
rect 23548 18676 23604 20526
rect 24332 20578 24388 20590
rect 24332 20526 24334 20578
rect 24386 20526 24388 20578
rect 24220 20132 24276 20142
rect 24220 20038 24276 20076
rect 23548 18610 23604 18620
rect 22204 18564 22260 18574
rect 21644 18562 22260 18564
rect 21644 18510 22206 18562
rect 22258 18510 22260 18562
rect 21644 18508 22260 18510
rect 21420 18452 21476 18462
rect 21420 18358 21476 18396
rect 21308 18162 21364 18172
rect 21532 18340 21588 18350
rect 20972 17948 21364 18004
rect 20972 17444 21028 17948
rect 21308 17666 21364 17948
rect 21308 17614 21310 17666
rect 21362 17614 21364 17666
rect 21308 17602 21364 17614
rect 21532 17666 21588 18284
rect 21532 17614 21534 17666
rect 21586 17614 21588 17666
rect 21532 17602 21588 17614
rect 20972 17378 21028 17388
rect 21644 17332 21700 18508
rect 22204 18498 22260 18508
rect 22988 18450 23044 18462
rect 22988 18398 22990 18450
rect 23042 18398 23044 18450
rect 21868 17892 21924 17930
rect 21868 17826 21924 17836
rect 21868 17668 21924 17678
rect 21868 17574 21924 17612
rect 21756 17444 21812 17454
rect 21756 17350 21812 17388
rect 21532 17276 21700 17332
rect 21084 16884 21140 16894
rect 20860 16882 21140 16884
rect 20860 16830 21086 16882
rect 21138 16830 21140 16882
rect 20860 16828 21140 16830
rect 21084 16818 21140 16828
rect 20524 16210 20692 16212
rect 20524 16158 20526 16210
rect 20578 16158 20692 16210
rect 20524 16156 20692 16158
rect 20524 16146 20580 16156
rect 19180 16100 19236 16110
rect 18732 15262 18734 15314
rect 18786 15262 18788 15314
rect 18732 15250 18788 15262
rect 19068 15314 19124 15326
rect 19068 15262 19070 15314
rect 19122 15262 19124 15314
rect 16268 14644 16324 14654
rect 16268 13972 16324 14588
rect 16380 14642 16436 15148
rect 16380 14590 16382 14642
rect 16434 14590 16436 14642
rect 16380 14578 16436 14590
rect 17612 15092 17780 15148
rect 17836 15204 17892 15242
rect 18844 15202 18900 15214
rect 18844 15150 18846 15202
rect 18898 15150 18900 15202
rect 18844 15148 18900 15150
rect 17836 15138 17892 15148
rect 18284 15092 18900 15148
rect 17612 14644 17668 15092
rect 16380 13972 16436 13982
rect 16828 13972 16884 13982
rect 16268 13970 16884 13972
rect 16268 13918 16382 13970
rect 16434 13918 16830 13970
rect 16882 13918 16884 13970
rect 16268 13916 16884 13918
rect 16380 13906 16436 13916
rect 16828 13748 16884 13916
rect 16828 13682 16884 13692
rect 17500 13748 17556 13758
rect 17500 13654 17556 13692
rect 15932 13634 16100 13636
rect 15932 13582 15934 13634
rect 15986 13582 16100 13634
rect 15932 13580 16100 13582
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 15932 8428 15988 13580
rect 15932 8372 16436 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 16156 5236 16212 5246
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 16156 800 16212 5180
rect 16380 5122 16436 8372
rect 17388 5236 17444 5246
rect 17388 5142 17444 5180
rect 16380 5070 16382 5122
rect 16434 5070 16436 5122
rect 16380 5058 16436 5070
rect 17612 4338 17668 14588
rect 18284 13858 18340 15092
rect 19068 14754 19124 15262
rect 19068 14702 19070 14754
rect 19122 14702 19124 14754
rect 19068 14690 19124 14702
rect 18508 14644 18564 14654
rect 18508 14550 18564 14588
rect 19180 14530 19236 16044
rect 20636 15988 20692 16156
rect 20748 16118 20804 16156
rect 20636 15932 21028 15988
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20972 15426 21028 15932
rect 21532 15876 21588 17276
rect 21644 17108 21700 17118
rect 22988 17108 23044 18398
rect 21700 17052 21924 17108
rect 21644 17014 21700 17052
rect 21868 16210 21924 17052
rect 21868 16158 21870 16210
rect 21922 16158 21924 16210
rect 21868 16146 21924 16158
rect 22764 16882 22820 16894
rect 22764 16830 22766 16882
rect 22818 16830 22820 16882
rect 22764 16212 22820 16830
rect 22988 16882 23044 17052
rect 22988 16830 22990 16882
rect 23042 16830 23044 16882
rect 22988 16818 23044 16830
rect 24332 17892 24388 20526
rect 25004 20244 25060 20750
rect 25340 20692 25396 20702
rect 25452 20692 25508 21868
rect 26236 22258 26292 22270
rect 26236 22206 26238 22258
rect 26290 22206 26292 22258
rect 26236 21586 26292 22206
rect 26236 21534 26238 21586
rect 26290 21534 26292 21586
rect 25900 21476 25956 21486
rect 26236 21476 26292 21534
rect 25900 21474 26292 21476
rect 25900 21422 25902 21474
rect 25954 21422 26292 21474
rect 25900 21420 26292 21422
rect 25900 21362 25956 21420
rect 25900 21310 25902 21362
rect 25954 21310 25956 21362
rect 25340 20690 25508 20692
rect 25340 20638 25342 20690
rect 25394 20638 25508 20690
rect 25340 20636 25508 20638
rect 25788 20804 25844 20814
rect 25900 20804 25956 21310
rect 25788 20802 25956 20804
rect 25788 20750 25790 20802
rect 25842 20750 25956 20802
rect 25788 20748 25956 20750
rect 25340 20626 25396 20636
rect 25004 20178 25060 20188
rect 24556 20132 24612 20142
rect 24556 20038 24612 20076
rect 25564 20020 25620 20030
rect 25564 19926 25620 19964
rect 25676 19908 25732 19918
rect 25676 19814 25732 19852
rect 25788 18450 25844 20748
rect 26348 20468 26404 23102
rect 26684 23042 26740 23054
rect 26684 22990 26686 23042
rect 26738 22990 26740 23042
rect 26572 21924 26628 21934
rect 26236 20412 26404 20468
rect 26460 20690 26516 20702
rect 26460 20638 26462 20690
rect 26514 20638 26516 20690
rect 25900 20244 25956 20254
rect 25900 20130 25956 20188
rect 25900 20078 25902 20130
rect 25954 20078 25956 20130
rect 25900 20066 25956 20078
rect 26124 20132 26180 20142
rect 26236 20132 26292 20412
rect 26348 20244 26404 20254
rect 26460 20244 26516 20638
rect 26348 20242 26516 20244
rect 26348 20190 26350 20242
rect 26402 20190 26516 20242
rect 26348 20188 26516 20190
rect 26348 20178 26404 20188
rect 26180 20130 26292 20132
rect 26180 20078 26238 20130
rect 26290 20078 26292 20130
rect 26180 20076 26292 20078
rect 26124 19234 26180 20076
rect 26236 20066 26292 20076
rect 26460 20020 26516 20030
rect 26460 19926 26516 19964
rect 26124 19182 26126 19234
rect 26178 19182 26180 19234
rect 26124 18564 26180 19182
rect 26348 19908 26404 19918
rect 26348 19236 26404 19852
rect 26348 19180 26516 19236
rect 26460 19122 26516 19180
rect 26460 19070 26462 19122
rect 26514 19070 26516 19122
rect 26460 19058 26516 19070
rect 26572 19124 26628 21868
rect 26684 21812 26740 22990
rect 28140 22594 28196 23212
rect 37660 23044 37716 23054
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 28140 22542 28142 22594
rect 28194 22542 28196 22594
rect 28140 22530 28196 22542
rect 37660 22370 37716 22988
rect 37660 22318 37662 22370
rect 37714 22318 37716 22370
rect 37660 22306 37716 22318
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 28252 22258 28308 22270
rect 28252 22206 28254 22258
rect 28306 22206 28308 22258
rect 26684 21756 27076 21812
rect 27020 21698 27076 21756
rect 27020 21646 27022 21698
rect 27074 21646 27076 21698
rect 27020 21634 27076 21646
rect 28252 21476 28308 22206
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 37660 21588 37716 21598
rect 37660 21494 37716 21532
rect 40012 21588 40068 21598
rect 28252 21410 28308 21420
rect 29148 21476 29204 21486
rect 29148 21382 29204 21420
rect 40012 21474 40068 21532
rect 40012 21422 40014 21474
rect 40066 21422 40068 21474
rect 40012 21410 40068 21422
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 27916 20916 27972 20926
rect 27916 20130 27972 20860
rect 28588 20916 28644 20926
rect 28588 20822 28644 20860
rect 40012 20916 40068 20926
rect 40012 20822 40068 20860
rect 37660 20804 37716 20814
rect 37660 20710 37716 20748
rect 27916 20078 27918 20130
rect 27970 20078 27972 20130
rect 27916 20066 27972 20078
rect 27804 20020 27860 20030
rect 27804 19926 27860 19964
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 26572 19122 26852 19124
rect 26572 19070 26574 19122
rect 26626 19070 26852 19122
rect 26572 19068 26852 19070
rect 26572 19058 26628 19068
rect 26236 19010 26292 19022
rect 26236 18958 26238 19010
rect 26290 18958 26292 19010
rect 26236 18676 26292 18958
rect 26348 19010 26404 19022
rect 26348 18958 26350 19010
rect 26402 18958 26404 19010
rect 26348 18788 26404 18958
rect 26348 18732 26740 18788
rect 26236 18620 26628 18676
rect 26124 18508 26516 18564
rect 25788 18398 25790 18450
rect 25842 18398 25844 18450
rect 24668 18340 24724 18350
rect 24780 18340 24836 18350
rect 24668 18338 24780 18340
rect 24668 18286 24670 18338
rect 24722 18286 24780 18338
rect 24668 18284 24780 18286
rect 24668 18274 24724 18284
rect 23212 16772 23268 16782
rect 23212 16770 23492 16772
rect 23212 16718 23214 16770
rect 23266 16718 23492 16770
rect 23212 16716 23492 16718
rect 23212 16706 23268 16716
rect 21532 15810 21588 15820
rect 20972 15374 20974 15426
rect 21026 15374 21028 15426
rect 20972 15362 21028 15374
rect 20300 15316 20356 15326
rect 20300 15222 20356 15260
rect 22764 15204 22820 16156
rect 23436 15426 23492 16716
rect 23996 16212 24052 16222
rect 24332 16212 24388 17836
rect 23772 16210 24388 16212
rect 23772 16158 23998 16210
rect 24050 16158 24388 16210
rect 23772 16156 24388 16158
rect 23772 15538 23828 16156
rect 23996 16146 24052 16156
rect 23772 15486 23774 15538
rect 23826 15486 23828 15538
rect 23772 15474 23828 15486
rect 24780 16100 24836 18284
rect 25228 18338 25284 18350
rect 25228 18286 25230 18338
rect 25282 18286 25284 18338
rect 25228 17444 25284 18286
rect 25788 18340 25844 18398
rect 25788 18274 25844 18284
rect 25340 18228 25396 18238
rect 25340 18226 25732 18228
rect 25340 18174 25342 18226
rect 25394 18174 25732 18226
rect 25340 18172 25732 18174
rect 25340 18162 25396 18172
rect 25676 17666 25732 18172
rect 26124 17780 26180 17790
rect 25676 17614 25678 17666
rect 25730 17614 25732 17666
rect 25676 17602 25732 17614
rect 26012 17778 26180 17780
rect 26012 17726 26126 17778
rect 26178 17726 26180 17778
rect 26012 17724 26180 17726
rect 25228 17378 25284 17388
rect 26012 16994 26068 17724
rect 26124 17714 26180 17724
rect 26460 17666 26516 18508
rect 26572 18562 26628 18620
rect 26572 18510 26574 18562
rect 26626 18510 26628 18562
rect 26572 18498 26628 18510
rect 26684 17892 26740 18732
rect 26684 17826 26740 17836
rect 26460 17614 26462 17666
rect 26514 17614 26516 17666
rect 26460 17602 26516 17614
rect 26124 17556 26180 17566
rect 26124 17462 26180 17500
rect 26236 17554 26292 17566
rect 26236 17502 26238 17554
rect 26290 17502 26292 17554
rect 26236 17444 26292 17502
rect 26796 17556 26852 19068
rect 37660 18452 37716 18462
rect 37660 18358 37716 18396
rect 27804 18340 27860 18350
rect 27692 17892 27748 17902
rect 27692 17798 27748 17836
rect 27804 17778 27860 18284
rect 28700 18340 28756 18350
rect 28700 18246 28756 18284
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 27804 17726 27806 17778
rect 27858 17726 27860 17778
rect 27804 17714 27860 17726
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 27132 17668 27188 17678
rect 27132 17574 27188 17612
rect 28140 17668 28196 17678
rect 26796 17490 26852 17500
rect 26236 17378 26292 17388
rect 27020 17444 27076 17454
rect 27020 17350 27076 17388
rect 26012 16942 26014 16994
rect 26066 16942 26068 16994
rect 26012 16930 26068 16942
rect 25228 16884 25284 16894
rect 25228 16100 25284 16828
rect 28140 16770 28196 17612
rect 37660 17668 37716 17678
rect 37660 17574 37716 17612
rect 28588 16884 28644 16894
rect 28588 16790 28644 16828
rect 40012 16884 40068 17726
rect 40012 16818 40068 16828
rect 28140 16718 28142 16770
rect 28194 16718 28196 16770
rect 28140 16706 28196 16718
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 24780 16098 25284 16100
rect 24780 16046 24782 16098
rect 24834 16046 25230 16098
rect 25282 16046 25284 16098
rect 24780 16044 25284 16046
rect 23436 15374 23438 15426
rect 23490 15374 23492 15426
rect 23436 15362 23492 15374
rect 24220 15316 24276 15326
rect 24220 15222 24276 15260
rect 24780 15316 24836 16044
rect 25228 16034 25284 16044
rect 24780 15250 24836 15260
rect 23100 15204 23156 15214
rect 22764 15202 23156 15204
rect 22764 15150 23102 15202
rect 23154 15150 23156 15202
rect 22764 15148 23156 15150
rect 23100 15138 23156 15148
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 19180 14478 19182 14530
rect 19234 14478 19236 14530
rect 19180 14466 19236 14478
rect 19068 14308 19124 14318
rect 19068 14214 19124 14252
rect 19628 14306 19684 14318
rect 19628 14254 19630 14306
rect 19682 14254 19684 14306
rect 18284 13806 18286 13858
rect 18338 13806 18340 13858
rect 18284 13794 18340 13806
rect 19628 13748 19684 14254
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20748 13860 20804 13870
rect 20524 13858 20804 13860
rect 20524 13806 20750 13858
rect 20802 13806 20804 13858
rect 20524 13804 20804 13806
rect 19628 13682 19684 13692
rect 19852 13748 19908 13758
rect 19852 12740 19908 13692
rect 20412 13748 20468 13758
rect 20412 13634 20468 13692
rect 20412 13582 20414 13634
rect 20466 13582 20468 13634
rect 20412 13570 20468 13582
rect 17612 4286 17614 4338
rect 17666 4286 17668 4338
rect 17612 4274 17668 4286
rect 19628 12738 19908 12740
rect 19628 12686 19854 12738
rect 19906 12686 19908 12738
rect 19628 12684 19908 12686
rect 18508 4116 18564 4126
rect 18172 4114 18564 4116
rect 18172 4062 18510 4114
rect 18562 4062 18564 4114
rect 18172 4060 18564 4062
rect 18172 800 18228 4060
rect 18508 4050 18564 4060
rect 19628 3556 19684 12684
rect 19852 12674 19908 12684
rect 20188 12740 20244 12750
rect 20188 12646 20244 12684
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20524 8428 20580 13804
rect 20748 13794 20804 13804
rect 20972 13748 21028 13758
rect 20972 13654 21028 13692
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 20860 12740 20916 12750
rect 20916 12684 21140 12740
rect 20860 12674 20916 12684
rect 20412 8372 20580 8428
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 20412 4338 20468 8372
rect 20412 4286 20414 4338
rect 20466 4286 20468 4338
rect 20412 4274 20468 4286
rect 20188 4116 20244 4126
rect 19740 3556 19796 3566
rect 19628 3554 19796 3556
rect 19628 3502 19742 3554
rect 19794 3502 19796 3554
rect 19628 3500 19796 3502
rect 19740 3490 19796 3500
rect 19180 3332 19236 3342
rect 19180 3330 19572 3332
rect 19180 3278 19182 3330
rect 19234 3278 19572 3330
rect 19180 3276 19572 3278
rect 19180 3266 19236 3276
rect 19516 800 19572 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 800 20244 4060
rect 20860 3668 20916 3678
rect 20860 800 20916 3612
rect 21084 3554 21140 12684
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 40236 11170 40292 11182
rect 40236 11118 40238 11170
rect 40290 11118 40292 11170
rect 40236 10836 40292 11118
rect 40236 10770 40292 10780
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 21420 4116 21476 4126
rect 21420 4022 21476 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 22092 3668 22148 3678
rect 22092 3574 22148 3612
rect 21084 3502 21086 3554
rect 21138 3502 21140 3554
rect 21084 3490 21140 3502
rect 16128 0 16240 800
rect 18144 0 18256 800
rect 19488 0 19600 800
rect 20160 0 20272 800
rect 20832 0 20944 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 16156 36652 16212 36708
rect 17388 36706 17444 36708
rect 17388 36654 17390 36706
rect 17390 36654 17442 36706
rect 17442 36654 17444 36706
rect 17388 36652 17444 36654
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 16380 28476 16436 28532
rect 4172 28252 4228 28308
rect 1932 25564 1988 25620
rect 1932 24498 1988 24500
rect 1932 24446 1934 24498
rect 1934 24446 1986 24498
rect 1986 24446 1988 24498
rect 1932 24444 1988 24446
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4284 26290 4340 26292
rect 4284 26238 4286 26290
rect 4286 26238 4338 26290
rect 4338 26238 4340 26290
rect 4284 26236 4340 26238
rect 12012 26236 12068 26292
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 12012 25340 12068 25396
rect 13580 26908 13636 26964
rect 4284 24722 4340 24724
rect 4284 24670 4286 24722
rect 4286 24670 4338 24722
rect 4338 24670 4340 24722
rect 4284 24668 4340 24670
rect 14252 26178 14308 26180
rect 14252 26126 14254 26178
rect 14254 26126 14306 26178
rect 14306 26126 14308 26178
rect 14252 26124 14308 26126
rect 14812 26908 14868 26964
rect 16828 28476 16884 28532
rect 15820 26124 15876 26180
rect 15372 25394 15428 25396
rect 15372 25342 15374 25394
rect 15374 25342 15426 25394
rect 15426 25342 15428 25394
rect 15372 25340 15428 25342
rect 14364 25228 14420 25284
rect 14588 24780 14644 24836
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 10556 24332 10612 24388
rect 4684 24276 4740 24278
rect 12348 23938 12404 23940
rect 12348 23886 12350 23938
rect 12350 23886 12402 23938
rect 12402 23886 12404 23938
rect 12348 23884 12404 23886
rect 10668 22988 10724 23044
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4172 22092 4228 22148
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 13804 24444 13860 24500
rect 13916 24332 13972 24388
rect 13804 23884 13860 23940
rect 14364 23826 14420 23828
rect 14364 23774 14366 23826
rect 14366 23774 14418 23826
rect 14418 23774 14420 23826
rect 14364 23772 14420 23774
rect 14140 22540 14196 22596
rect 9996 20018 10052 20020
rect 9996 19966 9998 20018
rect 9998 19966 10050 20018
rect 10050 19966 10052 20018
rect 9996 19964 10052 19966
rect 12684 19964 12740 20020
rect 10668 19906 10724 19908
rect 10668 19854 10670 19906
rect 10670 19854 10722 19906
rect 10722 19854 10724 19906
rect 10668 19852 10724 19854
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 11676 18620 11732 18676
rect 4284 18450 4340 18452
rect 4284 18398 4286 18450
rect 4286 18398 4338 18450
rect 4338 18398 4340 18450
rect 4284 18396 4340 18398
rect 9884 18396 9940 18452
rect 1932 18226 1988 18228
rect 1932 18174 1934 18226
rect 1934 18174 1986 18226
rect 1986 18174 1988 18226
rect 1932 18172 1988 18174
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 1932 17778 1988 17780
rect 1932 17726 1934 17778
rect 1934 17726 1986 17778
rect 1986 17726 1988 17778
rect 1932 17724 1988 17726
rect 12572 18674 12628 18676
rect 12572 18622 12574 18674
rect 12574 18622 12626 18674
rect 12626 18622 12628 18674
rect 12572 18620 12628 18622
rect 4284 17666 4340 17668
rect 4284 17614 4286 17666
rect 4286 17614 4338 17666
rect 4338 17614 4340 17666
rect 4284 17612 4340 17614
rect 13244 20018 13300 20020
rect 13244 19966 13246 20018
rect 13246 19966 13298 20018
rect 13298 19966 13300 20018
rect 13244 19964 13300 19966
rect 15484 24892 15540 24948
rect 16044 24946 16100 24948
rect 16044 24894 16046 24946
rect 16046 24894 16098 24946
rect 16098 24894 16100 24946
rect 16044 24892 16100 24894
rect 17388 27692 17444 27748
rect 15484 24444 15540 24500
rect 16604 24722 16660 24724
rect 16604 24670 16606 24722
rect 16606 24670 16658 24722
rect 16658 24670 16660 24722
rect 16604 24668 16660 24670
rect 16156 22876 16212 22932
rect 16268 23772 16324 23828
rect 14812 22540 14868 22596
rect 14140 21420 14196 21476
rect 16492 23154 16548 23156
rect 16492 23102 16494 23154
rect 16494 23102 16546 23154
rect 16546 23102 16548 23154
rect 16492 23100 16548 23102
rect 16380 23042 16436 23044
rect 16380 22990 16382 23042
rect 16382 22990 16434 23042
rect 16434 22990 16436 23042
rect 16380 22988 16436 22990
rect 16268 22428 16324 22484
rect 15820 21868 15876 21924
rect 15820 21532 15876 21588
rect 14140 20130 14196 20132
rect 14140 20078 14142 20130
rect 14142 20078 14194 20130
rect 14194 20078 14196 20130
rect 14140 20076 14196 20078
rect 13468 19740 13524 19796
rect 12796 19292 12852 19348
rect 13132 19404 13188 19460
rect 14028 19906 14084 19908
rect 14028 19854 14030 19906
rect 14030 19854 14082 19906
rect 14082 19854 14084 19906
rect 14028 19852 14084 19854
rect 14700 19852 14756 19908
rect 13916 19628 13972 19684
rect 13692 19404 13748 19460
rect 14028 19346 14084 19348
rect 14028 19294 14030 19346
rect 14030 19294 14082 19346
rect 14082 19294 14084 19346
rect 14028 19292 14084 19294
rect 14476 19292 14532 19348
rect 14140 19234 14196 19236
rect 14140 19182 14142 19234
rect 14142 19182 14194 19234
rect 14194 19182 14196 19234
rect 14140 19180 14196 19182
rect 14812 19516 14868 19572
rect 13468 18956 13524 19012
rect 13692 18450 13748 18452
rect 13692 18398 13694 18450
rect 13694 18398 13746 18450
rect 13746 18398 13748 18450
rect 13692 18396 13748 18398
rect 12908 18338 12964 18340
rect 12908 18286 12910 18338
rect 12910 18286 12962 18338
rect 12962 18286 12964 18338
rect 12908 18284 12964 18286
rect 13580 18338 13636 18340
rect 13580 18286 13582 18338
rect 13582 18286 13634 18338
rect 13634 18286 13636 18338
rect 13580 18284 13636 18286
rect 13468 17612 13524 17668
rect 14140 18284 14196 18340
rect 15148 21474 15204 21476
rect 15148 21422 15150 21474
rect 15150 21422 15202 21474
rect 15202 21422 15204 21474
rect 15148 21420 15204 21422
rect 15708 20636 15764 20692
rect 15596 20188 15652 20244
rect 14924 18284 14980 18340
rect 15484 20076 15540 20132
rect 15484 19852 15540 19908
rect 15372 19234 15428 19236
rect 15372 19182 15374 19234
rect 15374 19182 15426 19234
rect 15426 19182 15428 19234
rect 15372 19180 15428 19182
rect 15820 20188 15876 20244
rect 15932 19180 15988 19236
rect 16044 19516 16100 19572
rect 15036 17836 15092 17892
rect 15148 19010 15204 19012
rect 15148 18958 15150 19010
rect 15150 18958 15202 19010
rect 15202 18958 15204 19010
rect 15148 18956 15204 18958
rect 15932 19010 15988 19012
rect 15932 18958 15934 19010
rect 15934 18958 15986 19010
rect 15986 18958 15988 19010
rect 15932 18956 15988 18958
rect 4284 16882 4340 16884
rect 4284 16830 4286 16882
rect 4286 16830 4338 16882
rect 4338 16830 4340 16882
rect 4284 16828 4340 16830
rect 11564 16828 11620 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 1932 16156 1988 16212
rect 17724 27858 17780 27860
rect 17724 27806 17726 27858
rect 17726 27806 17778 27858
rect 17778 27806 17780 27858
rect 17724 27804 17780 27806
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 21532 38220 21588 38276
rect 22428 38274 22484 38276
rect 22428 38222 22430 38274
rect 22430 38222 22482 38274
rect 22482 38222 22484 38274
rect 22428 38220 22484 38222
rect 25564 38444 25620 38500
rect 24220 38220 24276 38276
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 20188 37436 20244 37492
rect 21420 37490 21476 37492
rect 21420 37438 21422 37490
rect 21422 37438 21474 37490
rect 21474 37438 21476 37490
rect 21420 37436 21476 37438
rect 18956 29426 19012 29428
rect 18956 29374 18958 29426
rect 18958 29374 19010 29426
rect 19010 29374 19012 29426
rect 18956 29372 19012 29374
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19628 28530 19684 28532
rect 19628 28478 19630 28530
rect 19630 28478 19682 28530
rect 19682 28478 19684 28530
rect 19628 28476 19684 28478
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 18844 27858 18900 27860
rect 18844 27806 18846 27858
rect 18846 27806 18898 27858
rect 18898 27806 18900 27858
rect 18844 27804 18900 27806
rect 19180 27858 19236 27860
rect 19180 27806 19182 27858
rect 19182 27806 19234 27858
rect 19234 27806 19236 27858
rect 19180 27804 19236 27806
rect 17836 27692 17892 27748
rect 18956 27692 19012 27748
rect 17388 25340 17444 25396
rect 16828 23324 16884 23380
rect 16828 22204 16884 22260
rect 16716 21868 16772 21924
rect 16828 21586 16884 21588
rect 16828 21534 16830 21586
rect 16830 21534 16882 21586
rect 16882 21534 16884 21586
rect 16828 21532 16884 21534
rect 16380 20188 16436 20244
rect 16268 20076 16324 20132
rect 16380 19458 16436 19460
rect 16380 19406 16382 19458
rect 16382 19406 16434 19458
rect 16434 19406 16436 19458
rect 16380 19404 16436 19406
rect 17052 23100 17108 23156
rect 17052 22146 17108 22148
rect 17052 22094 17054 22146
rect 17054 22094 17106 22146
rect 17106 22094 17108 22146
rect 17052 22092 17108 22094
rect 17052 21532 17108 21588
rect 16716 20076 16772 20132
rect 16828 19964 16884 20020
rect 16716 19458 16772 19460
rect 16716 19406 16718 19458
rect 16718 19406 16770 19458
rect 16770 19406 16772 19458
rect 16716 19404 16772 19406
rect 17724 24946 17780 24948
rect 17724 24894 17726 24946
rect 17726 24894 17778 24946
rect 17778 24894 17780 24946
rect 17724 24892 17780 24894
rect 21868 29372 21924 29428
rect 20860 27858 20916 27860
rect 20860 27806 20862 27858
rect 20862 27806 20914 27858
rect 20914 27806 20916 27858
rect 20860 27804 20916 27806
rect 22316 29426 22372 29428
rect 22316 29374 22318 29426
rect 22318 29374 22370 29426
rect 22370 29374 22372 29426
rect 22316 29372 22372 29374
rect 23324 27804 23380 27860
rect 18844 24892 18900 24948
rect 19516 24892 19572 24948
rect 17612 23324 17668 23380
rect 17836 23212 17892 23268
rect 19516 23378 19572 23380
rect 19516 23326 19518 23378
rect 19518 23326 19570 23378
rect 19570 23326 19572 23378
rect 19516 23324 19572 23326
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20300 26124 20356 26180
rect 19740 25452 19796 25508
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20188 24946 20244 24948
rect 20188 24894 20190 24946
rect 20190 24894 20242 24946
rect 20242 24894 20244 24946
rect 20188 24892 20244 24894
rect 20300 24722 20356 24724
rect 20300 24670 20302 24722
rect 20302 24670 20354 24722
rect 20354 24670 20356 24722
rect 20300 24668 20356 24670
rect 20748 26178 20804 26180
rect 20748 26126 20750 26178
rect 20750 26126 20802 26178
rect 20802 26126 20804 26178
rect 20748 26124 20804 26126
rect 21644 25452 21700 25508
rect 20748 25228 20804 25284
rect 21532 25004 21588 25060
rect 23212 27692 23268 27748
rect 26236 37884 26292 37940
rect 26796 38444 26852 38500
rect 27468 37938 27524 37940
rect 27468 37886 27470 37938
rect 27470 37886 27522 37938
rect 27522 37886 27524 37938
rect 27468 37884 27524 37886
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 24556 27746 24612 27748
rect 24556 27694 24558 27746
rect 24558 27694 24610 27746
rect 24610 27694 24612 27746
rect 24556 27692 24612 27694
rect 21868 25452 21924 25508
rect 22092 25394 22148 25396
rect 22092 25342 22094 25394
rect 22094 25342 22146 25394
rect 22146 25342 22148 25394
rect 22092 25340 22148 25342
rect 21756 25228 21812 25284
rect 22876 25228 22932 25284
rect 21868 25116 21924 25172
rect 21644 24892 21700 24948
rect 22764 25004 22820 25060
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20188 23436 20244 23492
rect 20300 23324 20356 23380
rect 20188 23266 20244 23268
rect 20188 23214 20190 23266
rect 20190 23214 20242 23266
rect 20242 23214 20244 23266
rect 20188 23212 20244 23214
rect 19068 23154 19124 23156
rect 19068 23102 19070 23154
rect 19070 23102 19122 23154
rect 19122 23102 19124 23154
rect 19068 23100 19124 23102
rect 17836 22428 17892 22484
rect 17388 21980 17444 22036
rect 17612 21868 17668 21924
rect 18284 22316 18340 22372
rect 18396 22204 18452 22260
rect 18172 21868 18228 21924
rect 19180 22594 19236 22596
rect 19180 22542 19182 22594
rect 19182 22542 19234 22594
rect 19234 22542 19236 22594
rect 19180 22540 19236 22542
rect 20300 22876 20356 22932
rect 18732 22204 18788 22260
rect 18620 21868 18676 21924
rect 18956 21868 19012 21924
rect 18508 21756 18564 21812
rect 18284 21586 18340 21588
rect 18284 21534 18286 21586
rect 18286 21534 18338 21586
rect 18338 21534 18340 21586
rect 18284 21532 18340 21534
rect 18844 20188 18900 20244
rect 19628 22370 19684 22372
rect 19628 22318 19630 22370
rect 19630 22318 19682 22370
rect 19682 22318 19684 22370
rect 19628 22316 19684 22318
rect 19068 20524 19124 20580
rect 19068 20130 19124 20132
rect 19068 20078 19070 20130
rect 19070 20078 19122 20130
rect 19122 20078 19124 20130
rect 19068 20076 19124 20078
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 21532 24834 21588 24836
rect 21532 24782 21534 24834
rect 21534 24782 21586 24834
rect 21586 24782 21588 24834
rect 21532 24780 21588 24782
rect 20524 22540 20580 22596
rect 20300 21868 20356 21924
rect 20300 21644 20356 21700
rect 20300 20524 20356 20580
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19964 20188 20020 20244
rect 19740 20076 19796 20132
rect 17948 20018 18004 20020
rect 17948 19966 17950 20018
rect 17950 19966 18002 20018
rect 18002 19966 18004 20018
rect 17948 19964 18004 19966
rect 18956 19964 19012 20020
rect 17724 19852 17780 19908
rect 17500 19404 17556 19460
rect 18620 19458 18676 19460
rect 18620 19406 18622 19458
rect 18622 19406 18674 19458
rect 18674 19406 18676 19458
rect 18620 19404 18676 19406
rect 17388 19180 17444 19236
rect 19852 20018 19908 20020
rect 19852 19966 19854 20018
rect 19854 19966 19906 20018
rect 19906 19966 19908 20018
rect 19852 19964 19908 19966
rect 19628 19516 19684 19572
rect 19180 19404 19236 19460
rect 20076 20076 20132 20132
rect 20412 19404 20468 19460
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20188 18732 20244 18788
rect 19404 18674 19460 18676
rect 19404 18622 19406 18674
rect 19406 18622 19458 18674
rect 19458 18622 19460 18674
rect 19404 18620 19460 18622
rect 18956 18508 19012 18564
rect 17836 18172 17892 18228
rect 18060 17612 18116 17668
rect 14924 16828 14980 16884
rect 15484 16882 15540 16884
rect 15484 16830 15486 16882
rect 15486 16830 15538 16882
rect 15538 16830 15540 16882
rect 15484 16828 15540 16830
rect 16044 17442 16100 17444
rect 16044 17390 16046 17442
rect 16046 17390 16098 17442
rect 16098 17390 16100 17442
rect 16044 17388 16100 17390
rect 16268 17276 16324 17332
rect 13020 15036 13076 15092
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 15036 16098 15092 16100
rect 15036 16046 15038 16098
rect 15038 16046 15090 16098
rect 15090 16046 15092 16098
rect 15036 16044 15092 16046
rect 13468 15036 13524 15092
rect 13804 15148 13860 15204
rect 15484 16044 15540 16100
rect 15932 16044 15988 16100
rect 16156 16044 16212 16100
rect 15484 15202 15540 15204
rect 15484 15150 15486 15202
rect 15486 15150 15538 15202
rect 15538 15150 15540 15202
rect 15484 15148 15540 15150
rect 14364 15036 14420 15092
rect 14700 14642 14756 14644
rect 14700 14590 14702 14642
rect 14702 14590 14754 14642
rect 14754 14590 14756 14642
rect 14700 14588 14756 14590
rect 15596 14588 15652 14644
rect 17724 17388 17780 17444
rect 17836 16044 17892 16100
rect 20412 18732 20468 18788
rect 20412 18508 20468 18564
rect 19852 17442 19908 17444
rect 19852 17390 19854 17442
rect 19854 17390 19906 17442
rect 19906 17390 19908 17442
rect 19852 17388 19908 17390
rect 20860 23436 20916 23492
rect 21644 24610 21700 24612
rect 21644 24558 21646 24610
rect 21646 24558 21698 24610
rect 21698 24558 21700 24610
rect 21644 24556 21700 24558
rect 20748 21532 20804 21588
rect 20636 19794 20692 19796
rect 20636 19742 20638 19794
rect 20638 19742 20690 19794
rect 20690 19742 20692 19794
rect 20636 19740 20692 19742
rect 20972 22092 21028 22148
rect 20972 21868 21028 21924
rect 20524 18396 20580 18452
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 18732 16828 18788 16884
rect 17388 15426 17444 15428
rect 17388 15374 17390 15426
rect 17390 15374 17442 15426
rect 17442 15374 17444 15426
rect 17388 15372 17444 15374
rect 17612 15820 17668 15876
rect 16380 15148 16436 15204
rect 18060 15372 18116 15428
rect 20860 18508 20916 18564
rect 22428 24892 22484 24948
rect 22428 23884 22484 23940
rect 22540 23324 22596 23380
rect 21084 21532 21140 21588
rect 21308 22988 21364 23044
rect 21084 20130 21140 20132
rect 21084 20078 21086 20130
rect 21086 20078 21138 20130
rect 21138 20078 21140 20130
rect 21084 20076 21140 20078
rect 21196 18508 21252 18564
rect 21756 23042 21812 23044
rect 21756 22990 21758 23042
rect 21758 22990 21810 23042
rect 21810 22990 21812 23042
rect 21756 22988 21812 22990
rect 21756 21698 21812 21700
rect 21756 21646 21758 21698
rect 21758 21646 21810 21698
rect 21810 21646 21812 21698
rect 21756 21644 21812 21646
rect 22988 24610 23044 24612
rect 22988 24558 22990 24610
rect 22990 24558 23042 24610
rect 23042 24558 23044 24610
rect 22988 24556 23044 24558
rect 23660 25452 23716 25508
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 25228 25452 25284 25508
rect 26236 25452 26292 25508
rect 26124 25394 26180 25396
rect 26124 25342 26126 25394
rect 26126 25342 26178 25394
rect 26178 25342 26180 25394
rect 26124 25340 26180 25342
rect 28140 25452 28196 25508
rect 25340 24892 25396 24948
rect 22764 23548 22820 23604
rect 23436 23548 23492 23604
rect 22876 21532 22932 21588
rect 21644 20578 21700 20580
rect 21644 20526 21646 20578
rect 21646 20526 21698 20578
rect 21698 20526 21700 20578
rect 21644 20524 21700 20526
rect 21868 20188 21924 20244
rect 21756 20076 21812 20132
rect 22652 20748 22708 20804
rect 22428 20690 22484 20692
rect 22428 20638 22430 20690
rect 22430 20638 22482 20690
rect 22482 20638 22484 20690
rect 22428 20636 22484 20638
rect 22764 21308 22820 21364
rect 21868 19458 21924 19460
rect 21868 19406 21870 19458
rect 21870 19406 21922 19458
rect 21922 19406 21924 19458
rect 21868 19404 21924 19406
rect 21420 18620 21476 18676
rect 22092 19516 22148 19572
rect 22652 20130 22708 20132
rect 22652 20078 22654 20130
rect 22654 20078 22706 20130
rect 22706 20078 22708 20130
rect 22652 20076 22708 20078
rect 24444 23212 24500 23268
rect 24332 22092 24388 22148
rect 24220 21362 24276 21364
rect 24220 21310 24222 21362
rect 24222 21310 24274 21362
rect 24274 21310 24276 21362
rect 24220 21308 24276 21310
rect 23212 20636 23268 20692
rect 23100 19906 23156 19908
rect 23100 19854 23102 19906
rect 23102 19854 23154 19906
rect 23154 19854 23156 19906
rect 23100 19852 23156 19854
rect 23884 20748 23940 20804
rect 24668 23154 24724 23156
rect 24668 23102 24670 23154
rect 24670 23102 24722 23154
rect 24722 23102 24724 23154
rect 24668 23100 24724 23102
rect 25676 23938 25732 23940
rect 25676 23886 25678 23938
rect 25678 23886 25730 23938
rect 25730 23886 25732 23938
rect 25676 23884 25732 23886
rect 26796 24892 26852 24948
rect 37660 25506 37716 25508
rect 37660 25454 37662 25506
rect 37662 25454 37714 25506
rect 37714 25454 37716 25506
rect 37660 25452 37716 25454
rect 28588 24946 28644 24948
rect 28588 24894 28590 24946
rect 28590 24894 28642 24946
rect 28642 24894 28644 24946
rect 28588 24892 28644 24894
rect 40012 24892 40068 24948
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 25340 23100 25396 23156
rect 25004 21756 25060 21812
rect 25452 23436 25508 23492
rect 26796 23436 26852 23492
rect 26684 23324 26740 23380
rect 26572 23266 26628 23268
rect 26572 23214 26574 23266
rect 26574 23214 26626 23266
rect 26626 23214 26628 23266
rect 26572 23212 26628 23214
rect 28140 23212 28196 23268
rect 25452 21868 25508 21924
rect 24108 20690 24164 20692
rect 24108 20638 24110 20690
rect 24110 20638 24162 20690
rect 24162 20638 24164 20690
rect 24108 20636 24164 20638
rect 23436 19740 23492 19796
rect 22652 19404 22708 19460
rect 22540 18732 22596 18788
rect 22876 18620 22932 18676
rect 24220 20130 24276 20132
rect 24220 20078 24222 20130
rect 24222 20078 24274 20130
rect 24274 20078 24276 20130
rect 24220 20076 24276 20078
rect 23548 18620 23604 18676
rect 21420 18450 21476 18452
rect 21420 18398 21422 18450
rect 21422 18398 21474 18450
rect 21474 18398 21476 18450
rect 21420 18396 21476 18398
rect 21308 18172 21364 18228
rect 21532 18284 21588 18340
rect 20972 17388 21028 17444
rect 21868 17890 21924 17892
rect 21868 17838 21870 17890
rect 21870 17838 21922 17890
rect 21922 17838 21924 17890
rect 21868 17836 21924 17838
rect 21868 17666 21924 17668
rect 21868 17614 21870 17666
rect 21870 17614 21922 17666
rect 21922 17614 21924 17666
rect 21868 17612 21924 17614
rect 21756 17442 21812 17444
rect 21756 17390 21758 17442
rect 21758 17390 21810 17442
rect 21810 17390 21812 17442
rect 21756 17388 21812 17390
rect 19180 16044 19236 16100
rect 16268 14588 16324 14644
rect 17836 15202 17892 15204
rect 17836 15150 17838 15202
rect 17838 15150 17890 15202
rect 17890 15150 17892 15202
rect 17836 15148 17892 15150
rect 17612 14588 17668 14644
rect 16828 13692 16884 13748
rect 17500 13746 17556 13748
rect 17500 13694 17502 13746
rect 17502 13694 17554 13746
rect 17554 13694 17556 13746
rect 17500 13692 17556 13694
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 16156 5180 16212 5236
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 17388 5234 17444 5236
rect 17388 5182 17390 5234
rect 17390 5182 17442 5234
rect 17442 5182 17444 5234
rect 17388 5180 17444 5182
rect 18508 14642 18564 14644
rect 18508 14590 18510 14642
rect 18510 14590 18562 14642
rect 18562 14590 18564 14642
rect 18508 14588 18564 14590
rect 20748 16210 20804 16212
rect 20748 16158 20750 16210
rect 20750 16158 20802 16210
rect 20802 16158 20804 16210
rect 20748 16156 20804 16158
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 21644 17106 21700 17108
rect 21644 17054 21646 17106
rect 21646 17054 21698 17106
rect 21698 17054 21700 17106
rect 21644 17052 21700 17054
rect 22988 17052 23044 17108
rect 25004 20188 25060 20244
rect 24556 20130 24612 20132
rect 24556 20078 24558 20130
rect 24558 20078 24610 20130
rect 24610 20078 24612 20130
rect 24556 20076 24612 20078
rect 25564 20018 25620 20020
rect 25564 19966 25566 20018
rect 25566 19966 25618 20018
rect 25618 19966 25620 20018
rect 25564 19964 25620 19966
rect 25676 19906 25732 19908
rect 25676 19854 25678 19906
rect 25678 19854 25730 19906
rect 25730 19854 25732 19906
rect 25676 19852 25732 19854
rect 26572 21868 26628 21924
rect 25900 20188 25956 20244
rect 26124 20076 26180 20132
rect 26460 20018 26516 20020
rect 26460 19966 26462 20018
rect 26462 19966 26514 20018
rect 26514 19966 26516 20018
rect 26460 19964 26516 19966
rect 26348 19852 26404 19908
rect 37660 22988 37716 23044
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 40012 22204 40068 22260
rect 37660 21586 37716 21588
rect 37660 21534 37662 21586
rect 37662 21534 37714 21586
rect 37714 21534 37716 21586
rect 37660 21532 37716 21534
rect 40012 21532 40068 21588
rect 28252 21420 28308 21476
rect 29148 21474 29204 21476
rect 29148 21422 29150 21474
rect 29150 21422 29202 21474
rect 29202 21422 29204 21474
rect 29148 21420 29204 21422
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 27916 20860 27972 20916
rect 28588 20914 28644 20916
rect 28588 20862 28590 20914
rect 28590 20862 28642 20914
rect 28642 20862 28644 20914
rect 28588 20860 28644 20862
rect 40012 20914 40068 20916
rect 40012 20862 40014 20914
rect 40014 20862 40066 20914
rect 40066 20862 40068 20914
rect 40012 20860 40068 20862
rect 37660 20802 37716 20804
rect 37660 20750 37662 20802
rect 37662 20750 37714 20802
rect 37714 20750 37716 20802
rect 37660 20748 37716 20750
rect 27804 20018 27860 20020
rect 27804 19966 27806 20018
rect 27806 19966 27858 20018
rect 27858 19966 27860 20018
rect 27804 19964 27860 19966
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 24780 18284 24836 18340
rect 24332 17836 24388 17892
rect 22764 16156 22820 16212
rect 21532 15820 21588 15876
rect 20300 15314 20356 15316
rect 20300 15262 20302 15314
rect 20302 15262 20354 15314
rect 20354 15262 20356 15314
rect 20300 15260 20356 15262
rect 25788 18284 25844 18340
rect 25228 17388 25284 17444
rect 26684 17836 26740 17892
rect 26124 17554 26180 17556
rect 26124 17502 26126 17554
rect 26126 17502 26178 17554
rect 26178 17502 26180 17554
rect 26124 17500 26180 17502
rect 37660 18450 37716 18452
rect 37660 18398 37662 18450
rect 37662 18398 37714 18450
rect 37714 18398 37716 18450
rect 37660 18396 37716 18398
rect 27804 18284 27860 18340
rect 27692 17890 27748 17892
rect 27692 17838 27694 17890
rect 27694 17838 27746 17890
rect 27746 17838 27748 17890
rect 27692 17836 27748 17838
rect 28700 18338 28756 18340
rect 28700 18286 28702 18338
rect 28702 18286 28754 18338
rect 28754 18286 28756 18338
rect 28700 18284 28756 18286
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 27132 17666 27188 17668
rect 27132 17614 27134 17666
rect 27134 17614 27186 17666
rect 27186 17614 27188 17666
rect 27132 17612 27188 17614
rect 28140 17612 28196 17668
rect 26796 17500 26852 17556
rect 26236 17388 26292 17444
rect 27020 17442 27076 17444
rect 27020 17390 27022 17442
rect 27022 17390 27074 17442
rect 27074 17390 27076 17442
rect 27020 17388 27076 17390
rect 25228 16882 25284 16884
rect 25228 16830 25230 16882
rect 25230 16830 25282 16882
rect 25282 16830 25284 16882
rect 25228 16828 25284 16830
rect 37660 17666 37716 17668
rect 37660 17614 37662 17666
rect 37662 17614 37714 17666
rect 37714 17614 37716 17666
rect 37660 17612 37716 17614
rect 28588 16882 28644 16884
rect 28588 16830 28590 16882
rect 28590 16830 28642 16882
rect 28642 16830 28644 16882
rect 28588 16828 28644 16830
rect 40012 16828 40068 16884
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 24220 15314 24276 15316
rect 24220 15262 24222 15314
rect 24222 15262 24274 15314
rect 24274 15262 24276 15314
rect 24220 15260 24276 15262
rect 24780 15260 24836 15316
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 19068 14306 19124 14308
rect 19068 14254 19070 14306
rect 19070 14254 19122 14306
rect 19122 14254 19124 14306
rect 19068 14252 19124 14254
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19628 13692 19684 13748
rect 19852 13692 19908 13748
rect 20412 13692 20468 13748
rect 20188 12738 20244 12740
rect 20188 12686 20190 12738
rect 20190 12686 20242 12738
rect 20242 12686 20244 12738
rect 20188 12684 20244 12686
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 20972 13746 21028 13748
rect 20972 13694 20974 13746
rect 20974 13694 21026 13746
rect 21026 13694 21028 13746
rect 20972 13692 21028 13694
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 20860 12684 20916 12740
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20188 4060 20244 4116
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 20860 3612 20916 3668
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 40236 10780 40292 10836
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 21420 4114 21476 4116
rect 21420 4062 21422 4114
rect 21422 4062 21474 4114
rect 21474 4062 21476 4114
rect 21420 4060 21476 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 22092 3666 22148 3668
rect 22092 3614 22094 3666
rect 22094 3614 22146 3666
rect 22146 3614 22148 3666
rect 22092 3612 22148 3614
<< metal3 >>
rect 25554 38444 25564 38500
rect 25620 38444 26796 38500
rect 26852 38444 26862 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 21522 38220 21532 38276
rect 21588 38220 22428 38276
rect 22484 38220 22494 38276
rect 24210 38220 24220 38276
rect 24276 38220 25564 38276
rect 25620 38220 25630 38276
rect 26226 37884 26236 37940
rect 26292 37884 27468 37940
rect 27524 37884 27534 37940
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 20178 37436 20188 37492
rect 20244 37436 21420 37492
rect 21476 37436 21486 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 16146 36652 16156 36708
rect 16212 36652 17388 36708
rect 17444 36652 17454 36708
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 18946 29372 18956 29428
rect 19012 29372 21868 29428
rect 21924 29372 22316 29428
rect 22372 29372 22382 29428
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 16370 28476 16380 28532
rect 16436 28476 16828 28532
rect 16884 28476 19628 28532
rect 19684 28476 19694 28532
rect 0 28308 800 28336
rect 0 28252 4172 28308
rect 4228 28252 4238 28308
rect 0 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 17714 27804 17724 27860
rect 17780 27804 18844 27860
rect 18900 27804 18910 27860
rect 19170 27804 19180 27860
rect 19236 27804 20860 27860
rect 20916 27804 23324 27860
rect 23380 27804 23390 27860
rect 17378 27692 17388 27748
rect 17444 27692 17836 27748
rect 17892 27692 18956 27748
rect 19012 27692 19022 27748
rect 23202 27692 23212 27748
rect 23268 27692 24556 27748
rect 24612 27692 24622 27748
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 13570 26908 13580 26964
rect 13636 26908 14812 26964
rect 14868 26908 14878 26964
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 4274 26236 4284 26292
rect 4340 26236 12012 26292
rect 12068 26236 12078 26292
rect 14242 26124 14252 26180
rect 14308 26124 15820 26180
rect 15876 26124 15886 26180
rect 20290 26124 20300 26180
rect 20356 26124 20748 26180
rect 20804 26124 20814 26180
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 0 25620 800 25648
rect 0 25564 1932 25620
rect 1988 25564 1998 25620
rect 0 25536 800 25564
rect 19730 25452 19740 25508
rect 19796 25452 21644 25508
rect 21700 25452 21868 25508
rect 21924 25452 21934 25508
rect 23650 25452 23660 25508
rect 23716 25452 25228 25508
rect 25284 25452 25294 25508
rect 26226 25452 26236 25508
rect 26292 25452 28140 25508
rect 28196 25452 37660 25508
rect 37716 25452 37726 25508
rect 12002 25340 12012 25396
rect 12068 25340 15372 25396
rect 15428 25340 15438 25396
rect 17378 25340 17388 25396
rect 17444 25340 22092 25396
rect 22148 25340 26124 25396
rect 26180 25340 26190 25396
rect 14354 25228 14364 25284
rect 14420 25228 20580 25284
rect 20738 25228 20748 25284
rect 20804 25228 21756 25284
rect 21812 25228 22876 25284
rect 22932 25228 23548 25284
rect 20524 25172 20580 25228
rect 20524 25116 21868 25172
rect 21924 25116 21934 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 21522 25004 21532 25060
rect 21588 25004 22764 25060
rect 22820 25004 22830 25060
rect 23492 24948 23548 25228
rect 41200 24948 42000 24976
rect 15474 24892 15484 24948
rect 15540 24892 16044 24948
rect 16100 24892 17724 24948
rect 17780 24892 18844 24948
rect 18900 24892 18910 24948
rect 19506 24892 19516 24948
rect 19572 24892 20188 24948
rect 20244 24892 20254 24948
rect 21634 24892 21644 24948
rect 21700 24892 22428 24948
rect 22484 24892 22494 24948
rect 23492 24892 25340 24948
rect 25396 24892 26796 24948
rect 26852 24892 28588 24948
rect 28644 24892 28654 24948
rect 40002 24892 40012 24948
rect 40068 24892 42000 24948
rect 41200 24864 42000 24892
rect 14578 24780 14588 24836
rect 14644 24780 21532 24836
rect 21588 24780 21598 24836
rect 4274 24668 4284 24724
rect 4340 24668 8428 24724
rect 16594 24668 16604 24724
rect 16660 24668 20300 24724
rect 20356 24668 20366 24724
rect 1922 24444 1932 24500
rect 1988 24444 1998 24500
rect 0 24276 800 24304
rect 1932 24276 1988 24444
rect 8372 24388 8428 24668
rect 21634 24556 21644 24612
rect 21700 24556 22988 24612
rect 23044 24556 23054 24612
rect 13794 24444 13804 24500
rect 13860 24444 15484 24500
rect 15540 24444 15550 24500
rect 8372 24332 10556 24388
rect 10612 24332 13916 24388
rect 13972 24332 13982 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 0 24220 1988 24276
rect 0 24192 800 24220
rect 12338 23884 12348 23940
rect 12404 23884 13804 23940
rect 13860 23884 13870 23940
rect 22418 23884 22428 23940
rect 22484 23884 25676 23940
rect 25732 23884 25742 23940
rect 14354 23772 14364 23828
rect 14420 23772 16268 23828
rect 16324 23772 16334 23828
rect 22754 23548 22764 23604
rect 22820 23548 23436 23604
rect 23492 23548 23502 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 20178 23436 20188 23492
rect 20244 23436 20860 23492
rect 20916 23436 20926 23492
rect 25442 23436 25452 23492
rect 25508 23436 26796 23492
rect 26852 23436 26862 23492
rect 16818 23324 16828 23380
rect 16884 23324 17612 23380
rect 17668 23324 17678 23380
rect 19506 23324 19516 23380
rect 19572 23324 20300 23380
rect 20356 23324 20366 23380
rect 22530 23324 22540 23380
rect 22596 23324 26684 23380
rect 26740 23324 26750 23380
rect 17826 23212 17836 23268
rect 17892 23212 20188 23268
rect 20244 23212 24444 23268
rect 24500 23212 24510 23268
rect 26562 23212 26572 23268
rect 26628 23212 28140 23268
rect 28196 23212 28206 23268
rect 16482 23100 16492 23156
rect 16548 23100 17052 23156
rect 17108 23100 19068 23156
rect 19124 23100 19134 23156
rect 24658 23100 24668 23156
rect 24724 23100 25340 23156
rect 25396 23100 25406 23156
rect 10658 22988 10668 23044
rect 10724 22988 16380 23044
rect 16436 22988 16446 23044
rect 21298 22988 21308 23044
rect 21364 22988 21756 23044
rect 21812 22988 37660 23044
rect 37716 22988 37726 23044
rect 16146 22876 16156 22932
rect 16212 22876 20300 22932
rect 20356 22876 20366 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 14130 22540 14140 22596
rect 14196 22540 14812 22596
rect 14868 22540 15148 22596
rect 19170 22540 19180 22596
rect 19236 22540 20524 22596
rect 20580 22540 20590 22596
rect 15092 22372 15148 22540
rect 16258 22428 16268 22484
rect 16324 22428 17836 22484
rect 17892 22428 17902 22484
rect 15092 22316 18284 22372
rect 18340 22316 19628 22372
rect 19684 22316 19694 22372
rect 41200 22260 42000 22288
rect 16818 22204 16828 22260
rect 16884 22204 18396 22260
rect 18452 22204 18732 22260
rect 18788 22204 18798 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 41200 22176 42000 22204
rect 4162 22092 4172 22148
rect 4228 22092 17052 22148
rect 17108 22092 17118 22148
rect 20962 22092 20972 22148
rect 21028 22092 24332 22148
rect 24388 22092 24398 22148
rect 15820 21980 17388 22036
rect 17444 21980 17454 22036
rect 15820 21924 15876 21980
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 15810 21868 15820 21924
rect 15876 21868 15886 21924
rect 16706 21868 16716 21924
rect 16772 21868 17612 21924
rect 17668 21868 17678 21924
rect 18162 21868 18172 21924
rect 18228 21868 18620 21924
rect 18676 21868 18956 21924
rect 19012 21868 19022 21924
rect 20290 21868 20300 21924
rect 20356 21868 20972 21924
rect 21028 21868 21038 21924
rect 25442 21868 25452 21924
rect 25508 21868 26572 21924
rect 26628 21868 26638 21924
rect 18498 21756 18508 21812
rect 18564 21756 25004 21812
rect 25060 21756 25070 21812
rect 20290 21644 20300 21700
rect 20356 21644 21756 21700
rect 21812 21644 21822 21700
rect 41200 21588 42000 21616
rect 15810 21532 15820 21588
rect 15876 21532 16828 21588
rect 16884 21532 16894 21588
rect 17042 21532 17052 21588
rect 17108 21532 18284 21588
rect 18340 21532 18350 21588
rect 20738 21532 20748 21588
rect 20804 21532 21084 21588
rect 21140 21532 22876 21588
rect 22932 21532 22942 21588
rect 31892 21532 37660 21588
rect 37716 21532 37726 21588
rect 40002 21532 40012 21588
rect 40068 21532 42000 21588
rect 31892 21476 31948 21532
rect 41200 21504 42000 21532
rect 14130 21420 14140 21476
rect 14196 21420 15148 21476
rect 15204 21420 15214 21476
rect 28242 21420 28252 21476
rect 28308 21420 29148 21476
rect 29204 21420 31948 21476
rect 22754 21308 22764 21364
rect 22820 21308 24220 21364
rect 24276 21308 24286 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 41200 20916 42000 20944
rect 27906 20860 27916 20916
rect 27972 20860 28588 20916
rect 28644 20860 31948 20916
rect 40002 20860 40012 20916
rect 40068 20860 42000 20916
rect 31892 20804 31948 20860
rect 41200 20832 42000 20860
rect 22642 20748 22652 20804
rect 22708 20748 23884 20804
rect 23940 20748 23950 20804
rect 31892 20748 37660 20804
rect 37716 20748 37726 20804
rect 15698 20636 15708 20692
rect 15764 20636 22428 20692
rect 22484 20636 22494 20692
rect 23202 20636 23212 20692
rect 23268 20636 24108 20692
rect 24164 20636 24174 20692
rect 19058 20524 19068 20580
rect 19124 20524 20300 20580
rect 20356 20524 21644 20580
rect 21700 20524 21710 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 15092 20188 15596 20244
rect 15652 20188 15662 20244
rect 15810 20188 15820 20244
rect 15876 20188 16380 20244
rect 16436 20188 16446 20244
rect 18834 20188 18844 20244
rect 18900 20188 19964 20244
rect 20020 20188 21868 20244
rect 21924 20188 21934 20244
rect 24994 20188 25004 20244
rect 25060 20188 25900 20244
rect 25956 20188 25966 20244
rect 15092 20132 15148 20188
rect 18844 20132 18900 20188
rect 14130 20076 14140 20132
rect 14196 20076 15148 20132
rect 15474 20076 15484 20132
rect 15540 20076 16268 20132
rect 16324 20076 16334 20132
rect 16706 20076 16716 20132
rect 16772 20076 18900 20132
rect 19058 20076 19068 20132
rect 19124 20076 19740 20132
rect 19796 20076 20076 20132
rect 20132 20076 21084 20132
rect 21140 20076 21150 20132
rect 21746 20076 21756 20132
rect 21812 20076 22652 20132
rect 22708 20076 24220 20132
rect 24276 20076 24286 20132
rect 24546 20076 24556 20132
rect 24612 20076 26124 20132
rect 26180 20076 26190 20132
rect 9986 19964 9996 20020
rect 10052 19964 12684 20020
rect 12740 19964 13244 20020
rect 13300 19964 16828 20020
rect 16884 19964 16894 20020
rect 10658 19852 10668 19908
rect 10724 19852 14028 19908
rect 14084 19852 14094 19908
rect 14690 19852 14700 19908
rect 14756 19852 15484 19908
rect 15540 19852 15550 19908
rect 17052 19796 17108 20076
rect 17938 19964 17948 20020
rect 18004 19964 18956 20020
rect 19012 19964 19852 20020
rect 19908 19964 19918 20020
rect 20076 19964 25564 20020
rect 25620 19964 25630 20020
rect 26450 19964 26460 20020
rect 26516 19964 27804 20020
rect 27860 19964 27870 20020
rect 20076 19908 20132 19964
rect 17714 19852 17724 19908
rect 17780 19852 20132 19908
rect 23090 19852 23100 19908
rect 23156 19852 25676 19908
rect 25732 19852 26348 19908
rect 26404 19852 26414 19908
rect 13458 19740 13468 19796
rect 13524 19740 17108 19796
rect 17724 19684 17780 19852
rect 20626 19740 20636 19796
rect 20692 19740 23436 19796
rect 23492 19740 23502 19796
rect 13906 19628 13916 19684
rect 13972 19628 17780 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 14802 19516 14812 19572
rect 14868 19516 16044 19572
rect 16100 19516 19628 19572
rect 19684 19516 22092 19572
rect 22148 19516 22158 19572
rect 13122 19404 13132 19460
rect 13188 19404 13692 19460
rect 13748 19404 16380 19460
rect 16436 19404 16446 19460
rect 16706 19404 16716 19460
rect 16772 19404 17500 19460
rect 17556 19404 18620 19460
rect 18676 19404 18686 19460
rect 19170 19404 19180 19460
rect 19236 19404 20412 19460
rect 20468 19404 20478 19460
rect 21858 19404 21868 19460
rect 21924 19404 22652 19460
rect 22708 19404 22718 19460
rect 12786 19292 12796 19348
rect 12852 19292 14028 19348
rect 14084 19292 14476 19348
rect 14532 19292 14542 19348
rect 14130 19180 14140 19236
rect 14196 19180 15372 19236
rect 15428 19180 15932 19236
rect 15988 19180 17388 19236
rect 17444 19180 17454 19236
rect 13458 18956 13468 19012
rect 13524 18956 15148 19012
rect 15204 18956 15932 19012
rect 15988 18956 15998 19012
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 20178 18732 20188 18788
rect 20244 18732 20412 18788
rect 20468 18732 22540 18788
rect 22596 18732 22606 18788
rect 11666 18620 11676 18676
rect 11732 18620 12572 18676
rect 12628 18620 12638 18676
rect 19394 18620 19404 18676
rect 19460 18620 21420 18676
rect 21476 18620 22876 18676
rect 22932 18620 23548 18676
rect 23604 18620 23614 18676
rect 18946 18508 18956 18564
rect 19012 18508 20412 18564
rect 20468 18508 20860 18564
rect 20916 18508 21196 18564
rect 21252 18508 21262 18564
rect 4274 18396 4284 18452
rect 4340 18396 9884 18452
rect 9940 18396 13692 18452
rect 13748 18396 13758 18452
rect 20514 18396 20524 18452
rect 20580 18396 21420 18452
rect 21476 18396 21486 18452
rect 31892 18396 37660 18452
rect 37716 18396 37726 18452
rect 31892 18340 31948 18396
rect 12898 18284 12908 18340
rect 12964 18284 13580 18340
rect 13636 18284 13646 18340
rect 14130 18284 14140 18340
rect 14196 18284 14924 18340
rect 14980 18284 21532 18340
rect 21588 18284 21598 18340
rect 24770 18284 24780 18340
rect 24836 18284 25788 18340
rect 25844 18284 25854 18340
rect 27794 18284 27804 18340
rect 27860 18284 28700 18340
rect 28756 18284 31948 18340
rect 0 18228 800 18256
rect 41200 18228 42000 18256
rect 0 18172 1932 18228
rect 1988 18172 1998 18228
rect 17826 18172 17836 18228
rect 17892 18172 21308 18228
rect 21364 18172 21374 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 0 18144 800 18172
rect 41200 18144 42000 18172
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 15026 17836 15036 17892
rect 1922 17724 1932 17780
rect 1988 17724 1998 17780
rect 0 17556 800 17584
rect 1932 17556 1988 17724
rect 4274 17612 4284 17668
rect 4340 17612 13468 17668
rect 13524 17612 13534 17668
rect 0 17500 1988 17556
rect 0 17472 800 17500
rect 15092 17444 15148 17892
rect 21858 17836 21868 17892
rect 21924 17836 24332 17892
rect 24388 17836 24398 17892
rect 26674 17836 26684 17892
rect 26740 17836 27692 17892
rect 27748 17836 27758 17892
rect 18050 17612 18060 17668
rect 18116 17612 21868 17668
rect 21924 17612 21934 17668
rect 27122 17612 27132 17668
rect 27188 17612 28140 17668
rect 28196 17612 37660 17668
rect 37716 17612 37726 17668
rect 26114 17500 26124 17556
rect 26180 17500 26796 17556
rect 26852 17500 26862 17556
rect 15092 17388 16044 17444
rect 16100 17388 17724 17444
rect 17780 17388 17790 17444
rect 17948 17388 19852 17444
rect 19908 17388 20972 17444
rect 21028 17388 21038 17444
rect 21746 17388 21756 17444
rect 21812 17388 25228 17444
rect 25284 17388 25294 17444
rect 26226 17388 26236 17444
rect 26292 17388 27020 17444
rect 27076 17388 27086 17444
rect 17948 17332 18004 17388
rect 16258 17276 16268 17332
rect 16324 17276 18004 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 21634 17052 21644 17108
rect 21700 17052 22988 17108
rect 23044 17052 23054 17108
rect 41200 16884 42000 16912
rect 4274 16828 4284 16884
rect 4340 16828 11564 16884
rect 11620 16828 14924 16884
rect 14980 16828 14990 16884
rect 15474 16828 15484 16884
rect 15540 16828 18732 16884
rect 18788 16828 18798 16884
rect 25218 16828 25228 16884
rect 25284 16828 28588 16884
rect 28644 16828 28654 16884
rect 40002 16828 40012 16884
rect 40068 16828 42000 16884
rect 41200 16800 42000 16828
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 0 16212 800 16240
rect 0 16156 1932 16212
rect 1988 16156 1998 16212
rect 20738 16156 20748 16212
rect 20804 16156 22764 16212
rect 22820 16156 22830 16212
rect 0 16128 800 16156
rect 15026 16044 15036 16100
rect 15092 16044 15484 16100
rect 15540 16044 15932 16100
rect 15988 16044 15998 16100
rect 16146 16044 16156 16100
rect 16212 16044 17836 16100
rect 17892 16044 19180 16100
rect 19236 16044 19246 16100
rect 17602 15820 17612 15876
rect 17668 15820 21532 15876
rect 21588 15820 21598 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 17378 15372 17388 15428
rect 17444 15372 18060 15428
rect 18116 15372 18126 15428
rect 20290 15260 20300 15316
rect 20356 15260 24220 15316
rect 24276 15260 24780 15316
rect 24836 15260 24846 15316
rect 13794 15148 13804 15204
rect 13860 15148 15484 15204
rect 15540 15148 15550 15204
rect 16370 15148 16380 15204
rect 16436 15148 17836 15204
rect 17892 15148 17902 15204
rect 13010 15036 13020 15092
rect 13076 15036 13468 15092
rect 13524 15036 14364 15092
rect 14420 15036 14430 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 14690 14588 14700 14644
rect 14756 14588 15596 14644
rect 15652 14588 16268 14644
rect 16324 14588 16334 14644
rect 17602 14588 17612 14644
rect 17668 14588 18508 14644
rect 18564 14588 18574 14644
rect 19058 14252 19068 14308
rect 19124 14252 20244 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 20188 13748 20244 14252
rect 16818 13692 16828 13748
rect 16884 13692 17500 13748
rect 17556 13692 19628 13748
rect 19684 13692 19694 13748
rect 19842 13692 19852 13748
rect 19908 13692 20412 13748
rect 20468 13692 20972 13748
rect 21028 13692 21038 13748
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 20178 12684 20188 12740
rect 20244 12684 20860 12740
rect 20916 12684 20926 12740
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 41200 10836 42000 10864
rect 40226 10780 40236 10836
rect 40292 10780 42000 10836
rect 41200 10752 42000 10780
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 16146 5180 16156 5236
rect 16212 5180 17388 5236
rect 17444 5180 17454 5236
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 20178 4060 20188 4116
rect 20244 4060 21420 4116
rect 21476 4060 21486 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 20850 3612 20860 3668
rect 20916 3612 22092 3668
rect 22148 3612 22158 3668
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22064 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23296 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _105_
timestamp 1698175906
transform 1 0 13216 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15008 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _107_
timestamp 1698175906
transform 1 0 15120 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16352 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_
timestamp 1698175906
transform -1 0 20944 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21840 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19376 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_
timestamp 1698175906
transform 1 0 14336 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _114_
timestamp 1698175906
transform 1 0 12768 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15904 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17808 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16128 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _118_
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform -1 0 15680 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _120_
timestamp 1698175906
transform 1 0 14000 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _121_
timestamp 1698175906
transform -1 0 16240 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _122_
timestamp 1698175906
transform 1 0 15232 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16912 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14336 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _125_
timestamp 1698175906
transform 1 0 15568 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform 1 0 21952 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _127_
timestamp 1698175906
transform -1 0 19376 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _128_
timestamp 1698175906
transform -1 0 17920 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_
timestamp 1698175906
transform 1 0 14560 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _130_
timestamp 1698175906
transform -1 0 16352 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform 1 0 17584 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _132_
timestamp 1698175906
transform -1 0 16352 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _133_
timestamp 1698175906
transform 1 0 19600 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _134_
timestamp 1698175906
transform -1 0 16352 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _135_
timestamp 1698175906
transform -1 0 15792 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _136_
timestamp 1698175906
transform 1 0 13888 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _137_
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19600 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _139_
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _140_
timestamp 1698175906
transform -1 0 15680 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _141_
timestamp 1698175906
transform 1 0 14224 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _142_
timestamp 1698175906
transform 1 0 13664 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _143_
timestamp 1698175906
transform -1 0 20496 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _144_
timestamp 1698175906
transform -1 0 23184 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _145_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18592 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _146_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18928 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _147_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21392 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _148_
timestamp 1698175906
transform 1 0 18704 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _149_
timestamp 1698175906
transform -1 0 18928 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _150_
timestamp 1698175906
transform -1 0 21056 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _151_
timestamp 1698175906
transform -1 0 20384 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _152_
timestamp 1698175906
transform -1 0 27328 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _153_
timestamp 1698175906
transform -1 0 22064 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _154_
timestamp 1698175906
transform 1 0 24080 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _155_
timestamp 1698175906
transform 1 0 18032 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _156_
timestamp 1698175906
transform 1 0 24864 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _157_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _158_
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _159_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 26656 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _160_
timestamp 1698175906
transform -1 0 28000 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _161_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _162_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21504 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _163_
timestamp 1698175906
transform 1 0 25984 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _164_
timestamp 1698175906
transform -1 0 28112 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _165_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25424 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _166_
timestamp 1698175906
transform -1 0 28448 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _167_
timestamp 1698175906
transform 1 0 22400 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _168_
timestamp 1698175906
transform 1 0 23408 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _169_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _170_
timestamp 1698175906
transform -1 0 24640 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _171_
timestamp 1698175906
transform 1 0 22288 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _172_
timestamp 1698175906
transform 1 0 26208 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _173_
timestamp 1698175906
transform -1 0 15456 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _174_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18816 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _175_
timestamp 1698175906
transform 1 0 14560 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _176_
timestamp 1698175906
transform 1 0 14672 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _177_
timestamp 1698175906
transform 1 0 13328 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _178_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13328 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _179_
timestamp 1698175906
transform 1 0 11536 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _180_
timestamp 1698175906
transform -1 0 19376 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _181_
timestamp 1698175906
transform -1 0 19152 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _182_
timestamp 1698175906
transform 1 0 16352 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _183_
timestamp 1698175906
transform -1 0 16800 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _184_
timestamp 1698175906
transform -1 0 16128 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _185_
timestamp 1698175906
transform 1 0 25984 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _186_
timestamp 1698175906
transform 1 0 25312 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _187_
timestamp 1698175906
transform -1 0 23520 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _188_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _189_
timestamp 1698175906
transform 1 0 21392 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _190_
timestamp 1698175906
transform 1 0 22288 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _191_
timestamp 1698175906
transform -1 0 14560 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _192_
timestamp 1698175906
transform 1 0 12208 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _193_
timestamp 1698175906
transform -1 0 25536 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _194_
timestamp 1698175906
transform -1 0 21952 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _195_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22400 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _196_
timestamp 1698175906
transform -1 0 20944 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _197_
timestamp 1698175906
transform 1 0 19936 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _198_
timestamp 1698175906
transform 1 0 18704 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _199_
timestamp 1698175906
transform 1 0 19152 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _200_
timestamp 1698175906
transform 1 0 17472 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _201_
timestamp 1698175906
transform -1 0 18144 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _202_
timestamp 1698175906
transform 1 0 20720 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _203_
timestamp 1698175906
transform -1 0 24640 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform -1 0 24976 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform 1 0 9744 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform 1 0 9744 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform 1 0 16128 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform 1 0 12880 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform -1 0 15120 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 17136 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 18704 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 25648 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 25536 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 26096 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform -1 0 14672 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform -1 0 12992 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 17360 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 13328 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 21504 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform -1 0 13664 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 22624 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform -1 0 20496 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 15456 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform -1 0 24864 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _231_
timestamp 1698175906
transform 1 0 19712 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _232_
timestamp 1698175906
transform -1 0 21280 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _233_
timestamp 1698175906
transform -1 0 14000 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24192 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 25200 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 13552 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 13216 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 19600 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 15344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 16912 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform -1 0 22400 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 28560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 25872 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 14672 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 12992 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 28560 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 13888 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 26768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 20720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 19600 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 17024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18144 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 20496 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 21728 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698175906
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698175906
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_195 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23184 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_203
timestamp 1698175906
transform 1 0 24080 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_107 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_123
timestamp 1698175906
transform 1 0 15120 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_131
timestamp 1698175906
transform 1 0 16016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_159
timestamp 1698175906
transform 1 0 19152 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_333
timestamp 1698175906
transform 1 0 38640 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_341
timestamp 1698175906
transform 1 0 39536 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_139
timestamp 1698175906
transform 1 0 16912 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_155
timestamp 1698175906
transform 1 0 18704 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_163
timestamp 1698175906
transform 1 0 19600 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_170
timestamp 1698175906
transform 1 0 20384 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_88
timestamp 1698175906
transform 1 0 11200 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_96
timestamp 1698175906
transform 1 0 12096 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_100
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_102
timestamp 1698175906
transform 1 0 12768 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_132
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_178
timestamp 1698175906
transform 1 0 21280 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_115
timestamp 1698175906
transform 1 0 14224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_121
timestamp 1698175906
transform 1 0 14896 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_125
timestamp 1698175906
transform 1 0 15344 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_155
timestamp 1698175906
transform 1 0 18704 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_161
timestamp 1698175906
transform 1 0 19376 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_165
timestamp 1698175906
transform 1 0 19824 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698175906
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_88
timestamp 1698175906
transform 1 0 11200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_119
timestamp 1698175906
transform 1 0 14672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_134
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698175906
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_150
timestamp 1698175906
transform 1 0 18144 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_159
timestamp 1698175906
transform 1 0 19152 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_202
timestamp 1698175906
transform 1 0 23968 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698175906
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_115
timestamp 1698175906
transform 1 0 14224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_127
timestamp 1698175906
transform 1 0 15568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_143
timestamp 1698175906
transform 1 0 17360 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_149
timestamp 1698175906
transform 1 0 18032 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_165
timestamp 1698175906
transform 1 0 19824 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_181
timestamp 1698175906
transform 1 0 21616 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_211
timestamp 1698175906
transform 1 0 24976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_215
timestamp 1698175906
transform 1 0 25424 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_231
timestamp 1698175906
transform 1 0 27216 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_239
timestamp 1698175906
transform 1 0 28112 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 4480 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_106
timestamp 1698175906
transform 1 0 13216 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_114
timestamp 1698175906
transform 1 0 14112 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_134
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698175906
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_158
timestamp 1698175906
transform 1 0 19040 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_166
timestamp 1698175906
transform 1 0 19936 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_168
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_183
timestamp 1698175906
transform 1 0 21840 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_197
timestamp 1698175906
transform 1 0 23408 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_205
timestamp 1698175906
transform 1 0 24304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_241
timestamp 1698175906
transform 1 0 28336 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_245
timestamp 1698175906
transform 1 0 28784 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698175906
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_69
timestamp 1698175906
transform 1 0 9072 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_73
timestamp 1698175906
transform 1 0 9520 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1698175906
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_113
timestamp 1698175906
transform 1 0 14000 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_126
timestamp 1698175906
transform 1 0 15456 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_128
timestamp 1698175906
transform 1 0 15680 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_140
timestamp 1698175906
transform 1 0 17024 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_144
timestamp 1698175906
transform 1 0 17472 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_151
timestamp 1698175906
transform 1 0 18256 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_159
timestamp 1698175906
transform 1 0 19152 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698175906
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_187
timestamp 1698175906
transform 1 0 22288 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_203
timestamp 1698175906
transform 1 0 24080 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_211
timestamp 1698175906
transform 1 0 24976 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_215
timestamp 1698175906
transform 1 0 25424 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_226
timestamp 1698175906
transform 1 0 26656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_232
timestamp 1698175906
transform 1 0 27328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_238
timestamp 1698175906
transform 1 0 28000 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_242
timestamp 1698175906
transform 1 0 28448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 4480 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 8064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_88
timestamp 1698175906
transform 1 0 11200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_90
timestamp 1698175906
transform 1 0 11424 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_95
timestamp 1698175906
transform 1 0 11984 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_115
timestamp 1698175906
transform 1 0 14224 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_131
timestamp 1698175906
transform 1 0 16016 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_150
timestamp 1698175906
transform 1 0 18144 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_154
timestamp 1698175906
transform 1 0 18592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_195
timestamp 1698175906
transform 1 0 23184 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_203
timestamp 1698175906
transform 1 0 24080 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_207
timestamp 1698175906
transform 1 0 24528 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_216
timestamp 1698175906
transform 1 0 25536 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_246
timestamp 1698175906
transform 1 0 28896 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_111
timestamp 1698175906
transform 1 0 13776 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_139
timestamp 1698175906
transform 1 0 16912 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_147
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_151
timestamp 1698175906
transform 1 0 18256 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_194
timestamp 1698175906
transform 1 0 23072 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_210
timestamp 1698175906
transform 1 0 24864 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_218
timestamp 1698175906
transform 1 0 25760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_230
timestamp 1698175906
transform 1 0 27104 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_238
timestamp 1698175906
transform 1 0 28000 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_242
timestamp 1698175906
transform 1 0 28448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_74
timestamp 1698175906
transform 1 0 9632 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_104
timestamp 1698175906
transform 1 0 12992 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_116
timestamp 1698175906
transform 1 0 14336 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_150
timestamp 1698175906
transform 1 0 18144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_154
timestamp 1698175906
transform 1 0 18592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_179
timestamp 1698175906
transform 1 0 21392 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_198
timestamp 1698175906
transform 1 0 23520 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_202
timestamp 1698175906
transform 1 0 23968 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_214
timestamp 1698175906
transform 1 0 25312 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_227
timestamp 1698175906
transform 1 0 26768 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_239
timestamp 1698175906
transform 1 0 28112 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_271
timestamp 1698175906
transform 1 0 31696 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 40320 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_111
timestamp 1698175906
transform 1 0 13776 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698175906
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_185
timestamp 1698175906
transform 1 0 22064 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_208
timestamp 1698175906
transform 1 0 24640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_88
timestamp 1698175906
transform 1 0 11200 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_96
timestamp 1698175906
transform 1 0 12096 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_100
timestamp 1698175906
transform 1 0 12544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_126
timestamp 1698175906
transform 1 0 15456 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_133
timestamp 1698175906
transform 1 0 16240 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_148
timestamp 1698175906
transform 1 0 17920 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698175906
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_216
timestamp 1698175906
transform 1 0 25536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_218
timestamp 1698175906
transform 1 0 25760 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_250
timestamp 1698175906
transform 1 0 29344 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_266
timestamp 1698175906
transform 1 0 31136 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_274
timestamp 1698175906
transform 1 0 32032 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_69
timestamp 1698175906
transform 1 0 9072 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_73
timestamp 1698175906
transform 1 0 9520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_104
timestamp 1698175906
transform 1 0 12992 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_111
timestamp 1698175906
transform 1 0 13776 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_118
timestamp 1698175906
transform 1 0 14560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_122
timestamp 1698175906
transform 1 0 15008 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_129
timestamp 1698175906
transform 1 0 15792 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_137
timestamp 1698175906
transform 1 0 16688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_139
timestamp 1698175906
transform 1 0 16912 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_147
timestamp 1698175906
transform 1 0 17808 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_177
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_181
timestamp 1698175906
transform 1 0 21616 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_232
timestamp 1698175906
transform 1 0 27328 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_236
timestamp 1698175906
transform 1 0 27776 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_242
timestamp 1698175906
transform 1 0 28448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_104
timestamp 1698175906
transform 1 0 12992 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_112
timestamp 1698175906
transform 1 0 13888 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_128
timestamp 1698175906
transform 1 0 15680 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_146
timestamp 1698175906
transform 1 0 17696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_148
timestamp 1698175906
transform 1 0 17920 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_171
timestamp 1698175906
transform 1 0 20496 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_216
timestamp 1698175906
transform 1 0 25536 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_220
timestamp 1698175906
transform 1 0 25984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_232
timestamp 1698175906
transform 1 0 27328 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_264
timestamp 1698175906
transform 1 0 30912 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 40320 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_69
timestamp 1698175906
transform 1 0 9072 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_85
timestamp 1698175906
transform 1 0 10864 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_93
timestamp 1698175906
transform 1 0 11760 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_118
timestamp 1698175906
transform 1 0 14560 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_134
timestamp 1698175906
transform 1 0 16352 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_138
timestamp 1698175906
transform 1 0 16800 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_170
timestamp 1698175906
transform 1 0 20384 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_209
timestamp 1698175906
transform 1 0 24752 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_213
timestamp 1698175906
transform 1 0 25200 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_222
timestamp 1698175906
transform 1 0 26208 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_238
timestamp 1698175906
transform 1 0 28000 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698175906
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 4480 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 8064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_80
timestamp 1698175906
transform 1 0 10304 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_110
timestamp 1698175906
transform 1 0 13664 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_114
timestamp 1698175906
transform 1 0 14112 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_122
timestamp 1698175906
transform 1 0 15008 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_126
timestamp 1698175906
transform 1 0 15456 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_128
timestamp 1698175906
transform 1 0 15680 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_148
timestamp 1698175906
transform 1 0 17920 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_164
timestamp 1698175906
transform 1 0 19712 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_174
timestamp 1698175906
transform 1 0 20832 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_184
timestamp 1698175906
transform 1 0 21952 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_199
timestamp 1698175906
transform 1 0 23632 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_207
timestamp 1698175906
transform 1 0 24528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698175906
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_241
timestamp 1698175906
transform 1 0 28336 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_245
timestamp 1698175906
transform 1 0 28784 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698175906
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_132
timestamp 1698175906
transform 1 0 16128 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_148
timestamp 1698175906
transform 1 0 17920 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_156
timestamp 1698175906
transform 1 0 18816 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_158
timestamp 1698175906
transform 1 0 19040 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_166
timestamp 1698175906
transform 1 0 19936 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_219
timestamp 1698175906
transform 1 0 25872 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_225
timestamp 1698175906
transform 1 0 26544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_229
timestamp 1698175906
transform 1 0 26992 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 4480 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_104
timestamp 1698175906
transform 1 0 12992 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_106
timestamp 1698175906
transform 1 0 13216 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_136
timestamp 1698175906
transform 1 0 16576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_171
timestamp 1698175906
transform 1 0 20496 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_175
timestamp 1698175906
transform 1 0 20944 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698175906
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_216
timestamp 1698175906
transform 1 0 25536 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_139
timestamp 1698175906
transform 1 0 16912 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_160
timestamp 1698175906
transform 1 0 19264 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_168
timestamp 1698175906
transform 1 0 20160 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_172
timestamp 1698175906
transform 1 0 20608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698175906
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_185
timestamp 1698175906
transform 1 0 22064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_192
timestamp 1698175906
transform 1 0 22848 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_198
timestamp 1698175906
transform 1 0 23520 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_230
timestamp 1698175906
transform 1 0 27104 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698175906
transform 1 0 28000 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_88
timestamp 1698175906
transform 1 0 11200 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_92
timestamp 1698175906
transform 1 0 11648 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_123
timestamp 1698175906
transform 1 0 15120 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_127
timestamp 1698175906
transform 1 0 15568 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_135
timestamp 1698175906
transform 1 0 16464 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698175906
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_148
timestamp 1698175906
transform 1 0 17920 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_161
timestamp 1698175906
transform 1 0 19376 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_170
timestamp 1698175906
transform 1 0 20384 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_176
timestamp 1698175906
transform 1 0 21056 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_216
timestamp 1698175906
transform 1 0 25536 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_123
timestamp 1698175906
transform 1 0 15120 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_131
timestamp 1698175906
transform 1 0 16016 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_161
timestamp 1698175906
transform 1 0 19376 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_165
timestamp 1698175906
transform 1 0 19824 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_173
timestamp 1698175906
transform 1 0 20720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_150
timestamp 1698175906
transform 1 0 18144 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_154
timestamp 1698175906
transform 1 0 18592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_184
timestamp 1698175906
transform 1 0 21952 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_188
timestamp 1698175906
transform 1 0 22400 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_204
timestamp 1698175906
transform 1 0 24192 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_208
timestamp 1698175906
transform 1 0 24640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_123
timestamp 1698175906
transform 1 0 15120 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_131
timestamp 1698175906
transform 1 0 16016 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_159
timestamp 1698175906
transform 1 0 19152 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_195
timestamp 1698175906
transform 1 0 23184 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698175906
transform 1 0 24080 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 25536 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_243
timestamp 1698175906
transform 1 0 28560 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698175906
transform 1 0 32144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_244
timestamp 1698175906
transform 1 0 28672 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_260
timestamp 1698175906
transform 1 0 30464 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_268
timestamp 1698175906
transform 1 0 31360 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita57_24 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 28672 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita57_25
timestamp 1698175906
transform 1 0 39984 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita57_26
timestamp 1698175906
transform -1 0 27776 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform -1 0 4480 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 20944 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 4480 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 20384 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 4480 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 25648 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 21280 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 37520 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 20272 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 4480 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 20272 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 16240 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 20272 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 17360 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 4480 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 16240 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 26880 41200 26992 42000 0 FreeSans 448 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 19488 41200 19600 42000 0 FreeSans 448 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 41200 21504 42000 21616 0 FreeSans 448 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 41200 10752 42000 10864 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 26208 41200 26320 42000 0 FreeSans 448 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 41200 16800 42000 16912 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 25536 41200 25648 42000 0 FreeSans 448 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 21504 41200 21616 42000 0 FreeSans 448 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 41200 24864 42000 24976 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 24192 41200 24304 42000 0 FreeSans 448 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 20160 41200 20272 42000 0 FreeSans 448 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 18816 41200 18928 42000 0 FreeSans 448 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 16128 41200 16240 42000 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 27048 21728 27048 21728 0 _000_
rlabel metal2 13720 15624 13720 15624 0 _001_
rlabel metal2 12040 17976 12040 17976 0 _002_
rlabel metal2 18312 14476 18312 14476 0 _003_
rlabel metal2 15848 25928 15848 25928 0 _004_
rlabel metal2 25592 24304 25592 24304 0 _005_
rlabel metal2 22568 27496 22568 27496 0 _006_
rlabel metal2 12488 24360 12488 24360 0 _007_
rlabel metal2 23352 25144 23352 25144 0 _008_
rlabel metal2 19544 25872 19544 25872 0 _009_
rlabel metal3 17136 15176 17136 15176 0 _010_
rlabel metal2 23912 22344 23912 22344 0 _011_
rlabel metal3 19880 22568 19880 22568 0 _012_
rlabel metal2 24192 16184 24192 16184 0 _013_
rlabel metal2 10696 22736 10696 22736 0 _014_
rlabel metal3 12376 19880 12376 19880 0 _015_
rlabel metal2 17416 28280 17416 28280 0 _016_
rlabel metal2 13832 14504 13832 14504 0 _017_
rlabel metal2 14504 26656 14504 26656 0 _018_
rlabel metal2 18200 23520 18200 23520 0 _019_
rlabel metal2 19768 28056 19768 28056 0 _020_
rlabel metal2 26040 17360 26040 17360 0 _021_
rlabel metal2 26600 18592 26600 18592 0 _022_
rlabel metal2 26432 20216 26432 20216 0 _023_
rlabel metal3 22232 20104 22232 20104 0 _024_
rlabel metal2 26264 20272 26264 20272 0 _025_
rlabel metal2 25032 21280 25032 21280 0 _026_
rlabel metal2 26824 23352 26824 23352 0 _027_
rlabel metal3 23520 17416 23520 17416 0 _028_
rlabel metal2 25704 17920 25704 17920 0 _029_
rlabel metal2 26712 18312 26712 18312 0 _030_
rlabel metal2 20664 21840 20664 21840 0 _031_
rlabel metal3 24416 19880 24416 19880 0 _032_
rlabel metal3 27160 19992 27160 19992 0 _033_
rlabel metal2 28168 22904 28168 22904 0 _034_
rlabel metal2 21448 18928 21448 18928 0 _035_
rlabel metal2 22456 24808 22456 24808 0 _036_
rlabel metal2 22792 20496 22792 20496 0 _037_
rlabel metal2 23240 20720 23240 20720 0 _038_
rlabel metal2 22568 22120 22568 22120 0 _039_
rlabel metal2 15064 17192 15064 17192 0 _040_
rlabel metal2 18760 16744 18760 16744 0 _041_
rlabel metal2 14840 16408 14840 16408 0 _042_
rlabel metal3 13272 18312 13272 18312 0 _043_
rlabel metal2 11704 18536 11704 18536 0 _044_
rlabel metal2 19096 15008 19096 15008 0 _045_
rlabel metal3 18480 24696 18480 24696 0 _046_
rlabel metal2 16016 24584 16016 24584 0 _047_
rlabel metal2 26264 23912 26264 23912 0 _048_
rlabel metal2 22568 26908 22568 26908 0 _049_
rlabel metal2 24024 21280 24024 21280 0 _050_
rlabel metal2 21672 25592 21672 25592 0 _051_
rlabel metal2 13832 23968 13832 23968 0 _052_
rlabel metal2 23464 24976 23464 24976 0 _053_
rlabel metal3 22344 24584 22344 24584 0 _054_
rlabel metal2 20888 21168 20888 21168 0 _055_
rlabel metal3 19880 24920 19880 24920 0 _056_
rlabel metal2 19208 26152 19208 26152 0 _057_
rlabel metal2 17976 15624 17976 15624 0 _058_
rlabel metal2 24360 21840 24360 21840 0 _059_
rlabel metal2 23464 16072 23464 16072 0 _060_
rlabel metal2 14056 22792 14056 22792 0 _061_
rlabel metal2 15288 22008 15288 22008 0 _062_
rlabel metal2 16520 21896 16520 21896 0 _063_
rlabel metal3 17808 23128 17808 23128 0 _064_
rlabel metal2 19208 19376 19208 19376 0 _065_
rlabel metal2 21224 19208 21224 19208 0 _066_
rlabel metal3 17696 19432 17696 19432 0 _067_
rlabel metal2 13944 19824 13944 19824 0 _068_
rlabel metal2 14392 20860 14392 20860 0 _069_
rlabel metal2 13496 20608 13496 20608 0 _070_
rlabel metal3 22344 23240 22344 23240 0 _071_
rlabel metal2 17584 22568 17584 22568 0 _072_
rlabel metal2 17416 19600 17416 19600 0 _073_
rlabel metal2 14728 17360 14728 17360 0 _074_
rlabel metal2 14784 20776 14784 20776 0 _075_
rlabel metal3 14644 20104 14644 20104 0 _076_
rlabel metal2 18368 22120 18368 22120 0 _077_
rlabel metal2 13720 19712 13720 19712 0 _078_
rlabel metal2 17416 23352 17416 23352 0 _079_
rlabel metal2 23184 24584 23184 24584 0 _080_
rlabel metal3 18312 27832 18312 27832 0 _081_
rlabel metal2 15064 18984 15064 18984 0 _082_
rlabel metal2 15848 17136 15848 17136 0 _083_
rlabel metal2 18088 17584 18088 17584 0 _084_
rlabel metal2 15736 15288 15736 15288 0 _085_
rlabel metal2 20328 23016 20328 23016 0 _086_
rlabel metal2 15400 16352 15400 16352 0 _087_
rlabel metal2 14616 25032 14616 25032 0 _088_
rlabel metal3 18928 19992 18928 19992 0 _089_
rlabel metal2 14392 25312 14392 25312 0 _090_
rlabel metal2 13720 24192 13720 24192 0 _091_
rlabel metal2 15064 25480 15064 25480 0 _092_
rlabel metal2 14840 22120 14840 22120 0 _093_
rlabel metal2 19824 23352 19824 23352 0 _094_
rlabel metal2 20272 19208 20272 19208 0 _095_
rlabel metal2 19320 22848 19320 22848 0 _096_
rlabel metal2 18536 23240 18536 23240 0 _097_
rlabel metal2 19096 19376 19096 19376 0 _098_
rlabel metal2 18200 22064 18200 22064 0 _099_
rlabel metal2 20384 27832 20384 27832 0 _100_
rlabel metal2 26264 17472 26264 17472 0 _101_
rlabel metal3 2478 28280 2478 28280 0 clk
rlabel metal2 21840 21672 21840 21672 0 clknet_0_clk
rlabel metal2 13608 22008 13608 22008 0 clknet_1_0__leaf_clk
rlabel metal3 22288 15288 22288 15288 0 clknet_1_1__leaf_clk
rlabel metal2 22792 16016 22792 16016 0 dut57.count\[0\]
rlabel metal2 23016 17640 23016 17640 0 dut57.count\[1\]
rlabel metal2 12824 22792 12824 22792 0 dut57.count\[2\]
rlabel metal3 13440 19320 13440 19320 0 dut57.count\[3\]
rlabel metal3 28280 20888 28280 20888 0 net1
rlabel metal2 27832 18032 27832 18032 0 net10
rlabel metal2 25760 25592 25760 25592 0 net11
rlabel metal2 21784 33656 21784 33656 0 net12
rlabel metal2 28168 25032 28168 25032 0 net13
rlabel metal2 24584 32872 24584 32872 0 net14
rlabel metal2 20328 24024 20328 24024 0 net15
rlabel metal2 12040 26544 12040 26544 0 net16
rlabel metal2 19208 32984 19208 32984 0 net17
rlabel metal2 16408 25536 16408 25536 0 net18
rlabel metal2 20440 6356 20440 6356 0 net19
rlabel metal3 17640 27720 17640 27720 0 net2
rlabel metal3 18088 14616 18088 14616 0 net20
rlabel metal2 13496 17584 13496 17584 0 net21
rlabel metal2 16408 6748 16408 6748 0 net22
rlabel metal2 37688 22680 37688 22680 0 net23
rlabel metal2 28392 38248 28392 38248 0 net24
rlabel metal2 40264 10976 40264 10976 0 net25
rlabel metal2 26264 39578 26264 39578 0 net26
rlabel metal2 11592 16016 11592 16016 0 net3
rlabel metal2 28280 21840 28280 21840 0 net4
rlabel metal2 21000 12712 21000 12712 0 net5
rlabel metal2 9912 18088 9912 18088 0 net6
rlabel metal3 20216 14000 20216 14000 0 net7
rlabel metal3 6356 24696 6356 24696 0 net8
rlabel metal2 28168 17192 28168 17192 0 net9
rlabel metal3 40642 20888 40642 20888 0 segm[10]
rlabel metal2 19544 39746 19544 39746 0 segm[11]
rlabel metal3 1358 16184 1358 16184 0 segm[12]
rlabel metal2 40040 21504 40040 21504 0 segm[13]
rlabel metal2 20888 2198 20888 2198 0 segm[1]
rlabel metal3 1358 18200 1358 18200 0 segm[2]
rlabel metal2 19544 2030 19544 2030 0 segm[4]
rlabel metal3 1358 24248 1358 24248 0 segm[6]
rlabel metal2 40040 17304 40040 17304 0 segm[7]
rlabel metal3 40642 18200 40642 18200 0 segm[8]
rlabel metal2 26824 37968 26824 37968 0 segm[9]
rlabel metal3 22008 38248 22008 38248 0 sel[0]
rlabel metal2 40040 25256 40040 25256 0 sel[10]
rlabel metal3 24920 38248 24920 38248 0 sel[11]
rlabel metal3 20832 37464 20832 37464 0 sel[1]
rlabel metal3 1358 25592 1358 25592 0 sel[2]
rlabel metal2 18872 39942 18872 39942 0 sel[3]
rlabel metal3 16800 36680 16800 36680 0 sel[4]
rlabel metal2 20216 2422 20216 2422 0 sel[5]
rlabel metal2 18200 2422 18200 2422 0 sel[6]
rlabel metal3 1358 17528 1358 17528 0 sel[7]
rlabel metal2 16184 2982 16184 2982 0 sel[8]
rlabel metal2 40040 22344 40040 22344 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
