magic
tech gf180mcuD
magscale 1 5
timestamp 1699641115
<< obsm1 >>
rect 672 1538 20328 19238
<< metal2 >>
rect 7728 20600 7784 21000
rect 9408 20600 9464 21000
rect 9744 20600 9800 21000
rect 10752 20600 10808 21000
rect 11088 20600 11144 21000
rect 12432 20600 12488 21000
rect 12768 20600 12824 21000
rect 15120 20600 15176 21000
rect 9408 0 9464 400
rect 9744 0 9800 400
rect 10080 0 10136 400
rect 11424 0 11480 400
rect 11760 0 11816 400
rect 17808 0 17864 400
<< obsm2 >>
rect 966 20570 7698 20600
rect 7814 20570 9378 20600
rect 9494 20570 9714 20600
rect 9830 20570 10722 20600
rect 10838 20570 11058 20600
rect 11174 20570 12402 20600
rect 12518 20570 12738 20600
rect 12854 20570 15090 20600
rect 15206 20570 20034 20600
rect 966 430 20034 20570
rect 966 400 9378 430
rect 9494 400 9714 430
rect 9830 400 10050 430
rect 10166 400 11394 430
rect 11510 400 11730 430
rect 11846 400 17778 430
rect 17894 400 20034 430
<< metal3 >>
rect 0 13776 400 13832
rect 0 13104 400 13160
rect 20600 12096 21000 12152
rect 20600 11760 21000 11816
rect 20600 11424 21000 11480
rect 20600 11088 21000 11144
rect 20600 10416 21000 10472
rect 20600 9744 21000 9800
rect 20600 9408 21000 9464
rect 0 9072 400 9128
rect 0 8064 400 8120
rect 20600 8064 21000 8120
rect 20600 7728 21000 7784
<< obsm3 >>
rect 400 13862 20600 19306
rect 430 13746 20600 13862
rect 400 13190 20600 13746
rect 430 13074 20600 13190
rect 400 12182 20600 13074
rect 400 12066 20570 12182
rect 400 11846 20600 12066
rect 400 11730 20570 11846
rect 400 11510 20600 11730
rect 400 11394 20570 11510
rect 400 11174 20600 11394
rect 400 11058 20570 11174
rect 400 10502 20600 11058
rect 400 10386 20570 10502
rect 400 9830 20600 10386
rect 400 9714 20570 9830
rect 400 9494 20600 9714
rect 400 9378 20570 9494
rect 400 9158 20600 9378
rect 430 9042 20600 9158
rect 400 8150 20600 9042
rect 430 8034 20570 8150
rect 400 7814 20600 8034
rect 400 7698 20570 7814
rect 400 1554 20600 7698
<< metal4 >>
rect 2224 1538 2384 19238
rect 9904 1538 10064 19238
rect 17584 1538 17744 19238
<< obsm4 >>
rect 13454 8241 13482 8559
<< labels >>
rlabel metal3 s 0 13776 400 13832 6 clk
port 1 nsew signal input
rlabel metal2 s 15120 20600 15176 21000 6 segm[0]
port 2 nsew signal output
rlabel metal3 s 20600 10416 21000 10472 6 segm[10]
port 3 nsew signal output
rlabel metal3 s 20600 11760 21000 11816 6 segm[11]
port 4 nsew signal output
rlabel metal3 s 20600 7728 21000 7784 6 segm[12]
port 5 nsew signal output
rlabel metal2 s 11424 0 11480 400 6 segm[13]
port 6 nsew signal output
rlabel metal2 s 11088 20600 11144 21000 6 segm[1]
port 7 nsew signal output
rlabel metal2 s 9744 0 9800 400 6 segm[2]
port 8 nsew signal output
rlabel metal2 s 9408 0 9464 400 6 segm[3]
port 9 nsew signal output
rlabel metal2 s 10752 20600 10808 21000 6 segm[4]
port 10 nsew signal output
rlabel metal2 s 17808 0 17864 400 6 segm[5]
port 11 nsew signal output
rlabel metal3 s 20600 8064 21000 8120 6 segm[6]
port 12 nsew signal output
rlabel metal3 s 20600 9744 21000 9800 6 segm[7]
port 13 nsew signal output
rlabel metal2 s 9408 20600 9464 21000 6 segm[8]
port 14 nsew signal output
rlabel metal3 s 20600 9408 21000 9464 6 segm[9]
port 15 nsew signal output
rlabel metal2 s 10080 0 10136 400 6 sel[0]
port 16 nsew signal output
rlabel metal2 s 12768 20600 12824 21000 6 sel[10]
port 17 nsew signal output
rlabel metal2 s 12432 20600 12488 21000 6 sel[11]
port 18 nsew signal output
rlabel metal2 s 7728 20600 7784 21000 6 sel[1]
port 19 nsew signal output
rlabel metal3 s 20600 12096 21000 12152 6 sel[2]
port 20 nsew signal output
rlabel metal3 s 0 13104 400 13160 6 sel[3]
port 21 nsew signal output
rlabel metal3 s 0 9072 400 9128 6 sel[4]
port 22 nsew signal output
rlabel metal3 s 20600 11424 21000 11480 6 sel[5]
port 23 nsew signal output
rlabel metal2 s 9744 20600 9800 21000 6 sel[6]
port 24 nsew signal output
rlabel metal3 s 0 8064 400 8120 6 sel[7]
port 25 nsew signal output
rlabel metal3 s 20600 11088 21000 11144 6 sel[8]
port 26 nsew signal output
rlabel metal2 s 11760 0 11816 400 6 sel[9]
port 27 nsew signal output
rlabel metal4 s 2224 1538 2384 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 19238 6 vss
port 29 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 21000 21000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 486930
string GDS_FILE /home/urielcho/Proyectos_caravel/ITA23_GFMPW1b/openlane/ita1/runs/23_11_10_12_29/results/signoff/ita1.magic.gds
string GDS_START 168908
<< end >>

