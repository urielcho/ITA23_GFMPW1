magic
tech gf180mcuD
magscale 1 5
timestamp 1699711247
<< obsm1 >>
rect 672 1538 31304 268617
<< metal2 >>
rect 560 269800 616 270200
rect 1120 269800 1176 270200
rect 1680 269800 1736 270200
rect 2240 269800 2296 270200
rect 2800 269800 2856 270200
rect 3360 269800 3416 270200
rect 3920 269800 3976 270200
rect 4480 269800 4536 270200
rect 5040 269800 5096 270200
rect 5600 269800 5656 270200
rect 6160 269800 6216 270200
rect 6720 269800 6776 270200
rect 7280 269800 7336 270200
rect 7840 269800 7896 270200
rect 8400 269800 8456 270200
rect 8960 269800 9016 270200
rect 9520 269800 9576 270200
rect 10080 269800 10136 270200
rect 10640 269800 10696 270200
rect 11200 269800 11256 270200
rect 11760 269800 11816 270200
rect 12320 269800 12376 270200
rect 12880 269800 12936 270200
rect 13440 269800 13496 270200
rect 14000 269800 14056 270200
rect 14560 269800 14616 270200
rect 15120 269800 15176 270200
rect 15680 269800 15736 270200
rect 16240 269800 16296 270200
rect 16800 269800 16856 270200
rect 17360 269800 17416 270200
rect 17920 269800 17976 270200
rect 18480 269800 18536 270200
rect 19040 269800 19096 270200
rect 19600 269800 19656 270200
rect 20160 269800 20216 270200
rect 20720 269800 20776 270200
rect 21280 269800 21336 270200
rect 21840 269800 21896 270200
rect 22400 269800 22456 270200
rect 22960 269800 23016 270200
rect 23520 269800 23576 270200
rect 24080 269800 24136 270200
rect 24640 269800 24696 270200
rect 25200 269800 25256 270200
rect 25760 269800 25816 270200
rect 26320 269800 26376 270200
rect 26880 269800 26936 270200
rect 27440 269800 27496 270200
rect 28000 269800 28056 270200
rect 28560 269800 28616 270200
rect 29120 269800 29176 270200
rect 29680 269800 29736 270200
rect 30240 269800 30296 270200
rect 30800 269800 30856 270200
rect 31360 269800 31416 270200
rect 1008 0 1064 400
rect 3136 0 3192 400
rect 5264 0 5320 400
rect 7392 0 7448 400
rect 9520 0 9576 400
rect 11648 0 11704 400
rect 13776 0 13832 400
rect 15904 0 15960 400
rect 18032 0 18088 400
rect 20160 0 20216 400
rect 22288 0 22344 400
rect 24416 0 24472 400
rect 26544 0 26600 400
rect 28672 0 28728 400
rect 30800 0 30856 400
<< obsm2 >>
rect 238 269770 530 269850
rect 646 269770 1090 269850
rect 1206 269770 1650 269850
rect 1766 269770 2210 269850
rect 2326 269770 2770 269850
rect 2886 269770 3330 269850
rect 3446 269770 3890 269850
rect 4006 269770 4450 269850
rect 4566 269770 5010 269850
rect 5126 269770 5570 269850
rect 5686 269770 6130 269850
rect 6246 269770 6690 269850
rect 6806 269770 7250 269850
rect 7366 269770 7810 269850
rect 7926 269770 8370 269850
rect 8486 269770 8930 269850
rect 9046 269770 9490 269850
rect 9606 269770 10050 269850
rect 10166 269770 10610 269850
rect 10726 269770 11170 269850
rect 11286 269770 11730 269850
rect 11846 269770 12290 269850
rect 12406 269770 12850 269850
rect 12966 269770 13410 269850
rect 13526 269770 13970 269850
rect 14086 269770 14530 269850
rect 14646 269770 15090 269850
rect 15206 269770 15650 269850
rect 15766 269770 16210 269850
rect 16326 269770 16770 269850
rect 16886 269770 17330 269850
rect 17446 269770 17890 269850
rect 18006 269770 18450 269850
rect 18566 269770 19010 269850
rect 19126 269770 19570 269850
rect 19686 269770 20130 269850
rect 20246 269770 20690 269850
rect 20806 269770 21250 269850
rect 21366 269770 21810 269850
rect 21926 269770 22370 269850
rect 22486 269770 22930 269850
rect 23046 269770 23490 269850
rect 23606 269770 24050 269850
rect 24166 269770 24610 269850
rect 24726 269770 25170 269850
rect 25286 269770 25730 269850
rect 25846 269770 26290 269850
rect 26406 269770 26850 269850
rect 26966 269770 27410 269850
rect 27526 269770 27970 269850
rect 28086 269770 28530 269850
rect 28646 269770 29090 269850
rect 29206 269770 29650 269850
rect 29766 269770 30210 269850
rect 30326 269770 30770 269850
rect 30886 269770 31330 269850
rect 31446 269770 31794 269850
rect 238 430 31794 269770
rect 238 350 978 430
rect 1094 350 3106 430
rect 3222 350 5234 430
rect 5350 350 7362 430
rect 7478 350 9490 430
rect 9606 350 11618 430
rect 11734 350 13746 430
rect 13862 350 15874 430
rect 15990 350 18002 430
rect 18118 350 20130 430
rect 20246 350 22258 430
rect 22374 350 24386 430
rect 24502 350 26514 430
rect 26630 350 28642 430
rect 28758 350 30770 430
rect 30886 350 31794 430
<< metal3 >>
rect 0 251160 400 251216
rect 31600 251160 32000 251216
rect 0 250880 400 250936
rect 31600 250880 32000 250936
rect 0 250600 400 250656
rect 31600 250600 32000 250656
rect 0 250320 400 250376
rect 31600 250320 32000 250376
rect 0 250040 400 250096
rect 31600 250040 32000 250096
rect 0 249760 400 249816
rect 31600 249760 32000 249816
rect 0 249480 400 249536
rect 31600 249480 32000 249536
rect 0 249200 400 249256
rect 31600 249200 32000 249256
rect 0 248920 400 248976
rect 31600 248920 32000 248976
rect 0 248640 400 248696
rect 31600 248640 32000 248696
rect 0 248360 400 248416
rect 31600 248360 32000 248416
rect 0 248080 400 248136
rect 31600 248080 32000 248136
rect 0 247800 400 247856
rect 31600 247800 32000 247856
rect 0 247520 400 247576
rect 31600 247520 32000 247576
rect 0 247240 400 247296
rect 31600 247240 32000 247296
rect 0 246960 400 247016
rect 31600 246960 32000 247016
rect 0 246680 400 246736
rect 31600 246680 32000 246736
rect 0 246400 400 246456
rect 31600 246400 32000 246456
rect 0 246120 400 246176
rect 31600 246120 32000 246176
rect 0 245840 400 245896
rect 31600 245840 32000 245896
rect 0 245560 400 245616
rect 31600 245560 32000 245616
rect 0 245280 400 245336
rect 31600 245280 32000 245336
rect 0 245000 400 245056
rect 31600 245000 32000 245056
rect 0 244720 400 244776
rect 31600 244720 32000 244776
rect 0 244440 400 244496
rect 31600 244440 32000 244496
rect 0 244160 400 244216
rect 31600 244160 32000 244216
rect 0 243880 400 243936
rect 31600 243880 32000 243936
rect 0 243600 400 243656
rect 31600 243600 32000 243656
rect 0 243320 400 243376
rect 31600 243320 32000 243376
rect 0 243040 400 243096
rect 31600 243040 32000 243096
rect 0 242760 400 242816
rect 31600 242760 32000 242816
rect 0 242480 400 242536
rect 31600 242480 32000 242536
rect 0 242200 400 242256
rect 31600 242200 32000 242256
rect 0 241920 400 241976
rect 31600 241920 32000 241976
rect 0 241640 400 241696
rect 31600 241640 32000 241696
rect 0 241360 400 241416
rect 31600 241360 32000 241416
rect 0 241080 400 241136
rect 31600 241080 32000 241136
rect 0 240800 400 240856
rect 31600 240800 32000 240856
rect 0 240520 400 240576
rect 31600 240520 32000 240576
rect 0 240240 400 240296
rect 31600 240240 32000 240296
rect 0 239960 400 240016
rect 31600 239960 32000 240016
rect 0 239680 400 239736
rect 31600 239680 32000 239736
rect 0 239400 400 239456
rect 31600 239400 32000 239456
rect 0 239120 400 239176
rect 31600 239120 32000 239176
rect 0 238840 400 238896
rect 31600 238840 32000 238896
rect 0 238560 400 238616
rect 31600 238560 32000 238616
rect 0 238280 400 238336
rect 31600 238280 32000 238336
rect 0 238000 400 238056
rect 31600 238000 32000 238056
rect 0 237720 400 237776
rect 31600 237720 32000 237776
rect 0 237440 400 237496
rect 31600 237440 32000 237496
rect 0 237160 400 237216
rect 31600 237160 32000 237216
rect 0 236880 400 236936
rect 31600 236880 32000 236936
rect 0 236600 400 236656
rect 31600 236600 32000 236656
rect 0 236320 400 236376
rect 31600 236320 32000 236376
rect 0 236040 400 236096
rect 31600 236040 32000 236096
rect 0 235760 400 235816
rect 31600 235760 32000 235816
rect 0 235480 400 235536
rect 31600 235480 32000 235536
rect 0 235200 400 235256
rect 31600 235200 32000 235256
rect 0 234920 400 234976
rect 31600 234920 32000 234976
rect 0 234640 400 234696
rect 31600 234640 32000 234696
rect 0 234360 400 234416
rect 31600 234360 32000 234416
rect 0 234080 400 234136
rect 31600 234080 32000 234136
rect 0 233800 400 233856
rect 31600 233800 32000 233856
rect 0 233520 400 233576
rect 31600 233520 32000 233576
rect 0 233240 400 233296
rect 31600 233240 32000 233296
rect 0 232960 400 233016
rect 31600 232960 32000 233016
rect 0 232680 400 232736
rect 31600 232680 32000 232736
rect 0 232400 400 232456
rect 31600 232400 32000 232456
rect 0 232120 400 232176
rect 31600 232120 32000 232176
rect 0 231840 400 231896
rect 31600 231840 32000 231896
rect 0 231560 400 231616
rect 31600 231560 32000 231616
rect 0 231280 400 231336
rect 31600 231280 32000 231336
rect 0 231000 400 231056
rect 31600 231000 32000 231056
rect 0 230720 400 230776
rect 31600 230720 32000 230776
rect 0 230440 400 230496
rect 31600 230440 32000 230496
rect 0 230160 400 230216
rect 31600 230160 32000 230216
rect 0 229880 400 229936
rect 31600 229880 32000 229936
rect 0 229600 400 229656
rect 31600 229600 32000 229656
rect 0 229320 400 229376
rect 31600 229320 32000 229376
rect 0 229040 400 229096
rect 31600 229040 32000 229096
rect 0 228760 400 228816
rect 31600 228760 32000 228816
rect 0 228480 400 228536
rect 31600 228480 32000 228536
rect 0 228200 400 228256
rect 31600 228200 32000 228256
rect 0 227920 400 227976
rect 31600 227920 32000 227976
rect 0 227640 400 227696
rect 31600 227640 32000 227696
rect 0 227360 400 227416
rect 31600 227360 32000 227416
rect 0 227080 400 227136
rect 31600 227080 32000 227136
rect 0 226800 400 226856
rect 31600 226800 32000 226856
rect 0 226520 400 226576
rect 31600 226520 32000 226576
rect 0 226240 400 226296
rect 31600 226240 32000 226296
rect 0 225960 400 226016
rect 31600 225960 32000 226016
rect 0 225680 400 225736
rect 31600 225680 32000 225736
rect 0 225400 400 225456
rect 31600 225400 32000 225456
rect 0 225120 400 225176
rect 31600 225120 32000 225176
rect 0 224840 400 224896
rect 31600 224840 32000 224896
rect 0 224560 400 224616
rect 31600 224560 32000 224616
rect 0 224280 400 224336
rect 31600 224280 32000 224336
rect 0 224000 400 224056
rect 31600 224000 32000 224056
rect 0 223720 400 223776
rect 31600 223720 32000 223776
rect 0 223440 400 223496
rect 31600 223440 32000 223496
rect 0 223160 400 223216
rect 31600 223160 32000 223216
rect 0 222880 400 222936
rect 31600 222880 32000 222936
rect 0 222600 400 222656
rect 31600 222600 32000 222656
rect 0 222320 400 222376
rect 31600 222320 32000 222376
rect 0 222040 400 222096
rect 31600 222040 32000 222096
rect 0 221760 400 221816
rect 31600 221760 32000 221816
rect 0 221480 400 221536
rect 31600 221480 32000 221536
rect 0 221200 400 221256
rect 31600 221200 32000 221256
rect 0 220920 400 220976
rect 31600 220920 32000 220976
rect 0 220640 400 220696
rect 31600 220640 32000 220696
rect 0 220360 400 220416
rect 31600 220360 32000 220416
rect 0 220080 400 220136
rect 31600 220080 32000 220136
rect 0 219800 400 219856
rect 31600 219800 32000 219856
rect 0 219520 400 219576
rect 31600 219520 32000 219576
rect 0 219240 400 219296
rect 31600 219240 32000 219296
rect 0 218960 400 219016
rect 31600 218960 32000 219016
rect 0 218680 400 218736
rect 31600 218680 32000 218736
rect 0 218400 400 218456
rect 31600 218400 32000 218456
rect 0 218120 400 218176
rect 31600 218120 32000 218176
rect 0 217840 400 217896
rect 31600 217840 32000 217896
rect 0 217560 400 217616
rect 31600 217560 32000 217616
rect 0 217280 400 217336
rect 31600 217280 32000 217336
rect 0 217000 400 217056
rect 31600 217000 32000 217056
rect 0 216720 400 216776
rect 31600 216720 32000 216776
rect 0 216440 400 216496
rect 31600 216440 32000 216496
rect 0 216160 400 216216
rect 31600 216160 32000 216216
rect 0 215880 400 215936
rect 31600 215880 32000 215936
rect 0 215600 400 215656
rect 31600 215600 32000 215656
rect 0 215320 400 215376
rect 31600 215320 32000 215376
rect 0 215040 400 215096
rect 31600 215040 32000 215096
rect 0 214760 400 214816
rect 31600 214760 32000 214816
rect 0 214480 400 214536
rect 31600 214480 32000 214536
rect 0 214200 400 214256
rect 31600 214200 32000 214256
rect 0 213920 400 213976
rect 31600 213920 32000 213976
rect 0 213640 400 213696
rect 31600 213640 32000 213696
rect 0 213360 400 213416
rect 31600 213360 32000 213416
rect 0 213080 400 213136
rect 31600 213080 32000 213136
rect 0 212800 400 212856
rect 31600 212800 32000 212856
rect 0 212520 400 212576
rect 31600 212520 32000 212576
rect 0 212240 400 212296
rect 31600 212240 32000 212296
rect 0 211960 400 212016
rect 31600 211960 32000 212016
rect 0 211680 400 211736
rect 31600 211680 32000 211736
rect 0 211400 400 211456
rect 31600 211400 32000 211456
rect 0 211120 400 211176
rect 31600 211120 32000 211176
rect 0 210840 400 210896
rect 31600 210840 32000 210896
rect 0 210560 400 210616
rect 31600 210560 32000 210616
rect 0 210280 400 210336
rect 31600 210280 32000 210336
rect 0 210000 400 210056
rect 31600 210000 32000 210056
rect 0 209720 400 209776
rect 31600 209720 32000 209776
rect 0 209440 400 209496
rect 31600 209440 32000 209496
rect 0 209160 400 209216
rect 31600 209160 32000 209216
rect 0 208880 400 208936
rect 31600 208880 32000 208936
rect 0 208600 400 208656
rect 31600 208600 32000 208656
rect 0 208320 400 208376
rect 31600 208320 32000 208376
rect 0 208040 400 208096
rect 31600 208040 32000 208096
rect 0 207760 400 207816
rect 31600 207760 32000 207816
rect 0 207480 400 207536
rect 31600 207480 32000 207536
rect 0 207200 400 207256
rect 31600 207200 32000 207256
rect 0 206920 400 206976
rect 31600 206920 32000 206976
rect 0 206640 400 206696
rect 31600 206640 32000 206696
rect 0 206360 400 206416
rect 31600 206360 32000 206416
rect 0 206080 400 206136
rect 31600 206080 32000 206136
rect 0 205800 400 205856
rect 31600 205800 32000 205856
rect 0 205520 400 205576
rect 31600 205520 32000 205576
rect 0 205240 400 205296
rect 31600 205240 32000 205296
rect 0 204960 400 205016
rect 31600 204960 32000 205016
rect 0 204680 400 204736
rect 31600 204680 32000 204736
rect 0 204400 400 204456
rect 31600 204400 32000 204456
rect 0 204120 400 204176
rect 31600 204120 32000 204176
rect 0 203840 400 203896
rect 31600 203840 32000 203896
rect 0 203560 400 203616
rect 31600 203560 32000 203616
rect 0 203280 400 203336
rect 31600 203280 32000 203336
rect 0 203000 400 203056
rect 31600 203000 32000 203056
rect 0 202720 400 202776
rect 31600 202720 32000 202776
rect 0 202440 400 202496
rect 31600 202440 32000 202496
rect 0 202160 400 202216
rect 31600 202160 32000 202216
rect 0 201880 400 201936
rect 31600 201880 32000 201936
rect 0 201600 400 201656
rect 31600 201600 32000 201656
rect 0 201320 400 201376
rect 31600 201320 32000 201376
rect 0 201040 400 201096
rect 31600 201040 32000 201096
rect 0 200760 400 200816
rect 31600 200760 32000 200816
rect 0 200480 400 200536
rect 31600 200480 32000 200536
rect 0 200200 400 200256
rect 31600 200200 32000 200256
rect 0 199920 400 199976
rect 31600 199920 32000 199976
rect 0 199640 400 199696
rect 31600 199640 32000 199696
rect 0 199360 400 199416
rect 31600 199360 32000 199416
rect 0 199080 400 199136
rect 31600 199080 32000 199136
rect 0 198800 400 198856
rect 31600 198800 32000 198856
rect 0 198520 400 198576
rect 31600 198520 32000 198576
rect 0 198240 400 198296
rect 31600 198240 32000 198296
rect 0 197960 400 198016
rect 31600 197960 32000 198016
rect 0 197680 400 197736
rect 31600 197680 32000 197736
rect 0 197400 400 197456
rect 31600 197400 32000 197456
rect 0 197120 400 197176
rect 31600 197120 32000 197176
rect 0 196840 400 196896
rect 31600 196840 32000 196896
rect 0 196560 400 196616
rect 31600 196560 32000 196616
rect 0 196280 400 196336
rect 31600 196280 32000 196336
rect 0 196000 400 196056
rect 31600 196000 32000 196056
rect 0 195720 400 195776
rect 31600 195720 32000 195776
rect 0 195440 400 195496
rect 31600 195440 32000 195496
rect 0 195160 400 195216
rect 31600 195160 32000 195216
rect 0 194880 400 194936
rect 31600 194880 32000 194936
rect 0 194600 400 194656
rect 31600 194600 32000 194656
rect 0 194320 400 194376
rect 31600 194320 32000 194376
rect 0 194040 400 194096
rect 31600 194040 32000 194096
rect 0 193760 400 193816
rect 31600 193760 32000 193816
rect 0 193480 400 193536
rect 31600 193480 32000 193536
rect 0 193200 400 193256
rect 31600 193200 32000 193256
rect 0 192920 400 192976
rect 31600 192920 32000 192976
rect 0 192640 400 192696
rect 31600 192640 32000 192696
rect 0 192360 400 192416
rect 31600 192360 32000 192416
rect 0 192080 400 192136
rect 31600 192080 32000 192136
rect 0 191800 400 191856
rect 31600 191800 32000 191856
rect 0 191520 400 191576
rect 31600 191520 32000 191576
rect 0 191240 400 191296
rect 31600 191240 32000 191296
rect 0 190960 400 191016
rect 31600 190960 32000 191016
rect 0 190680 400 190736
rect 31600 190680 32000 190736
rect 0 190400 400 190456
rect 31600 190400 32000 190456
rect 0 190120 400 190176
rect 31600 190120 32000 190176
rect 0 189840 400 189896
rect 31600 189840 32000 189896
rect 0 189560 400 189616
rect 31600 189560 32000 189616
rect 0 189280 400 189336
rect 31600 189280 32000 189336
rect 0 189000 400 189056
rect 31600 189000 32000 189056
rect 0 188720 400 188776
rect 31600 188720 32000 188776
rect 0 188440 400 188496
rect 31600 188440 32000 188496
rect 0 188160 400 188216
rect 31600 188160 32000 188216
rect 0 187880 400 187936
rect 31600 187880 32000 187936
rect 0 187600 400 187656
rect 31600 187600 32000 187656
rect 0 187320 400 187376
rect 31600 187320 32000 187376
rect 0 187040 400 187096
rect 31600 187040 32000 187096
rect 0 186760 400 186816
rect 31600 186760 32000 186816
rect 0 186480 400 186536
rect 31600 186480 32000 186536
rect 0 186200 400 186256
rect 31600 186200 32000 186256
rect 0 185920 400 185976
rect 31600 185920 32000 185976
rect 0 185640 400 185696
rect 31600 185640 32000 185696
rect 0 185360 400 185416
rect 31600 185360 32000 185416
rect 0 185080 400 185136
rect 31600 185080 32000 185136
rect 0 184800 400 184856
rect 31600 184800 32000 184856
rect 0 184520 400 184576
rect 31600 184520 32000 184576
rect 0 184240 400 184296
rect 31600 184240 32000 184296
rect 0 183960 400 184016
rect 31600 183960 32000 184016
rect 0 183680 400 183736
rect 31600 183680 32000 183736
rect 0 183400 400 183456
rect 31600 183400 32000 183456
rect 0 183120 400 183176
rect 31600 183120 32000 183176
rect 0 182840 400 182896
rect 31600 182840 32000 182896
rect 0 182560 400 182616
rect 31600 182560 32000 182616
rect 0 182280 400 182336
rect 31600 182280 32000 182336
rect 0 182000 400 182056
rect 31600 182000 32000 182056
rect 0 181720 400 181776
rect 31600 181720 32000 181776
rect 0 181440 400 181496
rect 31600 181440 32000 181496
rect 0 181160 400 181216
rect 31600 181160 32000 181216
rect 0 180880 400 180936
rect 31600 180880 32000 180936
rect 0 180600 400 180656
rect 31600 180600 32000 180656
rect 0 180320 400 180376
rect 31600 180320 32000 180376
rect 0 180040 400 180096
rect 31600 180040 32000 180096
rect 0 179760 400 179816
rect 31600 179760 32000 179816
rect 0 179480 400 179536
rect 31600 179480 32000 179536
rect 0 179200 400 179256
rect 31600 179200 32000 179256
rect 0 178920 400 178976
rect 31600 178920 32000 178976
rect 0 178640 400 178696
rect 31600 178640 32000 178696
rect 0 178360 400 178416
rect 31600 178360 32000 178416
rect 0 178080 400 178136
rect 31600 178080 32000 178136
rect 0 177800 400 177856
rect 31600 177800 32000 177856
rect 0 177520 400 177576
rect 31600 177520 32000 177576
rect 0 177240 400 177296
rect 31600 177240 32000 177296
rect 0 176960 400 177016
rect 31600 176960 32000 177016
rect 0 176680 400 176736
rect 31600 176680 32000 176736
rect 0 176400 400 176456
rect 31600 176400 32000 176456
rect 0 176120 400 176176
rect 31600 176120 32000 176176
rect 0 175840 400 175896
rect 31600 175840 32000 175896
rect 0 175560 400 175616
rect 31600 175560 32000 175616
rect 0 175280 400 175336
rect 31600 175280 32000 175336
rect 0 175000 400 175056
rect 31600 175000 32000 175056
rect 0 174720 400 174776
rect 31600 174720 32000 174776
rect 0 174440 400 174496
rect 31600 174440 32000 174496
rect 0 174160 400 174216
rect 31600 174160 32000 174216
rect 0 173880 400 173936
rect 31600 173880 32000 173936
rect 0 173600 400 173656
rect 31600 173600 32000 173656
rect 0 173320 400 173376
rect 31600 173320 32000 173376
rect 0 173040 400 173096
rect 31600 173040 32000 173096
rect 0 172760 400 172816
rect 31600 172760 32000 172816
rect 0 172480 400 172536
rect 31600 172480 32000 172536
rect 0 172200 400 172256
rect 31600 172200 32000 172256
rect 0 171920 400 171976
rect 31600 171920 32000 171976
rect 0 171640 400 171696
rect 31600 171640 32000 171696
rect 0 171360 400 171416
rect 31600 171360 32000 171416
rect 0 171080 400 171136
rect 31600 171080 32000 171136
rect 0 170800 400 170856
rect 31600 170800 32000 170856
rect 0 170520 400 170576
rect 31600 170520 32000 170576
rect 0 170240 400 170296
rect 31600 170240 32000 170296
rect 0 169960 400 170016
rect 31600 169960 32000 170016
rect 0 169680 400 169736
rect 31600 169680 32000 169736
rect 0 169400 400 169456
rect 31600 169400 32000 169456
rect 0 169120 400 169176
rect 31600 169120 32000 169176
rect 0 168840 400 168896
rect 31600 168840 32000 168896
rect 0 168560 400 168616
rect 31600 168560 32000 168616
rect 0 168280 400 168336
rect 31600 168280 32000 168336
rect 0 168000 400 168056
rect 31600 168000 32000 168056
rect 0 167720 400 167776
rect 31600 167720 32000 167776
rect 0 167440 400 167496
rect 31600 167440 32000 167496
rect 0 167160 400 167216
rect 31600 167160 32000 167216
rect 0 166880 400 166936
rect 31600 166880 32000 166936
rect 0 166600 400 166656
rect 31600 166600 32000 166656
rect 0 166320 400 166376
rect 31600 166320 32000 166376
rect 0 166040 400 166096
rect 31600 166040 32000 166096
rect 0 165760 400 165816
rect 31600 165760 32000 165816
rect 0 165480 400 165536
rect 31600 165480 32000 165536
rect 0 165200 400 165256
rect 31600 165200 32000 165256
rect 0 164920 400 164976
rect 31600 164920 32000 164976
rect 0 164640 400 164696
rect 31600 164640 32000 164696
rect 0 164360 400 164416
rect 31600 164360 32000 164416
rect 0 164080 400 164136
rect 31600 164080 32000 164136
rect 0 163800 400 163856
rect 31600 163800 32000 163856
rect 0 163520 400 163576
rect 31600 163520 32000 163576
rect 0 163240 400 163296
rect 31600 163240 32000 163296
rect 0 162960 400 163016
rect 31600 162960 32000 163016
rect 0 162680 400 162736
rect 31600 162680 32000 162736
rect 0 162400 400 162456
rect 31600 162400 32000 162456
rect 0 162120 400 162176
rect 31600 162120 32000 162176
rect 0 161840 400 161896
rect 31600 161840 32000 161896
rect 0 161560 400 161616
rect 31600 161560 32000 161616
rect 0 161280 400 161336
rect 31600 161280 32000 161336
rect 0 161000 400 161056
rect 31600 161000 32000 161056
rect 0 160720 400 160776
rect 31600 160720 32000 160776
rect 0 160440 400 160496
rect 31600 160440 32000 160496
rect 0 160160 400 160216
rect 31600 160160 32000 160216
rect 0 159880 400 159936
rect 31600 159880 32000 159936
rect 0 159600 400 159656
rect 31600 159600 32000 159656
rect 0 159320 400 159376
rect 31600 159320 32000 159376
rect 0 159040 400 159096
rect 31600 159040 32000 159096
rect 0 158760 400 158816
rect 31600 158760 32000 158816
rect 0 158480 400 158536
rect 31600 158480 32000 158536
rect 0 158200 400 158256
rect 31600 158200 32000 158256
rect 0 157920 400 157976
rect 31600 157920 32000 157976
rect 0 157640 400 157696
rect 31600 157640 32000 157696
rect 0 157360 400 157416
rect 31600 157360 32000 157416
rect 0 157080 400 157136
rect 31600 157080 32000 157136
rect 0 156800 400 156856
rect 31600 156800 32000 156856
rect 0 156520 400 156576
rect 31600 156520 32000 156576
rect 0 156240 400 156296
rect 31600 156240 32000 156296
rect 0 155960 400 156016
rect 31600 155960 32000 156016
rect 0 155680 400 155736
rect 31600 155680 32000 155736
rect 0 155400 400 155456
rect 31600 155400 32000 155456
rect 0 155120 400 155176
rect 31600 155120 32000 155176
rect 0 154840 400 154896
rect 31600 154840 32000 154896
rect 0 154560 400 154616
rect 31600 154560 32000 154616
rect 0 154280 400 154336
rect 31600 154280 32000 154336
rect 0 154000 400 154056
rect 31600 154000 32000 154056
rect 0 153720 400 153776
rect 31600 153720 32000 153776
rect 0 153440 400 153496
rect 31600 153440 32000 153496
rect 0 153160 400 153216
rect 31600 153160 32000 153216
rect 0 152880 400 152936
rect 31600 152880 32000 152936
rect 0 152600 400 152656
rect 31600 152600 32000 152656
rect 0 152320 400 152376
rect 31600 152320 32000 152376
rect 0 152040 400 152096
rect 31600 152040 32000 152096
rect 0 151760 400 151816
rect 31600 151760 32000 151816
rect 0 151480 400 151536
rect 31600 151480 32000 151536
rect 0 151200 400 151256
rect 31600 151200 32000 151256
rect 0 150920 400 150976
rect 31600 150920 32000 150976
rect 0 150640 400 150696
rect 31600 150640 32000 150696
rect 0 150360 400 150416
rect 31600 150360 32000 150416
rect 0 150080 400 150136
rect 31600 150080 32000 150136
rect 0 149800 400 149856
rect 31600 149800 32000 149856
rect 0 149520 400 149576
rect 31600 149520 32000 149576
rect 0 149240 400 149296
rect 31600 149240 32000 149296
rect 0 148960 400 149016
rect 31600 148960 32000 149016
rect 0 148680 400 148736
rect 31600 148680 32000 148736
rect 0 148400 400 148456
rect 31600 148400 32000 148456
rect 0 148120 400 148176
rect 31600 148120 32000 148176
rect 0 147840 400 147896
rect 31600 147840 32000 147896
rect 0 147560 400 147616
rect 31600 147560 32000 147616
rect 0 147280 400 147336
rect 31600 147280 32000 147336
rect 0 147000 400 147056
rect 31600 147000 32000 147056
rect 0 146720 400 146776
rect 31600 146720 32000 146776
rect 0 146440 400 146496
rect 31600 146440 32000 146496
rect 0 146160 400 146216
rect 31600 146160 32000 146216
rect 0 145880 400 145936
rect 31600 145880 32000 145936
rect 0 145600 400 145656
rect 31600 145600 32000 145656
rect 0 145320 400 145376
rect 31600 145320 32000 145376
rect 0 145040 400 145096
rect 31600 145040 32000 145096
rect 0 144760 400 144816
rect 31600 144760 32000 144816
rect 0 144480 400 144536
rect 31600 144480 32000 144536
rect 0 144200 400 144256
rect 31600 144200 32000 144256
rect 0 143920 400 143976
rect 31600 143920 32000 143976
rect 0 143640 400 143696
rect 31600 143640 32000 143696
rect 0 143360 400 143416
rect 31600 143360 32000 143416
rect 0 143080 400 143136
rect 31600 143080 32000 143136
rect 0 142800 400 142856
rect 31600 142800 32000 142856
rect 0 142520 400 142576
rect 31600 142520 32000 142576
rect 0 142240 400 142296
rect 31600 142240 32000 142296
rect 0 141960 400 142016
rect 31600 141960 32000 142016
rect 0 141680 400 141736
rect 31600 141680 32000 141736
rect 0 141400 400 141456
rect 31600 141400 32000 141456
rect 0 141120 400 141176
rect 31600 141120 32000 141176
rect 0 140840 400 140896
rect 31600 140840 32000 140896
rect 0 140560 400 140616
rect 31600 140560 32000 140616
rect 0 140280 400 140336
rect 31600 140280 32000 140336
rect 0 140000 400 140056
rect 31600 140000 32000 140056
rect 0 139720 400 139776
rect 31600 139720 32000 139776
rect 0 139440 400 139496
rect 31600 139440 32000 139496
rect 0 139160 400 139216
rect 31600 139160 32000 139216
rect 0 138880 400 138936
rect 31600 138880 32000 138936
rect 0 138600 400 138656
rect 31600 138600 32000 138656
rect 0 138320 400 138376
rect 31600 138320 32000 138376
rect 0 138040 400 138096
rect 31600 138040 32000 138096
rect 0 137760 400 137816
rect 31600 137760 32000 137816
rect 0 137480 400 137536
rect 31600 137480 32000 137536
rect 0 137200 400 137256
rect 31600 137200 32000 137256
rect 0 136920 400 136976
rect 31600 136920 32000 136976
rect 0 136640 400 136696
rect 31600 136640 32000 136696
rect 0 136360 400 136416
rect 31600 136360 32000 136416
rect 0 136080 400 136136
rect 31600 136080 32000 136136
rect 0 135800 400 135856
rect 31600 135800 32000 135856
rect 0 135520 400 135576
rect 31600 135520 32000 135576
rect 0 135240 400 135296
rect 31600 135240 32000 135296
rect 0 134960 400 135016
rect 31600 134960 32000 135016
rect 0 134680 400 134736
rect 31600 134680 32000 134736
rect 0 134400 400 134456
rect 31600 134400 32000 134456
rect 0 134120 400 134176
rect 31600 134120 32000 134176
rect 0 133840 400 133896
rect 31600 133840 32000 133896
rect 0 133560 400 133616
rect 31600 133560 32000 133616
rect 0 133280 400 133336
rect 31600 133280 32000 133336
rect 0 133000 400 133056
rect 31600 133000 32000 133056
rect 0 132720 400 132776
rect 31600 132720 32000 132776
rect 0 132440 400 132496
rect 31600 132440 32000 132496
rect 0 132160 400 132216
rect 31600 132160 32000 132216
rect 0 131880 400 131936
rect 31600 131880 32000 131936
rect 0 131600 400 131656
rect 31600 131600 32000 131656
rect 0 131320 400 131376
rect 31600 131320 32000 131376
rect 0 131040 400 131096
rect 31600 131040 32000 131096
rect 0 130760 400 130816
rect 31600 130760 32000 130816
rect 0 130480 400 130536
rect 31600 130480 32000 130536
rect 0 130200 400 130256
rect 31600 130200 32000 130256
rect 0 129920 400 129976
rect 31600 129920 32000 129976
rect 0 129640 400 129696
rect 31600 129640 32000 129696
rect 0 129360 400 129416
rect 31600 129360 32000 129416
rect 0 129080 400 129136
rect 31600 129080 32000 129136
rect 0 128800 400 128856
rect 31600 128800 32000 128856
rect 0 128520 400 128576
rect 31600 128520 32000 128576
rect 0 128240 400 128296
rect 31600 128240 32000 128296
rect 0 127960 400 128016
rect 31600 127960 32000 128016
rect 0 127680 400 127736
rect 31600 127680 32000 127736
rect 0 127400 400 127456
rect 31600 127400 32000 127456
rect 0 127120 400 127176
rect 31600 127120 32000 127176
rect 0 126840 400 126896
rect 31600 126840 32000 126896
rect 0 126560 400 126616
rect 31600 126560 32000 126616
rect 0 126280 400 126336
rect 31600 126280 32000 126336
rect 0 126000 400 126056
rect 31600 126000 32000 126056
rect 0 125720 400 125776
rect 31600 125720 32000 125776
rect 0 125440 400 125496
rect 31600 125440 32000 125496
rect 0 125160 400 125216
rect 31600 125160 32000 125216
rect 0 124880 400 124936
rect 31600 124880 32000 124936
rect 0 124600 400 124656
rect 31600 124600 32000 124656
rect 0 124320 400 124376
rect 31600 124320 32000 124376
rect 0 124040 400 124096
rect 31600 124040 32000 124096
rect 0 123760 400 123816
rect 31600 123760 32000 123816
rect 0 123480 400 123536
rect 31600 123480 32000 123536
rect 0 123200 400 123256
rect 31600 123200 32000 123256
rect 0 122920 400 122976
rect 31600 122920 32000 122976
rect 0 122640 400 122696
rect 31600 122640 32000 122696
rect 0 122360 400 122416
rect 31600 122360 32000 122416
rect 0 122080 400 122136
rect 31600 122080 32000 122136
rect 0 121800 400 121856
rect 31600 121800 32000 121856
rect 0 121520 400 121576
rect 31600 121520 32000 121576
rect 0 121240 400 121296
rect 31600 121240 32000 121296
rect 0 120960 400 121016
rect 31600 120960 32000 121016
rect 0 120680 400 120736
rect 31600 120680 32000 120736
rect 0 120400 400 120456
rect 31600 120400 32000 120456
rect 0 120120 400 120176
rect 31600 120120 32000 120176
rect 0 119840 400 119896
rect 31600 119840 32000 119896
rect 0 119560 400 119616
rect 31600 119560 32000 119616
rect 0 119280 400 119336
rect 31600 119280 32000 119336
rect 0 119000 400 119056
rect 31600 119000 32000 119056
rect 0 118720 400 118776
rect 31600 118720 32000 118776
rect 0 118440 400 118496
rect 31600 118440 32000 118496
rect 0 118160 400 118216
rect 31600 118160 32000 118216
rect 0 117880 400 117936
rect 31600 117880 32000 117936
rect 0 117600 400 117656
rect 31600 117600 32000 117656
rect 0 117320 400 117376
rect 31600 117320 32000 117376
rect 0 117040 400 117096
rect 31600 117040 32000 117096
rect 0 116760 400 116816
rect 31600 116760 32000 116816
rect 0 116480 400 116536
rect 31600 116480 32000 116536
rect 0 116200 400 116256
rect 31600 116200 32000 116256
rect 0 115920 400 115976
rect 31600 115920 32000 115976
rect 0 115640 400 115696
rect 31600 115640 32000 115696
rect 0 115360 400 115416
rect 31600 115360 32000 115416
rect 0 115080 400 115136
rect 31600 115080 32000 115136
rect 0 114800 400 114856
rect 31600 114800 32000 114856
rect 0 114520 400 114576
rect 31600 114520 32000 114576
rect 0 114240 400 114296
rect 31600 114240 32000 114296
rect 0 113960 400 114016
rect 31600 113960 32000 114016
rect 0 113680 400 113736
rect 31600 113680 32000 113736
rect 0 113400 400 113456
rect 31600 113400 32000 113456
rect 0 113120 400 113176
rect 31600 113120 32000 113176
rect 0 112840 400 112896
rect 31600 112840 32000 112896
rect 0 112560 400 112616
rect 31600 112560 32000 112616
rect 0 112280 400 112336
rect 31600 112280 32000 112336
rect 0 112000 400 112056
rect 31600 112000 32000 112056
rect 0 111720 400 111776
rect 31600 111720 32000 111776
rect 0 111440 400 111496
rect 31600 111440 32000 111496
rect 0 111160 400 111216
rect 31600 111160 32000 111216
rect 0 110880 400 110936
rect 31600 110880 32000 110936
rect 0 110600 400 110656
rect 31600 110600 32000 110656
rect 0 110320 400 110376
rect 31600 110320 32000 110376
rect 0 110040 400 110096
rect 31600 110040 32000 110096
rect 0 109760 400 109816
rect 31600 109760 32000 109816
rect 0 109480 400 109536
rect 31600 109480 32000 109536
rect 0 109200 400 109256
rect 31600 109200 32000 109256
rect 0 108920 400 108976
rect 31600 108920 32000 108976
rect 0 108640 400 108696
rect 31600 108640 32000 108696
rect 0 108360 400 108416
rect 31600 108360 32000 108416
rect 0 108080 400 108136
rect 31600 108080 32000 108136
rect 0 107800 400 107856
rect 31600 107800 32000 107856
rect 0 107520 400 107576
rect 31600 107520 32000 107576
rect 0 107240 400 107296
rect 31600 107240 32000 107296
rect 0 106960 400 107016
rect 31600 106960 32000 107016
rect 0 106680 400 106736
rect 31600 106680 32000 106736
rect 0 106400 400 106456
rect 31600 106400 32000 106456
rect 0 106120 400 106176
rect 31600 106120 32000 106176
rect 0 105840 400 105896
rect 31600 105840 32000 105896
rect 0 105560 400 105616
rect 31600 105560 32000 105616
rect 0 105280 400 105336
rect 31600 105280 32000 105336
rect 0 105000 400 105056
rect 31600 105000 32000 105056
rect 0 104720 400 104776
rect 31600 104720 32000 104776
rect 0 104440 400 104496
rect 31600 104440 32000 104496
rect 0 104160 400 104216
rect 31600 104160 32000 104216
rect 0 103880 400 103936
rect 31600 103880 32000 103936
rect 0 103600 400 103656
rect 31600 103600 32000 103656
rect 0 103320 400 103376
rect 31600 103320 32000 103376
rect 0 103040 400 103096
rect 31600 103040 32000 103096
rect 0 102760 400 102816
rect 31600 102760 32000 102816
rect 0 102480 400 102536
rect 31600 102480 32000 102536
rect 0 102200 400 102256
rect 31600 102200 32000 102256
rect 0 101920 400 101976
rect 31600 101920 32000 101976
rect 0 101640 400 101696
rect 31600 101640 32000 101696
rect 0 101360 400 101416
rect 31600 101360 32000 101416
rect 0 101080 400 101136
rect 31600 101080 32000 101136
rect 0 100800 400 100856
rect 31600 100800 32000 100856
rect 0 100520 400 100576
rect 31600 100520 32000 100576
rect 0 100240 400 100296
rect 31600 100240 32000 100296
rect 0 99960 400 100016
rect 31600 99960 32000 100016
rect 0 99680 400 99736
rect 31600 99680 32000 99736
rect 0 99400 400 99456
rect 31600 99400 32000 99456
rect 0 99120 400 99176
rect 31600 99120 32000 99176
rect 0 98840 400 98896
rect 31600 98840 32000 98896
rect 0 98560 400 98616
rect 31600 98560 32000 98616
rect 0 98280 400 98336
rect 31600 98280 32000 98336
rect 0 98000 400 98056
rect 31600 98000 32000 98056
rect 0 97720 400 97776
rect 31600 97720 32000 97776
rect 0 97440 400 97496
rect 31600 97440 32000 97496
rect 0 97160 400 97216
rect 31600 97160 32000 97216
rect 0 96880 400 96936
rect 31600 96880 32000 96936
rect 0 96600 400 96656
rect 31600 96600 32000 96656
rect 0 96320 400 96376
rect 31600 96320 32000 96376
rect 0 96040 400 96096
rect 31600 96040 32000 96096
rect 0 95760 400 95816
rect 31600 95760 32000 95816
rect 0 95480 400 95536
rect 31600 95480 32000 95536
rect 0 95200 400 95256
rect 31600 95200 32000 95256
rect 0 94920 400 94976
rect 31600 94920 32000 94976
rect 0 94640 400 94696
rect 31600 94640 32000 94696
rect 0 94360 400 94416
rect 31600 94360 32000 94416
rect 0 94080 400 94136
rect 31600 94080 32000 94136
rect 0 93800 400 93856
rect 31600 93800 32000 93856
rect 0 93520 400 93576
rect 31600 93520 32000 93576
rect 0 93240 400 93296
rect 31600 93240 32000 93296
rect 0 92960 400 93016
rect 31600 92960 32000 93016
rect 0 92680 400 92736
rect 31600 92680 32000 92736
rect 0 92400 400 92456
rect 31600 92400 32000 92456
rect 0 92120 400 92176
rect 31600 92120 32000 92176
rect 0 91840 400 91896
rect 31600 91840 32000 91896
rect 0 91560 400 91616
rect 31600 91560 32000 91616
rect 0 91280 400 91336
rect 31600 91280 32000 91336
rect 0 91000 400 91056
rect 31600 91000 32000 91056
rect 0 90720 400 90776
rect 31600 90720 32000 90776
rect 0 90440 400 90496
rect 31600 90440 32000 90496
rect 0 90160 400 90216
rect 31600 90160 32000 90216
rect 0 89880 400 89936
rect 31600 89880 32000 89936
rect 0 89600 400 89656
rect 31600 89600 32000 89656
rect 0 89320 400 89376
rect 31600 89320 32000 89376
rect 0 89040 400 89096
rect 31600 89040 32000 89096
rect 0 88760 400 88816
rect 31600 88760 32000 88816
rect 0 88480 400 88536
rect 31600 88480 32000 88536
rect 0 88200 400 88256
rect 31600 88200 32000 88256
rect 0 87920 400 87976
rect 31600 87920 32000 87976
rect 0 87640 400 87696
rect 31600 87640 32000 87696
rect 0 87360 400 87416
rect 31600 87360 32000 87416
rect 0 87080 400 87136
rect 31600 87080 32000 87136
rect 0 86800 400 86856
rect 31600 86800 32000 86856
rect 0 86520 400 86576
rect 31600 86520 32000 86576
rect 0 86240 400 86296
rect 31600 86240 32000 86296
rect 0 85960 400 86016
rect 31600 85960 32000 86016
rect 0 85680 400 85736
rect 31600 85680 32000 85736
rect 0 85400 400 85456
rect 31600 85400 32000 85456
rect 0 85120 400 85176
rect 31600 85120 32000 85176
rect 0 84840 400 84896
rect 31600 84840 32000 84896
rect 0 84560 400 84616
rect 31600 84560 32000 84616
rect 0 84280 400 84336
rect 31600 84280 32000 84336
rect 0 84000 400 84056
rect 31600 84000 32000 84056
rect 0 83720 400 83776
rect 31600 83720 32000 83776
rect 0 83440 400 83496
rect 31600 83440 32000 83496
rect 0 83160 400 83216
rect 31600 83160 32000 83216
rect 0 82880 400 82936
rect 31600 82880 32000 82936
rect 0 82600 400 82656
rect 31600 82600 32000 82656
rect 0 82320 400 82376
rect 31600 82320 32000 82376
rect 0 82040 400 82096
rect 31600 82040 32000 82096
rect 0 81760 400 81816
rect 31600 81760 32000 81816
rect 0 81480 400 81536
rect 31600 81480 32000 81536
rect 0 81200 400 81256
rect 31600 81200 32000 81256
rect 0 80920 400 80976
rect 31600 80920 32000 80976
rect 0 80640 400 80696
rect 31600 80640 32000 80696
rect 0 80360 400 80416
rect 31600 80360 32000 80416
rect 0 80080 400 80136
rect 31600 80080 32000 80136
rect 0 79800 400 79856
rect 31600 79800 32000 79856
rect 0 79520 400 79576
rect 31600 79520 32000 79576
rect 0 79240 400 79296
rect 31600 79240 32000 79296
rect 0 78960 400 79016
rect 31600 78960 32000 79016
rect 0 78680 400 78736
rect 31600 78680 32000 78736
rect 0 78400 400 78456
rect 31600 78400 32000 78456
rect 0 78120 400 78176
rect 31600 78120 32000 78176
rect 0 77840 400 77896
rect 31600 77840 32000 77896
rect 0 77560 400 77616
rect 31600 77560 32000 77616
rect 0 77280 400 77336
rect 31600 77280 32000 77336
rect 0 77000 400 77056
rect 31600 77000 32000 77056
rect 0 76720 400 76776
rect 31600 76720 32000 76776
rect 0 76440 400 76496
rect 31600 76440 32000 76496
rect 0 76160 400 76216
rect 31600 76160 32000 76216
rect 0 75880 400 75936
rect 31600 75880 32000 75936
rect 0 75600 400 75656
rect 31600 75600 32000 75656
rect 0 75320 400 75376
rect 31600 75320 32000 75376
rect 0 75040 400 75096
rect 31600 75040 32000 75096
rect 0 74760 400 74816
rect 31600 74760 32000 74816
rect 0 74480 400 74536
rect 31600 74480 32000 74536
rect 0 74200 400 74256
rect 31600 74200 32000 74256
rect 0 73920 400 73976
rect 31600 73920 32000 73976
rect 0 73640 400 73696
rect 31600 73640 32000 73696
rect 0 73360 400 73416
rect 31600 73360 32000 73416
rect 0 73080 400 73136
rect 31600 73080 32000 73136
rect 0 72800 400 72856
rect 31600 72800 32000 72856
rect 0 72520 400 72576
rect 31600 72520 32000 72576
rect 0 72240 400 72296
rect 31600 72240 32000 72296
rect 0 71960 400 72016
rect 31600 71960 32000 72016
rect 0 71680 400 71736
rect 31600 71680 32000 71736
rect 0 71400 400 71456
rect 31600 71400 32000 71456
rect 0 71120 400 71176
rect 31600 71120 32000 71176
rect 0 70840 400 70896
rect 31600 70840 32000 70896
rect 0 70560 400 70616
rect 31600 70560 32000 70616
rect 0 70280 400 70336
rect 31600 70280 32000 70336
rect 0 70000 400 70056
rect 31600 70000 32000 70056
rect 0 69720 400 69776
rect 31600 69720 32000 69776
rect 0 69440 400 69496
rect 31600 69440 32000 69496
rect 0 69160 400 69216
rect 31600 69160 32000 69216
rect 0 68880 400 68936
rect 31600 68880 32000 68936
rect 0 68600 400 68656
rect 31600 68600 32000 68656
rect 0 68320 400 68376
rect 31600 68320 32000 68376
rect 0 68040 400 68096
rect 31600 68040 32000 68096
rect 0 67760 400 67816
rect 31600 67760 32000 67816
rect 0 67480 400 67536
rect 31600 67480 32000 67536
rect 0 67200 400 67256
rect 31600 67200 32000 67256
rect 0 66920 400 66976
rect 31600 66920 32000 66976
rect 0 66640 400 66696
rect 31600 66640 32000 66696
rect 0 66360 400 66416
rect 31600 66360 32000 66416
rect 0 66080 400 66136
rect 31600 66080 32000 66136
rect 0 65800 400 65856
rect 31600 65800 32000 65856
rect 0 65520 400 65576
rect 31600 65520 32000 65576
rect 0 65240 400 65296
rect 31600 65240 32000 65296
rect 0 64960 400 65016
rect 31600 64960 32000 65016
rect 0 64680 400 64736
rect 31600 64680 32000 64736
rect 0 64400 400 64456
rect 31600 64400 32000 64456
rect 0 64120 400 64176
rect 31600 64120 32000 64176
rect 0 63840 400 63896
rect 31600 63840 32000 63896
rect 0 63560 400 63616
rect 31600 63560 32000 63616
rect 0 63280 400 63336
rect 31600 63280 32000 63336
rect 0 63000 400 63056
rect 31600 63000 32000 63056
rect 0 62720 400 62776
rect 31600 62720 32000 62776
rect 0 62440 400 62496
rect 31600 62440 32000 62496
rect 0 62160 400 62216
rect 31600 62160 32000 62216
rect 0 61880 400 61936
rect 31600 61880 32000 61936
rect 0 61600 400 61656
rect 31600 61600 32000 61656
rect 0 61320 400 61376
rect 31600 61320 32000 61376
rect 0 61040 400 61096
rect 31600 61040 32000 61096
rect 0 60760 400 60816
rect 31600 60760 32000 60816
rect 0 60480 400 60536
rect 31600 60480 32000 60536
rect 0 60200 400 60256
rect 31600 60200 32000 60256
rect 0 59920 400 59976
rect 31600 59920 32000 59976
rect 0 59640 400 59696
rect 31600 59640 32000 59696
rect 0 59360 400 59416
rect 31600 59360 32000 59416
rect 0 59080 400 59136
rect 31600 59080 32000 59136
rect 0 58800 400 58856
rect 31600 58800 32000 58856
rect 0 58520 400 58576
rect 31600 58520 32000 58576
rect 0 58240 400 58296
rect 31600 58240 32000 58296
rect 0 57960 400 58016
rect 31600 57960 32000 58016
rect 0 57680 400 57736
rect 31600 57680 32000 57736
rect 0 57400 400 57456
rect 31600 57400 32000 57456
rect 0 57120 400 57176
rect 31600 57120 32000 57176
rect 0 56840 400 56896
rect 31600 56840 32000 56896
rect 0 56560 400 56616
rect 31600 56560 32000 56616
rect 0 56280 400 56336
rect 31600 56280 32000 56336
rect 0 56000 400 56056
rect 31600 56000 32000 56056
rect 0 55720 400 55776
rect 31600 55720 32000 55776
rect 0 55440 400 55496
rect 31600 55440 32000 55496
rect 0 55160 400 55216
rect 31600 55160 32000 55216
rect 0 54880 400 54936
rect 31600 54880 32000 54936
rect 0 54600 400 54656
rect 31600 54600 32000 54656
rect 0 54320 400 54376
rect 31600 54320 32000 54376
rect 0 54040 400 54096
rect 31600 54040 32000 54096
rect 0 53760 400 53816
rect 31600 53760 32000 53816
rect 0 53480 400 53536
rect 31600 53480 32000 53536
rect 0 53200 400 53256
rect 31600 53200 32000 53256
rect 0 52920 400 52976
rect 31600 52920 32000 52976
rect 0 52640 400 52696
rect 31600 52640 32000 52696
rect 0 52360 400 52416
rect 31600 52360 32000 52416
rect 0 52080 400 52136
rect 31600 52080 32000 52136
rect 0 51800 400 51856
rect 31600 51800 32000 51856
rect 0 51520 400 51576
rect 31600 51520 32000 51576
rect 0 51240 400 51296
rect 31600 51240 32000 51296
rect 0 50960 400 51016
rect 31600 50960 32000 51016
rect 0 50680 400 50736
rect 31600 50680 32000 50736
rect 0 50400 400 50456
rect 31600 50400 32000 50456
rect 0 50120 400 50176
rect 31600 50120 32000 50176
rect 0 49840 400 49896
rect 31600 49840 32000 49896
rect 0 49560 400 49616
rect 31600 49560 32000 49616
rect 0 49280 400 49336
rect 31600 49280 32000 49336
rect 0 49000 400 49056
rect 31600 49000 32000 49056
rect 0 48720 400 48776
rect 31600 48720 32000 48776
rect 0 48440 400 48496
rect 31600 48440 32000 48496
rect 0 48160 400 48216
rect 31600 48160 32000 48216
rect 0 47880 400 47936
rect 31600 47880 32000 47936
rect 0 47600 400 47656
rect 31600 47600 32000 47656
rect 0 47320 400 47376
rect 31600 47320 32000 47376
rect 0 47040 400 47096
rect 31600 47040 32000 47096
rect 0 46760 400 46816
rect 31600 46760 32000 46816
rect 0 46480 400 46536
rect 31600 46480 32000 46536
rect 0 46200 400 46256
rect 31600 46200 32000 46256
rect 0 45920 400 45976
rect 31600 45920 32000 45976
rect 0 45640 400 45696
rect 31600 45640 32000 45696
rect 0 45360 400 45416
rect 31600 45360 32000 45416
rect 0 45080 400 45136
rect 31600 45080 32000 45136
rect 0 44800 400 44856
rect 31600 44800 32000 44856
rect 0 44520 400 44576
rect 31600 44520 32000 44576
rect 0 44240 400 44296
rect 31600 44240 32000 44296
rect 0 43960 400 44016
rect 31600 43960 32000 44016
rect 0 43680 400 43736
rect 31600 43680 32000 43736
rect 0 43400 400 43456
rect 31600 43400 32000 43456
rect 0 43120 400 43176
rect 31600 43120 32000 43176
rect 0 42840 400 42896
rect 31600 42840 32000 42896
rect 0 42560 400 42616
rect 31600 42560 32000 42616
rect 0 42280 400 42336
rect 31600 42280 32000 42336
rect 0 42000 400 42056
rect 31600 42000 32000 42056
rect 0 41720 400 41776
rect 31600 41720 32000 41776
rect 0 41440 400 41496
rect 31600 41440 32000 41496
rect 0 41160 400 41216
rect 31600 41160 32000 41216
rect 0 40880 400 40936
rect 31600 40880 32000 40936
rect 0 40600 400 40656
rect 31600 40600 32000 40656
rect 0 40320 400 40376
rect 31600 40320 32000 40376
rect 0 40040 400 40096
rect 31600 40040 32000 40096
rect 0 39760 400 39816
rect 31600 39760 32000 39816
rect 0 39480 400 39536
rect 31600 39480 32000 39536
rect 0 39200 400 39256
rect 31600 39200 32000 39256
rect 0 38920 400 38976
rect 31600 38920 32000 38976
rect 0 38640 400 38696
rect 31600 38640 32000 38696
rect 0 38360 400 38416
rect 31600 38360 32000 38416
rect 0 38080 400 38136
rect 31600 38080 32000 38136
rect 0 37800 400 37856
rect 31600 37800 32000 37856
rect 0 37520 400 37576
rect 31600 37520 32000 37576
rect 0 37240 400 37296
rect 31600 37240 32000 37296
rect 0 36960 400 37016
rect 31600 36960 32000 37016
rect 0 36680 400 36736
rect 31600 36680 32000 36736
rect 0 36400 400 36456
rect 31600 36400 32000 36456
rect 0 36120 400 36176
rect 31600 36120 32000 36176
rect 0 35840 400 35896
rect 31600 35840 32000 35896
rect 0 35560 400 35616
rect 31600 35560 32000 35616
rect 0 35280 400 35336
rect 31600 35280 32000 35336
rect 0 35000 400 35056
rect 31600 35000 32000 35056
rect 0 34720 400 34776
rect 31600 34720 32000 34776
rect 0 34440 400 34496
rect 31600 34440 32000 34496
rect 0 34160 400 34216
rect 31600 34160 32000 34216
rect 0 33880 400 33936
rect 31600 33880 32000 33936
rect 0 33600 400 33656
rect 31600 33600 32000 33656
rect 0 33320 400 33376
rect 31600 33320 32000 33376
rect 0 33040 400 33096
rect 31600 33040 32000 33096
rect 0 32760 400 32816
rect 31600 32760 32000 32816
rect 0 32480 400 32536
rect 31600 32480 32000 32536
rect 0 32200 400 32256
rect 31600 32200 32000 32256
rect 0 31920 400 31976
rect 31600 31920 32000 31976
rect 0 31640 400 31696
rect 31600 31640 32000 31696
rect 0 31360 400 31416
rect 31600 31360 32000 31416
rect 0 31080 400 31136
rect 31600 31080 32000 31136
rect 0 30800 400 30856
rect 31600 30800 32000 30856
rect 0 30520 400 30576
rect 31600 30520 32000 30576
rect 0 30240 400 30296
rect 31600 30240 32000 30296
rect 0 29960 400 30016
rect 31600 29960 32000 30016
rect 0 29680 400 29736
rect 31600 29680 32000 29736
rect 0 29400 400 29456
rect 31600 29400 32000 29456
rect 0 29120 400 29176
rect 31600 29120 32000 29176
rect 0 28840 400 28896
rect 31600 28840 32000 28896
rect 0 28560 400 28616
rect 31600 28560 32000 28616
rect 0 28280 400 28336
rect 31600 28280 32000 28336
rect 0 28000 400 28056
rect 31600 28000 32000 28056
rect 0 27720 400 27776
rect 31600 27720 32000 27776
rect 0 27440 400 27496
rect 31600 27440 32000 27496
rect 0 27160 400 27216
rect 31600 27160 32000 27216
rect 0 26880 400 26936
rect 31600 26880 32000 26936
rect 0 26600 400 26656
rect 31600 26600 32000 26656
rect 0 26320 400 26376
rect 31600 26320 32000 26376
rect 0 26040 400 26096
rect 31600 26040 32000 26096
rect 0 25760 400 25816
rect 31600 25760 32000 25816
rect 0 25480 400 25536
rect 31600 25480 32000 25536
rect 0 25200 400 25256
rect 31600 25200 32000 25256
rect 0 24920 400 24976
rect 31600 24920 32000 24976
rect 0 24640 400 24696
rect 31600 24640 32000 24696
rect 0 24360 400 24416
rect 31600 24360 32000 24416
rect 0 24080 400 24136
rect 31600 24080 32000 24136
rect 0 23800 400 23856
rect 31600 23800 32000 23856
rect 0 23520 400 23576
rect 31600 23520 32000 23576
rect 0 23240 400 23296
rect 31600 23240 32000 23296
rect 0 22960 400 23016
rect 31600 22960 32000 23016
rect 0 22680 400 22736
rect 31600 22680 32000 22736
rect 0 22400 400 22456
rect 31600 22400 32000 22456
rect 0 22120 400 22176
rect 31600 22120 32000 22176
rect 0 21840 400 21896
rect 31600 21840 32000 21896
rect 0 21560 400 21616
rect 31600 21560 32000 21616
rect 0 21280 400 21336
rect 31600 21280 32000 21336
rect 0 21000 400 21056
rect 31600 21000 32000 21056
rect 0 20720 400 20776
rect 31600 20720 32000 20776
rect 0 20440 400 20496
rect 31600 20440 32000 20496
rect 0 20160 400 20216
rect 31600 20160 32000 20216
rect 0 19880 400 19936
rect 31600 19880 32000 19936
rect 0 19600 400 19656
rect 31600 19600 32000 19656
rect 0 19320 400 19376
rect 31600 19320 32000 19376
rect 0 19040 400 19096
rect 31600 19040 32000 19096
rect 0 18760 400 18816
rect 31600 18760 32000 18816
rect 0 18480 400 18536
rect 31600 18480 32000 18536
<< obsm3 >>
rect 233 251246 31799 268534
rect 430 251130 31570 251246
rect 233 250966 31799 251130
rect 430 250850 31570 250966
rect 233 250686 31799 250850
rect 430 250570 31570 250686
rect 233 250406 31799 250570
rect 430 250290 31570 250406
rect 233 250126 31799 250290
rect 430 250010 31570 250126
rect 233 249846 31799 250010
rect 430 249730 31570 249846
rect 233 249566 31799 249730
rect 430 249450 31570 249566
rect 233 249286 31799 249450
rect 430 249170 31570 249286
rect 233 249006 31799 249170
rect 430 248890 31570 249006
rect 233 248726 31799 248890
rect 430 248610 31570 248726
rect 233 248446 31799 248610
rect 430 248330 31570 248446
rect 233 248166 31799 248330
rect 430 248050 31570 248166
rect 233 247886 31799 248050
rect 430 247770 31570 247886
rect 233 247606 31799 247770
rect 430 247490 31570 247606
rect 233 247326 31799 247490
rect 430 247210 31570 247326
rect 233 247046 31799 247210
rect 430 246930 31570 247046
rect 233 246766 31799 246930
rect 430 246650 31570 246766
rect 233 246486 31799 246650
rect 430 246370 31570 246486
rect 233 246206 31799 246370
rect 430 246090 31570 246206
rect 233 245926 31799 246090
rect 430 245810 31570 245926
rect 233 245646 31799 245810
rect 430 245530 31570 245646
rect 233 245366 31799 245530
rect 430 245250 31570 245366
rect 233 245086 31799 245250
rect 430 244970 31570 245086
rect 233 244806 31799 244970
rect 430 244690 31570 244806
rect 233 244526 31799 244690
rect 430 244410 31570 244526
rect 233 244246 31799 244410
rect 430 244130 31570 244246
rect 233 243966 31799 244130
rect 430 243850 31570 243966
rect 233 243686 31799 243850
rect 430 243570 31570 243686
rect 233 243406 31799 243570
rect 430 243290 31570 243406
rect 233 243126 31799 243290
rect 430 243010 31570 243126
rect 233 242846 31799 243010
rect 430 242730 31570 242846
rect 233 242566 31799 242730
rect 430 242450 31570 242566
rect 233 242286 31799 242450
rect 430 242170 31570 242286
rect 233 242006 31799 242170
rect 430 241890 31570 242006
rect 233 241726 31799 241890
rect 430 241610 31570 241726
rect 233 241446 31799 241610
rect 430 241330 31570 241446
rect 233 241166 31799 241330
rect 430 241050 31570 241166
rect 233 240886 31799 241050
rect 430 240770 31570 240886
rect 233 240606 31799 240770
rect 430 240490 31570 240606
rect 233 240326 31799 240490
rect 430 240210 31570 240326
rect 233 240046 31799 240210
rect 430 239930 31570 240046
rect 233 239766 31799 239930
rect 430 239650 31570 239766
rect 233 239486 31799 239650
rect 430 239370 31570 239486
rect 233 239206 31799 239370
rect 430 239090 31570 239206
rect 233 238926 31799 239090
rect 430 238810 31570 238926
rect 233 238646 31799 238810
rect 430 238530 31570 238646
rect 233 238366 31799 238530
rect 430 238250 31570 238366
rect 233 238086 31799 238250
rect 430 237970 31570 238086
rect 233 237806 31799 237970
rect 430 237690 31570 237806
rect 233 237526 31799 237690
rect 430 237410 31570 237526
rect 233 237246 31799 237410
rect 430 237130 31570 237246
rect 233 236966 31799 237130
rect 430 236850 31570 236966
rect 233 236686 31799 236850
rect 430 236570 31570 236686
rect 233 236406 31799 236570
rect 430 236290 31570 236406
rect 233 236126 31799 236290
rect 430 236010 31570 236126
rect 233 235846 31799 236010
rect 430 235730 31570 235846
rect 233 235566 31799 235730
rect 430 235450 31570 235566
rect 233 235286 31799 235450
rect 430 235170 31570 235286
rect 233 235006 31799 235170
rect 430 234890 31570 235006
rect 233 234726 31799 234890
rect 430 234610 31570 234726
rect 233 234446 31799 234610
rect 430 234330 31570 234446
rect 233 234166 31799 234330
rect 430 234050 31570 234166
rect 233 233886 31799 234050
rect 430 233770 31570 233886
rect 233 233606 31799 233770
rect 430 233490 31570 233606
rect 233 233326 31799 233490
rect 430 233210 31570 233326
rect 233 233046 31799 233210
rect 430 232930 31570 233046
rect 233 232766 31799 232930
rect 430 232650 31570 232766
rect 233 232486 31799 232650
rect 430 232370 31570 232486
rect 233 232206 31799 232370
rect 430 232090 31570 232206
rect 233 231926 31799 232090
rect 430 231810 31570 231926
rect 233 231646 31799 231810
rect 430 231530 31570 231646
rect 233 231366 31799 231530
rect 430 231250 31570 231366
rect 233 231086 31799 231250
rect 430 230970 31570 231086
rect 233 230806 31799 230970
rect 430 230690 31570 230806
rect 233 230526 31799 230690
rect 430 230410 31570 230526
rect 233 230246 31799 230410
rect 430 230130 31570 230246
rect 233 229966 31799 230130
rect 430 229850 31570 229966
rect 233 229686 31799 229850
rect 430 229570 31570 229686
rect 233 229406 31799 229570
rect 430 229290 31570 229406
rect 233 229126 31799 229290
rect 430 229010 31570 229126
rect 233 228846 31799 229010
rect 430 228730 31570 228846
rect 233 228566 31799 228730
rect 430 228450 31570 228566
rect 233 228286 31799 228450
rect 430 228170 31570 228286
rect 233 228006 31799 228170
rect 430 227890 31570 228006
rect 233 227726 31799 227890
rect 430 227610 31570 227726
rect 233 227446 31799 227610
rect 430 227330 31570 227446
rect 233 227166 31799 227330
rect 430 227050 31570 227166
rect 233 226886 31799 227050
rect 430 226770 31570 226886
rect 233 226606 31799 226770
rect 430 226490 31570 226606
rect 233 226326 31799 226490
rect 430 226210 31570 226326
rect 233 226046 31799 226210
rect 430 225930 31570 226046
rect 233 225766 31799 225930
rect 430 225650 31570 225766
rect 233 225486 31799 225650
rect 430 225370 31570 225486
rect 233 225206 31799 225370
rect 430 225090 31570 225206
rect 233 224926 31799 225090
rect 430 224810 31570 224926
rect 233 224646 31799 224810
rect 430 224530 31570 224646
rect 233 224366 31799 224530
rect 430 224250 31570 224366
rect 233 224086 31799 224250
rect 430 223970 31570 224086
rect 233 223806 31799 223970
rect 430 223690 31570 223806
rect 233 223526 31799 223690
rect 430 223410 31570 223526
rect 233 223246 31799 223410
rect 430 223130 31570 223246
rect 233 222966 31799 223130
rect 430 222850 31570 222966
rect 233 222686 31799 222850
rect 430 222570 31570 222686
rect 233 222406 31799 222570
rect 430 222290 31570 222406
rect 233 222126 31799 222290
rect 430 222010 31570 222126
rect 233 221846 31799 222010
rect 430 221730 31570 221846
rect 233 221566 31799 221730
rect 430 221450 31570 221566
rect 233 221286 31799 221450
rect 430 221170 31570 221286
rect 233 221006 31799 221170
rect 430 220890 31570 221006
rect 233 220726 31799 220890
rect 430 220610 31570 220726
rect 233 220446 31799 220610
rect 430 220330 31570 220446
rect 233 220166 31799 220330
rect 430 220050 31570 220166
rect 233 219886 31799 220050
rect 430 219770 31570 219886
rect 233 219606 31799 219770
rect 430 219490 31570 219606
rect 233 219326 31799 219490
rect 430 219210 31570 219326
rect 233 219046 31799 219210
rect 430 218930 31570 219046
rect 233 218766 31799 218930
rect 430 218650 31570 218766
rect 233 218486 31799 218650
rect 430 218370 31570 218486
rect 233 218206 31799 218370
rect 430 218090 31570 218206
rect 233 217926 31799 218090
rect 430 217810 31570 217926
rect 233 217646 31799 217810
rect 430 217530 31570 217646
rect 233 217366 31799 217530
rect 430 217250 31570 217366
rect 233 217086 31799 217250
rect 430 216970 31570 217086
rect 233 216806 31799 216970
rect 430 216690 31570 216806
rect 233 216526 31799 216690
rect 430 216410 31570 216526
rect 233 216246 31799 216410
rect 430 216130 31570 216246
rect 233 215966 31799 216130
rect 430 215850 31570 215966
rect 233 215686 31799 215850
rect 430 215570 31570 215686
rect 233 215406 31799 215570
rect 430 215290 31570 215406
rect 233 215126 31799 215290
rect 430 215010 31570 215126
rect 233 214846 31799 215010
rect 430 214730 31570 214846
rect 233 214566 31799 214730
rect 430 214450 31570 214566
rect 233 214286 31799 214450
rect 430 214170 31570 214286
rect 233 214006 31799 214170
rect 430 213890 31570 214006
rect 233 213726 31799 213890
rect 430 213610 31570 213726
rect 233 213446 31799 213610
rect 430 213330 31570 213446
rect 233 213166 31799 213330
rect 430 213050 31570 213166
rect 233 212886 31799 213050
rect 430 212770 31570 212886
rect 233 212606 31799 212770
rect 430 212490 31570 212606
rect 233 212326 31799 212490
rect 430 212210 31570 212326
rect 233 212046 31799 212210
rect 430 211930 31570 212046
rect 233 211766 31799 211930
rect 430 211650 31570 211766
rect 233 211486 31799 211650
rect 430 211370 31570 211486
rect 233 211206 31799 211370
rect 430 211090 31570 211206
rect 233 210926 31799 211090
rect 430 210810 31570 210926
rect 233 210646 31799 210810
rect 430 210530 31570 210646
rect 233 210366 31799 210530
rect 430 210250 31570 210366
rect 233 210086 31799 210250
rect 430 209970 31570 210086
rect 233 209806 31799 209970
rect 430 209690 31570 209806
rect 233 209526 31799 209690
rect 430 209410 31570 209526
rect 233 209246 31799 209410
rect 430 209130 31570 209246
rect 233 208966 31799 209130
rect 430 208850 31570 208966
rect 233 208686 31799 208850
rect 430 208570 31570 208686
rect 233 208406 31799 208570
rect 430 208290 31570 208406
rect 233 208126 31799 208290
rect 430 208010 31570 208126
rect 233 207846 31799 208010
rect 430 207730 31570 207846
rect 233 207566 31799 207730
rect 430 207450 31570 207566
rect 233 207286 31799 207450
rect 430 207170 31570 207286
rect 233 207006 31799 207170
rect 430 206890 31570 207006
rect 233 206726 31799 206890
rect 430 206610 31570 206726
rect 233 206446 31799 206610
rect 430 206330 31570 206446
rect 233 206166 31799 206330
rect 430 206050 31570 206166
rect 233 205886 31799 206050
rect 430 205770 31570 205886
rect 233 205606 31799 205770
rect 430 205490 31570 205606
rect 233 205326 31799 205490
rect 430 205210 31570 205326
rect 233 205046 31799 205210
rect 430 204930 31570 205046
rect 233 204766 31799 204930
rect 430 204650 31570 204766
rect 233 204486 31799 204650
rect 430 204370 31570 204486
rect 233 204206 31799 204370
rect 430 204090 31570 204206
rect 233 203926 31799 204090
rect 430 203810 31570 203926
rect 233 203646 31799 203810
rect 430 203530 31570 203646
rect 233 203366 31799 203530
rect 430 203250 31570 203366
rect 233 203086 31799 203250
rect 430 202970 31570 203086
rect 233 202806 31799 202970
rect 430 202690 31570 202806
rect 233 202526 31799 202690
rect 430 202410 31570 202526
rect 233 202246 31799 202410
rect 430 202130 31570 202246
rect 233 201966 31799 202130
rect 430 201850 31570 201966
rect 233 201686 31799 201850
rect 430 201570 31570 201686
rect 233 201406 31799 201570
rect 430 201290 31570 201406
rect 233 201126 31799 201290
rect 430 201010 31570 201126
rect 233 200846 31799 201010
rect 430 200730 31570 200846
rect 233 200566 31799 200730
rect 430 200450 31570 200566
rect 233 200286 31799 200450
rect 430 200170 31570 200286
rect 233 200006 31799 200170
rect 430 199890 31570 200006
rect 233 199726 31799 199890
rect 430 199610 31570 199726
rect 233 199446 31799 199610
rect 430 199330 31570 199446
rect 233 199166 31799 199330
rect 430 199050 31570 199166
rect 233 198886 31799 199050
rect 430 198770 31570 198886
rect 233 198606 31799 198770
rect 430 198490 31570 198606
rect 233 198326 31799 198490
rect 430 198210 31570 198326
rect 233 198046 31799 198210
rect 430 197930 31570 198046
rect 233 197766 31799 197930
rect 430 197650 31570 197766
rect 233 197486 31799 197650
rect 430 197370 31570 197486
rect 233 197206 31799 197370
rect 430 197090 31570 197206
rect 233 196926 31799 197090
rect 430 196810 31570 196926
rect 233 196646 31799 196810
rect 430 196530 31570 196646
rect 233 196366 31799 196530
rect 430 196250 31570 196366
rect 233 196086 31799 196250
rect 430 195970 31570 196086
rect 233 195806 31799 195970
rect 430 195690 31570 195806
rect 233 195526 31799 195690
rect 430 195410 31570 195526
rect 233 195246 31799 195410
rect 430 195130 31570 195246
rect 233 194966 31799 195130
rect 430 194850 31570 194966
rect 233 194686 31799 194850
rect 430 194570 31570 194686
rect 233 194406 31799 194570
rect 430 194290 31570 194406
rect 233 194126 31799 194290
rect 430 194010 31570 194126
rect 233 193846 31799 194010
rect 430 193730 31570 193846
rect 233 193566 31799 193730
rect 430 193450 31570 193566
rect 233 193286 31799 193450
rect 430 193170 31570 193286
rect 233 193006 31799 193170
rect 430 192890 31570 193006
rect 233 192726 31799 192890
rect 430 192610 31570 192726
rect 233 192446 31799 192610
rect 430 192330 31570 192446
rect 233 192166 31799 192330
rect 430 192050 31570 192166
rect 233 191886 31799 192050
rect 430 191770 31570 191886
rect 233 191606 31799 191770
rect 430 191490 31570 191606
rect 233 191326 31799 191490
rect 430 191210 31570 191326
rect 233 191046 31799 191210
rect 430 190930 31570 191046
rect 233 190766 31799 190930
rect 430 190650 31570 190766
rect 233 190486 31799 190650
rect 430 190370 31570 190486
rect 233 190206 31799 190370
rect 430 190090 31570 190206
rect 233 189926 31799 190090
rect 430 189810 31570 189926
rect 233 189646 31799 189810
rect 430 189530 31570 189646
rect 233 189366 31799 189530
rect 430 189250 31570 189366
rect 233 189086 31799 189250
rect 430 188970 31570 189086
rect 233 188806 31799 188970
rect 430 188690 31570 188806
rect 233 188526 31799 188690
rect 430 188410 31570 188526
rect 233 188246 31799 188410
rect 430 188130 31570 188246
rect 233 187966 31799 188130
rect 430 187850 31570 187966
rect 233 187686 31799 187850
rect 430 187570 31570 187686
rect 233 187406 31799 187570
rect 430 187290 31570 187406
rect 233 187126 31799 187290
rect 430 187010 31570 187126
rect 233 186846 31799 187010
rect 430 186730 31570 186846
rect 233 186566 31799 186730
rect 430 186450 31570 186566
rect 233 186286 31799 186450
rect 430 186170 31570 186286
rect 233 186006 31799 186170
rect 430 185890 31570 186006
rect 233 185726 31799 185890
rect 430 185610 31570 185726
rect 233 185446 31799 185610
rect 430 185330 31570 185446
rect 233 185166 31799 185330
rect 430 185050 31570 185166
rect 233 184886 31799 185050
rect 430 184770 31570 184886
rect 233 184606 31799 184770
rect 430 184490 31570 184606
rect 233 184326 31799 184490
rect 430 184210 31570 184326
rect 233 184046 31799 184210
rect 430 183930 31570 184046
rect 233 183766 31799 183930
rect 430 183650 31570 183766
rect 233 183486 31799 183650
rect 430 183370 31570 183486
rect 233 183206 31799 183370
rect 430 183090 31570 183206
rect 233 182926 31799 183090
rect 430 182810 31570 182926
rect 233 182646 31799 182810
rect 430 182530 31570 182646
rect 233 182366 31799 182530
rect 430 182250 31570 182366
rect 233 182086 31799 182250
rect 430 181970 31570 182086
rect 233 181806 31799 181970
rect 430 181690 31570 181806
rect 233 181526 31799 181690
rect 430 181410 31570 181526
rect 233 181246 31799 181410
rect 430 181130 31570 181246
rect 233 180966 31799 181130
rect 430 180850 31570 180966
rect 233 180686 31799 180850
rect 430 180570 31570 180686
rect 233 180406 31799 180570
rect 430 180290 31570 180406
rect 233 180126 31799 180290
rect 430 180010 31570 180126
rect 233 179846 31799 180010
rect 430 179730 31570 179846
rect 233 179566 31799 179730
rect 430 179450 31570 179566
rect 233 179286 31799 179450
rect 430 179170 31570 179286
rect 233 179006 31799 179170
rect 430 178890 31570 179006
rect 233 178726 31799 178890
rect 430 178610 31570 178726
rect 233 178446 31799 178610
rect 430 178330 31570 178446
rect 233 178166 31799 178330
rect 430 178050 31570 178166
rect 233 177886 31799 178050
rect 430 177770 31570 177886
rect 233 177606 31799 177770
rect 430 177490 31570 177606
rect 233 177326 31799 177490
rect 430 177210 31570 177326
rect 233 177046 31799 177210
rect 430 176930 31570 177046
rect 233 176766 31799 176930
rect 430 176650 31570 176766
rect 233 176486 31799 176650
rect 430 176370 31570 176486
rect 233 176206 31799 176370
rect 430 176090 31570 176206
rect 233 175926 31799 176090
rect 430 175810 31570 175926
rect 233 175646 31799 175810
rect 430 175530 31570 175646
rect 233 175366 31799 175530
rect 430 175250 31570 175366
rect 233 175086 31799 175250
rect 430 174970 31570 175086
rect 233 174806 31799 174970
rect 430 174690 31570 174806
rect 233 174526 31799 174690
rect 430 174410 31570 174526
rect 233 174246 31799 174410
rect 430 174130 31570 174246
rect 233 173966 31799 174130
rect 430 173850 31570 173966
rect 233 173686 31799 173850
rect 430 173570 31570 173686
rect 233 173406 31799 173570
rect 430 173290 31570 173406
rect 233 173126 31799 173290
rect 430 173010 31570 173126
rect 233 172846 31799 173010
rect 430 172730 31570 172846
rect 233 172566 31799 172730
rect 430 172450 31570 172566
rect 233 172286 31799 172450
rect 430 172170 31570 172286
rect 233 172006 31799 172170
rect 430 171890 31570 172006
rect 233 171726 31799 171890
rect 430 171610 31570 171726
rect 233 171446 31799 171610
rect 430 171330 31570 171446
rect 233 171166 31799 171330
rect 430 171050 31570 171166
rect 233 170886 31799 171050
rect 430 170770 31570 170886
rect 233 170606 31799 170770
rect 430 170490 31570 170606
rect 233 170326 31799 170490
rect 430 170210 31570 170326
rect 233 170046 31799 170210
rect 430 169930 31570 170046
rect 233 169766 31799 169930
rect 430 169650 31570 169766
rect 233 169486 31799 169650
rect 430 169370 31570 169486
rect 233 169206 31799 169370
rect 430 169090 31570 169206
rect 233 168926 31799 169090
rect 430 168810 31570 168926
rect 233 168646 31799 168810
rect 430 168530 31570 168646
rect 233 168366 31799 168530
rect 430 168250 31570 168366
rect 233 168086 31799 168250
rect 430 167970 31570 168086
rect 233 167806 31799 167970
rect 430 167690 31570 167806
rect 233 167526 31799 167690
rect 430 167410 31570 167526
rect 233 167246 31799 167410
rect 430 167130 31570 167246
rect 233 166966 31799 167130
rect 430 166850 31570 166966
rect 233 166686 31799 166850
rect 430 166570 31570 166686
rect 233 166406 31799 166570
rect 430 166290 31570 166406
rect 233 166126 31799 166290
rect 430 166010 31570 166126
rect 233 165846 31799 166010
rect 430 165730 31570 165846
rect 233 165566 31799 165730
rect 430 165450 31570 165566
rect 233 165286 31799 165450
rect 430 165170 31570 165286
rect 233 165006 31799 165170
rect 430 164890 31570 165006
rect 233 164726 31799 164890
rect 430 164610 31570 164726
rect 233 164446 31799 164610
rect 430 164330 31570 164446
rect 233 164166 31799 164330
rect 430 164050 31570 164166
rect 233 163886 31799 164050
rect 430 163770 31570 163886
rect 233 163606 31799 163770
rect 430 163490 31570 163606
rect 233 163326 31799 163490
rect 430 163210 31570 163326
rect 233 163046 31799 163210
rect 430 162930 31570 163046
rect 233 162766 31799 162930
rect 430 162650 31570 162766
rect 233 162486 31799 162650
rect 430 162370 31570 162486
rect 233 162206 31799 162370
rect 430 162090 31570 162206
rect 233 161926 31799 162090
rect 430 161810 31570 161926
rect 233 161646 31799 161810
rect 430 161530 31570 161646
rect 233 161366 31799 161530
rect 430 161250 31570 161366
rect 233 161086 31799 161250
rect 430 160970 31570 161086
rect 233 160806 31799 160970
rect 430 160690 31570 160806
rect 233 160526 31799 160690
rect 430 160410 31570 160526
rect 233 160246 31799 160410
rect 430 160130 31570 160246
rect 233 159966 31799 160130
rect 430 159850 31570 159966
rect 233 159686 31799 159850
rect 430 159570 31570 159686
rect 233 159406 31799 159570
rect 430 159290 31570 159406
rect 233 159126 31799 159290
rect 430 159010 31570 159126
rect 233 158846 31799 159010
rect 430 158730 31570 158846
rect 233 158566 31799 158730
rect 430 158450 31570 158566
rect 233 158286 31799 158450
rect 430 158170 31570 158286
rect 233 158006 31799 158170
rect 430 157890 31570 158006
rect 233 157726 31799 157890
rect 430 157610 31570 157726
rect 233 157446 31799 157610
rect 430 157330 31570 157446
rect 233 157166 31799 157330
rect 430 157050 31570 157166
rect 233 156886 31799 157050
rect 430 156770 31570 156886
rect 233 156606 31799 156770
rect 430 156490 31570 156606
rect 233 156326 31799 156490
rect 430 156210 31570 156326
rect 233 156046 31799 156210
rect 430 155930 31570 156046
rect 233 155766 31799 155930
rect 430 155650 31570 155766
rect 233 155486 31799 155650
rect 430 155370 31570 155486
rect 233 155206 31799 155370
rect 430 155090 31570 155206
rect 233 154926 31799 155090
rect 430 154810 31570 154926
rect 233 154646 31799 154810
rect 430 154530 31570 154646
rect 233 154366 31799 154530
rect 430 154250 31570 154366
rect 233 154086 31799 154250
rect 430 153970 31570 154086
rect 233 153806 31799 153970
rect 430 153690 31570 153806
rect 233 153526 31799 153690
rect 430 153410 31570 153526
rect 233 153246 31799 153410
rect 430 153130 31570 153246
rect 233 152966 31799 153130
rect 430 152850 31570 152966
rect 233 152686 31799 152850
rect 430 152570 31570 152686
rect 233 152406 31799 152570
rect 430 152290 31570 152406
rect 233 152126 31799 152290
rect 430 152010 31570 152126
rect 233 151846 31799 152010
rect 430 151730 31570 151846
rect 233 151566 31799 151730
rect 430 151450 31570 151566
rect 233 151286 31799 151450
rect 430 151170 31570 151286
rect 233 151006 31799 151170
rect 430 150890 31570 151006
rect 233 150726 31799 150890
rect 430 150610 31570 150726
rect 233 150446 31799 150610
rect 430 150330 31570 150446
rect 233 150166 31799 150330
rect 430 150050 31570 150166
rect 233 149886 31799 150050
rect 430 149770 31570 149886
rect 233 149606 31799 149770
rect 430 149490 31570 149606
rect 233 149326 31799 149490
rect 430 149210 31570 149326
rect 233 149046 31799 149210
rect 430 148930 31570 149046
rect 233 148766 31799 148930
rect 430 148650 31570 148766
rect 233 148486 31799 148650
rect 430 148370 31570 148486
rect 233 148206 31799 148370
rect 430 148090 31570 148206
rect 233 147926 31799 148090
rect 430 147810 31570 147926
rect 233 147646 31799 147810
rect 430 147530 31570 147646
rect 233 147366 31799 147530
rect 430 147250 31570 147366
rect 233 147086 31799 147250
rect 430 146970 31570 147086
rect 233 146806 31799 146970
rect 430 146690 31570 146806
rect 233 146526 31799 146690
rect 430 146410 31570 146526
rect 233 146246 31799 146410
rect 430 146130 31570 146246
rect 233 145966 31799 146130
rect 430 145850 31570 145966
rect 233 145686 31799 145850
rect 430 145570 31570 145686
rect 233 145406 31799 145570
rect 430 145290 31570 145406
rect 233 145126 31799 145290
rect 430 145010 31570 145126
rect 233 144846 31799 145010
rect 430 144730 31570 144846
rect 233 144566 31799 144730
rect 430 144450 31570 144566
rect 233 144286 31799 144450
rect 430 144170 31570 144286
rect 233 144006 31799 144170
rect 430 143890 31570 144006
rect 233 143726 31799 143890
rect 430 143610 31570 143726
rect 233 143446 31799 143610
rect 430 143330 31570 143446
rect 233 143166 31799 143330
rect 430 143050 31570 143166
rect 233 142886 31799 143050
rect 430 142770 31570 142886
rect 233 142606 31799 142770
rect 430 142490 31570 142606
rect 233 142326 31799 142490
rect 430 142210 31570 142326
rect 233 142046 31799 142210
rect 430 141930 31570 142046
rect 233 141766 31799 141930
rect 430 141650 31570 141766
rect 233 141486 31799 141650
rect 430 141370 31570 141486
rect 233 141206 31799 141370
rect 430 141090 31570 141206
rect 233 140926 31799 141090
rect 430 140810 31570 140926
rect 233 140646 31799 140810
rect 430 140530 31570 140646
rect 233 140366 31799 140530
rect 430 140250 31570 140366
rect 233 140086 31799 140250
rect 430 139970 31570 140086
rect 233 139806 31799 139970
rect 430 139690 31570 139806
rect 233 139526 31799 139690
rect 430 139410 31570 139526
rect 233 139246 31799 139410
rect 430 139130 31570 139246
rect 233 138966 31799 139130
rect 430 138850 31570 138966
rect 233 138686 31799 138850
rect 430 138570 31570 138686
rect 233 138406 31799 138570
rect 430 138290 31570 138406
rect 233 138126 31799 138290
rect 430 138010 31570 138126
rect 233 137846 31799 138010
rect 430 137730 31570 137846
rect 233 137566 31799 137730
rect 430 137450 31570 137566
rect 233 137286 31799 137450
rect 430 137170 31570 137286
rect 233 137006 31799 137170
rect 430 136890 31570 137006
rect 233 136726 31799 136890
rect 430 136610 31570 136726
rect 233 136446 31799 136610
rect 430 136330 31570 136446
rect 233 136166 31799 136330
rect 430 136050 31570 136166
rect 233 135886 31799 136050
rect 430 135770 31570 135886
rect 233 135606 31799 135770
rect 430 135490 31570 135606
rect 233 135326 31799 135490
rect 430 135210 31570 135326
rect 233 135046 31799 135210
rect 430 134930 31570 135046
rect 233 134766 31799 134930
rect 430 134650 31570 134766
rect 233 134486 31799 134650
rect 430 134370 31570 134486
rect 233 134206 31799 134370
rect 430 134090 31570 134206
rect 233 133926 31799 134090
rect 430 133810 31570 133926
rect 233 133646 31799 133810
rect 430 133530 31570 133646
rect 233 133366 31799 133530
rect 430 133250 31570 133366
rect 233 133086 31799 133250
rect 430 132970 31570 133086
rect 233 132806 31799 132970
rect 430 132690 31570 132806
rect 233 132526 31799 132690
rect 430 132410 31570 132526
rect 233 132246 31799 132410
rect 430 132130 31570 132246
rect 233 131966 31799 132130
rect 430 131850 31570 131966
rect 233 131686 31799 131850
rect 430 131570 31570 131686
rect 233 131406 31799 131570
rect 430 131290 31570 131406
rect 233 131126 31799 131290
rect 430 131010 31570 131126
rect 233 130846 31799 131010
rect 430 130730 31570 130846
rect 233 130566 31799 130730
rect 430 130450 31570 130566
rect 233 130286 31799 130450
rect 430 130170 31570 130286
rect 233 130006 31799 130170
rect 430 129890 31570 130006
rect 233 129726 31799 129890
rect 430 129610 31570 129726
rect 233 129446 31799 129610
rect 430 129330 31570 129446
rect 233 129166 31799 129330
rect 430 129050 31570 129166
rect 233 128886 31799 129050
rect 430 128770 31570 128886
rect 233 128606 31799 128770
rect 430 128490 31570 128606
rect 233 128326 31799 128490
rect 430 128210 31570 128326
rect 233 128046 31799 128210
rect 430 127930 31570 128046
rect 233 127766 31799 127930
rect 430 127650 31570 127766
rect 233 127486 31799 127650
rect 430 127370 31570 127486
rect 233 127206 31799 127370
rect 430 127090 31570 127206
rect 233 126926 31799 127090
rect 430 126810 31570 126926
rect 233 126646 31799 126810
rect 430 126530 31570 126646
rect 233 126366 31799 126530
rect 430 126250 31570 126366
rect 233 126086 31799 126250
rect 430 125970 31570 126086
rect 233 125806 31799 125970
rect 430 125690 31570 125806
rect 233 125526 31799 125690
rect 430 125410 31570 125526
rect 233 125246 31799 125410
rect 430 125130 31570 125246
rect 233 124966 31799 125130
rect 430 124850 31570 124966
rect 233 124686 31799 124850
rect 430 124570 31570 124686
rect 233 124406 31799 124570
rect 430 124290 31570 124406
rect 233 124126 31799 124290
rect 430 124010 31570 124126
rect 233 123846 31799 124010
rect 430 123730 31570 123846
rect 233 123566 31799 123730
rect 430 123450 31570 123566
rect 233 123286 31799 123450
rect 430 123170 31570 123286
rect 233 123006 31799 123170
rect 430 122890 31570 123006
rect 233 122726 31799 122890
rect 430 122610 31570 122726
rect 233 122446 31799 122610
rect 430 122330 31570 122446
rect 233 122166 31799 122330
rect 430 122050 31570 122166
rect 233 121886 31799 122050
rect 430 121770 31570 121886
rect 233 121606 31799 121770
rect 430 121490 31570 121606
rect 233 121326 31799 121490
rect 430 121210 31570 121326
rect 233 121046 31799 121210
rect 430 120930 31570 121046
rect 233 120766 31799 120930
rect 430 120650 31570 120766
rect 233 120486 31799 120650
rect 430 120370 31570 120486
rect 233 120206 31799 120370
rect 430 120090 31570 120206
rect 233 119926 31799 120090
rect 430 119810 31570 119926
rect 233 119646 31799 119810
rect 430 119530 31570 119646
rect 233 119366 31799 119530
rect 430 119250 31570 119366
rect 233 119086 31799 119250
rect 430 118970 31570 119086
rect 233 118806 31799 118970
rect 430 118690 31570 118806
rect 233 118526 31799 118690
rect 430 118410 31570 118526
rect 233 118246 31799 118410
rect 430 118130 31570 118246
rect 233 117966 31799 118130
rect 430 117850 31570 117966
rect 233 117686 31799 117850
rect 430 117570 31570 117686
rect 233 117406 31799 117570
rect 430 117290 31570 117406
rect 233 117126 31799 117290
rect 430 117010 31570 117126
rect 233 116846 31799 117010
rect 430 116730 31570 116846
rect 233 116566 31799 116730
rect 430 116450 31570 116566
rect 233 116286 31799 116450
rect 430 116170 31570 116286
rect 233 116006 31799 116170
rect 430 115890 31570 116006
rect 233 115726 31799 115890
rect 430 115610 31570 115726
rect 233 115446 31799 115610
rect 430 115330 31570 115446
rect 233 115166 31799 115330
rect 430 115050 31570 115166
rect 233 114886 31799 115050
rect 430 114770 31570 114886
rect 233 114606 31799 114770
rect 430 114490 31570 114606
rect 233 114326 31799 114490
rect 430 114210 31570 114326
rect 233 114046 31799 114210
rect 430 113930 31570 114046
rect 233 113766 31799 113930
rect 430 113650 31570 113766
rect 233 113486 31799 113650
rect 430 113370 31570 113486
rect 233 113206 31799 113370
rect 430 113090 31570 113206
rect 233 112926 31799 113090
rect 430 112810 31570 112926
rect 233 112646 31799 112810
rect 430 112530 31570 112646
rect 233 112366 31799 112530
rect 430 112250 31570 112366
rect 233 112086 31799 112250
rect 430 111970 31570 112086
rect 233 111806 31799 111970
rect 430 111690 31570 111806
rect 233 111526 31799 111690
rect 430 111410 31570 111526
rect 233 111246 31799 111410
rect 430 111130 31570 111246
rect 233 110966 31799 111130
rect 430 110850 31570 110966
rect 233 110686 31799 110850
rect 430 110570 31570 110686
rect 233 110406 31799 110570
rect 430 110290 31570 110406
rect 233 110126 31799 110290
rect 430 110010 31570 110126
rect 233 109846 31799 110010
rect 430 109730 31570 109846
rect 233 109566 31799 109730
rect 430 109450 31570 109566
rect 233 109286 31799 109450
rect 430 109170 31570 109286
rect 233 109006 31799 109170
rect 430 108890 31570 109006
rect 233 108726 31799 108890
rect 430 108610 31570 108726
rect 233 108446 31799 108610
rect 430 108330 31570 108446
rect 233 108166 31799 108330
rect 430 108050 31570 108166
rect 233 107886 31799 108050
rect 430 107770 31570 107886
rect 233 107606 31799 107770
rect 430 107490 31570 107606
rect 233 107326 31799 107490
rect 430 107210 31570 107326
rect 233 107046 31799 107210
rect 430 106930 31570 107046
rect 233 106766 31799 106930
rect 430 106650 31570 106766
rect 233 106486 31799 106650
rect 430 106370 31570 106486
rect 233 106206 31799 106370
rect 430 106090 31570 106206
rect 233 105926 31799 106090
rect 430 105810 31570 105926
rect 233 105646 31799 105810
rect 430 105530 31570 105646
rect 233 105366 31799 105530
rect 430 105250 31570 105366
rect 233 105086 31799 105250
rect 430 104970 31570 105086
rect 233 104806 31799 104970
rect 430 104690 31570 104806
rect 233 104526 31799 104690
rect 430 104410 31570 104526
rect 233 104246 31799 104410
rect 430 104130 31570 104246
rect 233 103966 31799 104130
rect 430 103850 31570 103966
rect 233 103686 31799 103850
rect 430 103570 31570 103686
rect 233 103406 31799 103570
rect 430 103290 31570 103406
rect 233 103126 31799 103290
rect 430 103010 31570 103126
rect 233 102846 31799 103010
rect 430 102730 31570 102846
rect 233 102566 31799 102730
rect 430 102450 31570 102566
rect 233 102286 31799 102450
rect 430 102170 31570 102286
rect 233 102006 31799 102170
rect 430 101890 31570 102006
rect 233 101726 31799 101890
rect 430 101610 31570 101726
rect 233 101446 31799 101610
rect 430 101330 31570 101446
rect 233 101166 31799 101330
rect 430 101050 31570 101166
rect 233 100886 31799 101050
rect 430 100770 31570 100886
rect 233 100606 31799 100770
rect 430 100490 31570 100606
rect 233 100326 31799 100490
rect 430 100210 31570 100326
rect 233 100046 31799 100210
rect 430 99930 31570 100046
rect 233 99766 31799 99930
rect 430 99650 31570 99766
rect 233 99486 31799 99650
rect 430 99370 31570 99486
rect 233 99206 31799 99370
rect 430 99090 31570 99206
rect 233 98926 31799 99090
rect 430 98810 31570 98926
rect 233 98646 31799 98810
rect 430 98530 31570 98646
rect 233 98366 31799 98530
rect 430 98250 31570 98366
rect 233 98086 31799 98250
rect 430 97970 31570 98086
rect 233 97806 31799 97970
rect 430 97690 31570 97806
rect 233 97526 31799 97690
rect 430 97410 31570 97526
rect 233 97246 31799 97410
rect 430 97130 31570 97246
rect 233 96966 31799 97130
rect 430 96850 31570 96966
rect 233 96686 31799 96850
rect 430 96570 31570 96686
rect 233 96406 31799 96570
rect 430 96290 31570 96406
rect 233 96126 31799 96290
rect 430 96010 31570 96126
rect 233 95846 31799 96010
rect 430 95730 31570 95846
rect 233 95566 31799 95730
rect 430 95450 31570 95566
rect 233 95286 31799 95450
rect 430 95170 31570 95286
rect 233 95006 31799 95170
rect 430 94890 31570 95006
rect 233 94726 31799 94890
rect 430 94610 31570 94726
rect 233 94446 31799 94610
rect 430 94330 31570 94446
rect 233 94166 31799 94330
rect 430 94050 31570 94166
rect 233 93886 31799 94050
rect 430 93770 31570 93886
rect 233 93606 31799 93770
rect 430 93490 31570 93606
rect 233 93326 31799 93490
rect 430 93210 31570 93326
rect 233 93046 31799 93210
rect 430 92930 31570 93046
rect 233 92766 31799 92930
rect 430 92650 31570 92766
rect 233 92486 31799 92650
rect 430 92370 31570 92486
rect 233 92206 31799 92370
rect 430 92090 31570 92206
rect 233 91926 31799 92090
rect 430 91810 31570 91926
rect 233 91646 31799 91810
rect 430 91530 31570 91646
rect 233 91366 31799 91530
rect 430 91250 31570 91366
rect 233 91086 31799 91250
rect 430 90970 31570 91086
rect 233 90806 31799 90970
rect 430 90690 31570 90806
rect 233 90526 31799 90690
rect 430 90410 31570 90526
rect 233 90246 31799 90410
rect 430 90130 31570 90246
rect 233 89966 31799 90130
rect 430 89850 31570 89966
rect 233 89686 31799 89850
rect 430 89570 31570 89686
rect 233 89406 31799 89570
rect 430 89290 31570 89406
rect 233 89126 31799 89290
rect 430 89010 31570 89126
rect 233 88846 31799 89010
rect 430 88730 31570 88846
rect 233 88566 31799 88730
rect 430 88450 31570 88566
rect 233 88286 31799 88450
rect 430 88170 31570 88286
rect 233 88006 31799 88170
rect 430 87890 31570 88006
rect 233 87726 31799 87890
rect 430 87610 31570 87726
rect 233 87446 31799 87610
rect 430 87330 31570 87446
rect 233 87166 31799 87330
rect 430 87050 31570 87166
rect 233 86886 31799 87050
rect 430 86770 31570 86886
rect 233 86606 31799 86770
rect 430 86490 31570 86606
rect 233 86326 31799 86490
rect 430 86210 31570 86326
rect 233 86046 31799 86210
rect 430 85930 31570 86046
rect 233 85766 31799 85930
rect 430 85650 31570 85766
rect 233 85486 31799 85650
rect 430 85370 31570 85486
rect 233 85206 31799 85370
rect 430 85090 31570 85206
rect 233 84926 31799 85090
rect 430 84810 31570 84926
rect 233 84646 31799 84810
rect 430 84530 31570 84646
rect 233 84366 31799 84530
rect 430 84250 31570 84366
rect 233 84086 31799 84250
rect 430 83970 31570 84086
rect 233 83806 31799 83970
rect 430 83690 31570 83806
rect 233 83526 31799 83690
rect 430 83410 31570 83526
rect 233 83246 31799 83410
rect 430 83130 31570 83246
rect 233 82966 31799 83130
rect 430 82850 31570 82966
rect 233 82686 31799 82850
rect 430 82570 31570 82686
rect 233 82406 31799 82570
rect 430 82290 31570 82406
rect 233 82126 31799 82290
rect 430 82010 31570 82126
rect 233 81846 31799 82010
rect 430 81730 31570 81846
rect 233 81566 31799 81730
rect 430 81450 31570 81566
rect 233 81286 31799 81450
rect 430 81170 31570 81286
rect 233 81006 31799 81170
rect 430 80890 31570 81006
rect 233 80726 31799 80890
rect 430 80610 31570 80726
rect 233 80446 31799 80610
rect 430 80330 31570 80446
rect 233 80166 31799 80330
rect 430 80050 31570 80166
rect 233 79886 31799 80050
rect 430 79770 31570 79886
rect 233 79606 31799 79770
rect 430 79490 31570 79606
rect 233 79326 31799 79490
rect 430 79210 31570 79326
rect 233 79046 31799 79210
rect 430 78930 31570 79046
rect 233 78766 31799 78930
rect 430 78650 31570 78766
rect 233 78486 31799 78650
rect 430 78370 31570 78486
rect 233 78206 31799 78370
rect 430 78090 31570 78206
rect 233 77926 31799 78090
rect 430 77810 31570 77926
rect 233 77646 31799 77810
rect 430 77530 31570 77646
rect 233 77366 31799 77530
rect 430 77250 31570 77366
rect 233 77086 31799 77250
rect 430 76970 31570 77086
rect 233 76806 31799 76970
rect 430 76690 31570 76806
rect 233 76526 31799 76690
rect 430 76410 31570 76526
rect 233 76246 31799 76410
rect 430 76130 31570 76246
rect 233 75966 31799 76130
rect 430 75850 31570 75966
rect 233 75686 31799 75850
rect 430 75570 31570 75686
rect 233 75406 31799 75570
rect 430 75290 31570 75406
rect 233 75126 31799 75290
rect 430 75010 31570 75126
rect 233 74846 31799 75010
rect 430 74730 31570 74846
rect 233 74566 31799 74730
rect 430 74450 31570 74566
rect 233 74286 31799 74450
rect 430 74170 31570 74286
rect 233 74006 31799 74170
rect 430 73890 31570 74006
rect 233 73726 31799 73890
rect 430 73610 31570 73726
rect 233 73446 31799 73610
rect 430 73330 31570 73446
rect 233 73166 31799 73330
rect 430 73050 31570 73166
rect 233 72886 31799 73050
rect 430 72770 31570 72886
rect 233 72606 31799 72770
rect 430 72490 31570 72606
rect 233 72326 31799 72490
rect 430 72210 31570 72326
rect 233 72046 31799 72210
rect 430 71930 31570 72046
rect 233 71766 31799 71930
rect 430 71650 31570 71766
rect 233 71486 31799 71650
rect 430 71370 31570 71486
rect 233 71206 31799 71370
rect 430 71090 31570 71206
rect 233 70926 31799 71090
rect 430 70810 31570 70926
rect 233 70646 31799 70810
rect 430 70530 31570 70646
rect 233 70366 31799 70530
rect 430 70250 31570 70366
rect 233 70086 31799 70250
rect 430 69970 31570 70086
rect 233 69806 31799 69970
rect 430 69690 31570 69806
rect 233 69526 31799 69690
rect 430 69410 31570 69526
rect 233 69246 31799 69410
rect 430 69130 31570 69246
rect 233 68966 31799 69130
rect 430 68850 31570 68966
rect 233 68686 31799 68850
rect 430 68570 31570 68686
rect 233 68406 31799 68570
rect 430 68290 31570 68406
rect 233 68126 31799 68290
rect 430 68010 31570 68126
rect 233 67846 31799 68010
rect 430 67730 31570 67846
rect 233 67566 31799 67730
rect 430 67450 31570 67566
rect 233 67286 31799 67450
rect 430 67170 31570 67286
rect 233 67006 31799 67170
rect 430 66890 31570 67006
rect 233 66726 31799 66890
rect 430 66610 31570 66726
rect 233 66446 31799 66610
rect 430 66330 31570 66446
rect 233 66166 31799 66330
rect 430 66050 31570 66166
rect 233 65886 31799 66050
rect 430 65770 31570 65886
rect 233 65606 31799 65770
rect 430 65490 31570 65606
rect 233 65326 31799 65490
rect 430 65210 31570 65326
rect 233 65046 31799 65210
rect 430 64930 31570 65046
rect 233 64766 31799 64930
rect 430 64650 31570 64766
rect 233 64486 31799 64650
rect 430 64370 31570 64486
rect 233 64206 31799 64370
rect 430 64090 31570 64206
rect 233 63926 31799 64090
rect 430 63810 31570 63926
rect 233 63646 31799 63810
rect 430 63530 31570 63646
rect 233 63366 31799 63530
rect 430 63250 31570 63366
rect 233 63086 31799 63250
rect 430 62970 31570 63086
rect 233 62806 31799 62970
rect 430 62690 31570 62806
rect 233 62526 31799 62690
rect 430 62410 31570 62526
rect 233 62246 31799 62410
rect 430 62130 31570 62246
rect 233 61966 31799 62130
rect 430 61850 31570 61966
rect 233 61686 31799 61850
rect 430 61570 31570 61686
rect 233 61406 31799 61570
rect 430 61290 31570 61406
rect 233 61126 31799 61290
rect 430 61010 31570 61126
rect 233 60846 31799 61010
rect 430 60730 31570 60846
rect 233 60566 31799 60730
rect 430 60450 31570 60566
rect 233 60286 31799 60450
rect 430 60170 31570 60286
rect 233 60006 31799 60170
rect 430 59890 31570 60006
rect 233 59726 31799 59890
rect 430 59610 31570 59726
rect 233 59446 31799 59610
rect 430 59330 31570 59446
rect 233 59166 31799 59330
rect 430 59050 31570 59166
rect 233 58886 31799 59050
rect 430 58770 31570 58886
rect 233 58606 31799 58770
rect 430 58490 31570 58606
rect 233 58326 31799 58490
rect 430 58210 31570 58326
rect 233 58046 31799 58210
rect 430 57930 31570 58046
rect 233 57766 31799 57930
rect 430 57650 31570 57766
rect 233 57486 31799 57650
rect 430 57370 31570 57486
rect 233 57206 31799 57370
rect 430 57090 31570 57206
rect 233 56926 31799 57090
rect 430 56810 31570 56926
rect 233 56646 31799 56810
rect 430 56530 31570 56646
rect 233 56366 31799 56530
rect 430 56250 31570 56366
rect 233 56086 31799 56250
rect 430 55970 31570 56086
rect 233 55806 31799 55970
rect 430 55690 31570 55806
rect 233 55526 31799 55690
rect 430 55410 31570 55526
rect 233 55246 31799 55410
rect 430 55130 31570 55246
rect 233 54966 31799 55130
rect 430 54850 31570 54966
rect 233 54686 31799 54850
rect 430 54570 31570 54686
rect 233 54406 31799 54570
rect 430 54290 31570 54406
rect 233 54126 31799 54290
rect 430 54010 31570 54126
rect 233 53846 31799 54010
rect 430 53730 31570 53846
rect 233 53566 31799 53730
rect 430 53450 31570 53566
rect 233 53286 31799 53450
rect 430 53170 31570 53286
rect 233 53006 31799 53170
rect 430 52890 31570 53006
rect 233 52726 31799 52890
rect 430 52610 31570 52726
rect 233 52446 31799 52610
rect 430 52330 31570 52446
rect 233 52166 31799 52330
rect 430 52050 31570 52166
rect 233 51886 31799 52050
rect 430 51770 31570 51886
rect 233 51606 31799 51770
rect 430 51490 31570 51606
rect 233 51326 31799 51490
rect 430 51210 31570 51326
rect 233 51046 31799 51210
rect 430 50930 31570 51046
rect 233 50766 31799 50930
rect 430 50650 31570 50766
rect 233 50486 31799 50650
rect 430 50370 31570 50486
rect 233 50206 31799 50370
rect 430 50090 31570 50206
rect 233 49926 31799 50090
rect 430 49810 31570 49926
rect 233 49646 31799 49810
rect 430 49530 31570 49646
rect 233 49366 31799 49530
rect 430 49250 31570 49366
rect 233 49086 31799 49250
rect 430 48970 31570 49086
rect 233 48806 31799 48970
rect 430 48690 31570 48806
rect 233 48526 31799 48690
rect 430 48410 31570 48526
rect 233 48246 31799 48410
rect 430 48130 31570 48246
rect 233 47966 31799 48130
rect 430 47850 31570 47966
rect 233 47686 31799 47850
rect 430 47570 31570 47686
rect 233 47406 31799 47570
rect 430 47290 31570 47406
rect 233 47126 31799 47290
rect 430 47010 31570 47126
rect 233 46846 31799 47010
rect 430 46730 31570 46846
rect 233 46566 31799 46730
rect 430 46450 31570 46566
rect 233 46286 31799 46450
rect 430 46170 31570 46286
rect 233 46006 31799 46170
rect 430 45890 31570 46006
rect 233 45726 31799 45890
rect 430 45610 31570 45726
rect 233 45446 31799 45610
rect 430 45330 31570 45446
rect 233 45166 31799 45330
rect 430 45050 31570 45166
rect 233 44886 31799 45050
rect 430 44770 31570 44886
rect 233 44606 31799 44770
rect 430 44490 31570 44606
rect 233 44326 31799 44490
rect 430 44210 31570 44326
rect 233 44046 31799 44210
rect 430 43930 31570 44046
rect 233 43766 31799 43930
rect 430 43650 31570 43766
rect 233 43486 31799 43650
rect 430 43370 31570 43486
rect 233 43206 31799 43370
rect 430 43090 31570 43206
rect 233 42926 31799 43090
rect 430 42810 31570 42926
rect 233 42646 31799 42810
rect 430 42530 31570 42646
rect 233 42366 31799 42530
rect 430 42250 31570 42366
rect 233 42086 31799 42250
rect 430 41970 31570 42086
rect 233 41806 31799 41970
rect 430 41690 31570 41806
rect 233 41526 31799 41690
rect 430 41410 31570 41526
rect 233 41246 31799 41410
rect 430 41130 31570 41246
rect 233 40966 31799 41130
rect 430 40850 31570 40966
rect 233 40686 31799 40850
rect 430 40570 31570 40686
rect 233 40406 31799 40570
rect 430 40290 31570 40406
rect 233 40126 31799 40290
rect 430 40010 31570 40126
rect 233 39846 31799 40010
rect 430 39730 31570 39846
rect 233 39566 31799 39730
rect 430 39450 31570 39566
rect 233 39286 31799 39450
rect 430 39170 31570 39286
rect 233 39006 31799 39170
rect 430 38890 31570 39006
rect 233 38726 31799 38890
rect 430 38610 31570 38726
rect 233 38446 31799 38610
rect 430 38330 31570 38446
rect 233 38166 31799 38330
rect 430 38050 31570 38166
rect 233 37886 31799 38050
rect 430 37770 31570 37886
rect 233 37606 31799 37770
rect 430 37490 31570 37606
rect 233 37326 31799 37490
rect 430 37210 31570 37326
rect 233 37046 31799 37210
rect 430 36930 31570 37046
rect 233 36766 31799 36930
rect 430 36650 31570 36766
rect 233 36486 31799 36650
rect 430 36370 31570 36486
rect 233 36206 31799 36370
rect 430 36090 31570 36206
rect 233 35926 31799 36090
rect 430 35810 31570 35926
rect 233 35646 31799 35810
rect 430 35530 31570 35646
rect 233 35366 31799 35530
rect 430 35250 31570 35366
rect 233 35086 31799 35250
rect 430 34970 31570 35086
rect 233 34806 31799 34970
rect 430 34690 31570 34806
rect 233 34526 31799 34690
rect 430 34410 31570 34526
rect 233 34246 31799 34410
rect 430 34130 31570 34246
rect 233 33966 31799 34130
rect 430 33850 31570 33966
rect 233 33686 31799 33850
rect 430 33570 31570 33686
rect 233 33406 31799 33570
rect 430 33290 31570 33406
rect 233 33126 31799 33290
rect 430 33010 31570 33126
rect 233 32846 31799 33010
rect 430 32730 31570 32846
rect 233 32566 31799 32730
rect 430 32450 31570 32566
rect 233 32286 31799 32450
rect 430 32170 31570 32286
rect 233 32006 31799 32170
rect 430 31890 31570 32006
rect 233 31726 31799 31890
rect 430 31610 31570 31726
rect 233 31446 31799 31610
rect 430 31330 31570 31446
rect 233 31166 31799 31330
rect 430 31050 31570 31166
rect 233 30886 31799 31050
rect 430 30770 31570 30886
rect 233 30606 31799 30770
rect 430 30490 31570 30606
rect 233 30326 31799 30490
rect 430 30210 31570 30326
rect 233 30046 31799 30210
rect 430 29930 31570 30046
rect 233 29766 31799 29930
rect 430 29650 31570 29766
rect 233 29486 31799 29650
rect 430 29370 31570 29486
rect 233 29206 31799 29370
rect 430 29090 31570 29206
rect 233 28926 31799 29090
rect 430 28810 31570 28926
rect 233 28646 31799 28810
rect 430 28530 31570 28646
rect 233 28366 31799 28530
rect 430 28250 31570 28366
rect 233 28086 31799 28250
rect 430 27970 31570 28086
rect 233 27806 31799 27970
rect 430 27690 31570 27806
rect 233 27526 31799 27690
rect 430 27410 31570 27526
rect 233 27246 31799 27410
rect 430 27130 31570 27246
rect 233 26966 31799 27130
rect 430 26850 31570 26966
rect 233 26686 31799 26850
rect 430 26570 31570 26686
rect 233 26406 31799 26570
rect 430 26290 31570 26406
rect 233 26126 31799 26290
rect 430 26010 31570 26126
rect 233 25846 31799 26010
rect 430 25730 31570 25846
rect 233 25566 31799 25730
rect 430 25450 31570 25566
rect 233 25286 31799 25450
rect 430 25170 31570 25286
rect 233 25006 31799 25170
rect 430 24890 31570 25006
rect 233 24726 31799 24890
rect 430 24610 31570 24726
rect 233 24446 31799 24610
rect 430 24330 31570 24446
rect 233 24166 31799 24330
rect 430 24050 31570 24166
rect 233 23886 31799 24050
rect 430 23770 31570 23886
rect 233 23606 31799 23770
rect 430 23490 31570 23606
rect 233 23326 31799 23490
rect 430 23210 31570 23326
rect 233 23046 31799 23210
rect 430 22930 31570 23046
rect 233 22766 31799 22930
rect 430 22650 31570 22766
rect 233 22486 31799 22650
rect 430 22370 31570 22486
rect 233 22206 31799 22370
rect 430 22090 31570 22206
rect 233 21926 31799 22090
rect 430 21810 31570 21926
rect 233 21646 31799 21810
rect 430 21530 31570 21646
rect 233 21366 31799 21530
rect 430 21250 31570 21366
rect 233 21086 31799 21250
rect 430 20970 31570 21086
rect 233 20806 31799 20970
rect 430 20690 31570 20806
rect 233 20526 31799 20690
rect 430 20410 31570 20526
rect 233 20246 31799 20410
rect 430 20130 31570 20246
rect 233 19966 31799 20130
rect 430 19850 31570 19966
rect 233 19686 31799 19850
rect 430 19570 31570 19686
rect 233 19406 31799 19570
rect 430 19290 31570 19406
rect 233 19126 31799 19290
rect 430 19010 31570 19126
rect 233 18846 31799 19010
rect 430 18730 31570 18846
rect 233 18566 31799 18730
rect 430 18450 31570 18566
rect 233 1554 31799 18450
<< metal4 >>
rect 2224 1538 2384 268550
rect 9904 1538 10064 268550
rect 17584 1538 17744 268550
rect 25264 1538 25424 268550
<< obsm4 >>
rect 742 20505 2194 267951
rect 2414 20505 9874 267951
rect 10094 20505 17554 267951
rect 17774 20505 25234 267951
rect 25454 20505 31402 267951
<< labels >>
rlabel metal2 s 1008 0 1064 400 6 clk
port 1 nsew signal input
rlabel metal2 s 10640 269800 10696 270200 6 io_oeb[0]
port 2 nsew signal output
rlabel metal2 s 16240 269800 16296 270200 6 io_oeb[10]
port 3 nsew signal output
rlabel metal2 s 16800 269800 16856 270200 6 io_oeb[11]
port 4 nsew signal output
rlabel metal2 s 17360 269800 17416 270200 6 io_oeb[12]
port 5 nsew signal output
rlabel metal2 s 17920 269800 17976 270200 6 io_oeb[13]
port 6 nsew signal output
rlabel metal2 s 18480 269800 18536 270200 6 io_oeb[14]
port 7 nsew signal output
rlabel metal2 s 19040 269800 19096 270200 6 io_oeb[15]
port 8 nsew signal output
rlabel metal2 s 19600 269800 19656 270200 6 io_oeb[16]
port 9 nsew signal output
rlabel metal2 s 20160 269800 20216 270200 6 io_oeb[17]
port 10 nsew signal output
rlabel metal2 s 20720 269800 20776 270200 6 io_oeb[18]
port 11 nsew signal output
rlabel metal2 s 21280 269800 21336 270200 6 io_oeb[19]
port 12 nsew signal output
rlabel metal2 s 11200 269800 11256 270200 6 io_oeb[1]
port 13 nsew signal output
rlabel metal2 s 21840 269800 21896 270200 6 io_oeb[20]
port 14 nsew signal output
rlabel metal2 s 22400 269800 22456 270200 6 io_oeb[21]
port 15 nsew signal output
rlabel metal2 s 22960 269800 23016 270200 6 io_oeb[22]
port 16 nsew signal output
rlabel metal2 s 23520 269800 23576 270200 6 io_oeb[23]
port 17 nsew signal output
rlabel metal2 s 24080 269800 24136 270200 6 io_oeb[24]
port 18 nsew signal output
rlabel metal2 s 24640 269800 24696 270200 6 io_oeb[25]
port 19 nsew signal output
rlabel metal2 s 25200 269800 25256 270200 6 io_oeb[26]
port 20 nsew signal output
rlabel metal2 s 25760 269800 25816 270200 6 io_oeb[27]
port 21 nsew signal output
rlabel metal2 s 26320 269800 26376 270200 6 io_oeb[28]
port 22 nsew signal output
rlabel metal2 s 26880 269800 26936 270200 6 io_oeb[29]
port 23 nsew signal output
rlabel metal2 s 11760 269800 11816 270200 6 io_oeb[2]
port 24 nsew signal output
rlabel metal2 s 27440 269800 27496 270200 6 io_oeb[30]
port 25 nsew signal output
rlabel metal2 s 28000 269800 28056 270200 6 io_oeb[31]
port 26 nsew signal output
rlabel metal2 s 28560 269800 28616 270200 6 io_oeb[32]
port 27 nsew signal output
rlabel metal2 s 29120 269800 29176 270200 6 io_oeb[33]
port 28 nsew signal output
rlabel metal2 s 29680 269800 29736 270200 6 io_oeb[34]
port 29 nsew signal output
rlabel metal2 s 30240 269800 30296 270200 6 io_oeb[35]
port 30 nsew signal output
rlabel metal2 s 30800 269800 30856 270200 6 io_oeb[36]
port 31 nsew signal output
rlabel metal2 s 31360 269800 31416 270200 6 io_oeb[37]
port 32 nsew signal output
rlabel metal2 s 12320 269800 12376 270200 6 io_oeb[3]
port 33 nsew signal output
rlabel metal2 s 12880 269800 12936 270200 6 io_oeb[4]
port 34 nsew signal output
rlabel metal2 s 13440 269800 13496 270200 6 io_oeb[5]
port 35 nsew signal output
rlabel metal2 s 14000 269800 14056 270200 6 io_oeb[6]
port 36 nsew signal output
rlabel metal2 s 14560 269800 14616 270200 6 io_oeb[7]
port 37 nsew signal output
rlabel metal2 s 15120 269800 15176 270200 6 io_oeb[8]
port 38 nsew signal output
rlabel metal2 s 15680 269800 15736 270200 6 io_oeb[9]
port 39 nsew signal output
rlabel metal3 s 0 31920 400 31976 6 itasegm[0]
port 40 nsew signal input
rlabel metal3 s 31600 44240 32000 44296 6 itasegm[100]
port 41 nsew signal input
rlabel metal3 s 31600 44520 32000 44576 6 itasegm[101]
port 42 nsew signal input
rlabel metal3 s 31600 44800 32000 44856 6 itasegm[102]
port 43 nsew signal input
rlabel metal3 s 31600 45080 32000 45136 6 itasegm[103]
port 44 nsew signal input
rlabel metal3 s 31600 45360 32000 45416 6 itasegm[104]
port 45 nsew signal input
rlabel metal3 s 31600 45640 32000 45696 6 itasegm[105]
port 46 nsew signal input
rlabel metal3 s 31600 45920 32000 45976 6 itasegm[106]
port 47 nsew signal input
rlabel metal3 s 31600 46200 32000 46256 6 itasegm[107]
port 48 nsew signal input
rlabel metal3 s 31600 46480 32000 46536 6 itasegm[108]
port 49 nsew signal input
rlabel metal3 s 31600 46760 32000 46816 6 itasegm[109]
port 50 nsew signal input
rlabel metal3 s 0 34720 400 34776 6 itasegm[10]
port 51 nsew signal input
rlabel metal3 s 31600 47040 32000 47096 6 itasegm[110]
port 52 nsew signal input
rlabel metal3 s 31600 47320 32000 47376 6 itasegm[111]
port 53 nsew signal input
rlabel metal3 s 0 61040 400 61096 6 itasegm[112]
port 54 nsew signal input
rlabel metal3 s 0 61320 400 61376 6 itasegm[113]
port 55 nsew signal input
rlabel metal3 s 0 61600 400 61656 6 itasegm[114]
port 56 nsew signal input
rlabel metal3 s 0 61880 400 61936 6 itasegm[115]
port 57 nsew signal input
rlabel metal3 s 0 62160 400 62216 6 itasegm[116]
port 58 nsew signal input
rlabel metal3 s 0 62440 400 62496 6 itasegm[117]
port 59 nsew signal input
rlabel metal3 s 0 62720 400 62776 6 itasegm[118]
port 60 nsew signal input
rlabel metal3 s 0 63000 400 63056 6 itasegm[119]
port 61 nsew signal input
rlabel metal3 s 0 35000 400 35056 6 itasegm[11]
port 62 nsew signal input
rlabel metal3 s 0 63280 400 63336 6 itasegm[120]
port 63 nsew signal input
rlabel metal3 s 0 63560 400 63616 6 itasegm[121]
port 64 nsew signal input
rlabel metal3 s 0 63840 400 63896 6 itasegm[122]
port 65 nsew signal input
rlabel metal3 s 0 64120 400 64176 6 itasegm[123]
port 66 nsew signal input
rlabel metal3 s 0 64400 400 64456 6 itasegm[124]
port 67 nsew signal input
rlabel metal3 s 0 64680 400 64736 6 itasegm[125]
port 68 nsew signal input
rlabel metal3 s 0 64960 400 65016 6 itasegm[126]
port 69 nsew signal input
rlabel metal3 s 0 65240 400 65296 6 itasegm[127]
port 70 nsew signal input
rlabel metal3 s 0 65520 400 65576 6 itasegm[128]
port 71 nsew signal input
rlabel metal3 s 0 65800 400 65856 6 itasegm[129]
port 72 nsew signal input
rlabel metal3 s 0 35280 400 35336 6 itasegm[12]
port 73 nsew signal input
rlabel metal3 s 0 66080 400 66136 6 itasegm[130]
port 74 nsew signal input
rlabel metal3 s 0 66360 400 66416 6 itasegm[131]
port 75 nsew signal input
rlabel metal3 s 0 66640 400 66696 6 itasegm[132]
port 76 nsew signal input
rlabel metal3 s 0 66920 400 66976 6 itasegm[133]
port 77 nsew signal input
rlabel metal3 s 0 67200 400 67256 6 itasegm[134]
port 78 nsew signal input
rlabel metal3 s 0 67480 400 67536 6 itasegm[135]
port 79 nsew signal input
rlabel metal3 s 0 67760 400 67816 6 itasegm[136]
port 80 nsew signal input
rlabel metal3 s 0 68040 400 68096 6 itasegm[137]
port 81 nsew signal input
rlabel metal3 s 0 68320 400 68376 6 itasegm[138]
port 82 nsew signal input
rlabel metal3 s 0 68600 400 68656 6 itasegm[139]
port 83 nsew signal input
rlabel metal3 s 0 35560 400 35616 6 itasegm[13]
port 84 nsew signal input
rlabel metal3 s 0 68880 400 68936 6 itasegm[140]
port 85 nsew signal input
rlabel metal3 s 0 69160 400 69216 6 itasegm[141]
port 86 nsew signal input
rlabel metal3 s 0 69440 400 69496 6 itasegm[142]
port 87 nsew signal input
rlabel metal3 s 0 69720 400 69776 6 itasegm[143]
port 88 nsew signal input
rlabel metal3 s 0 70000 400 70056 6 itasegm[144]
port 89 nsew signal input
rlabel metal3 s 0 70280 400 70336 6 itasegm[145]
port 90 nsew signal input
rlabel metal3 s 0 70560 400 70616 6 itasegm[146]
port 91 nsew signal input
rlabel metal3 s 0 70840 400 70896 6 itasegm[147]
port 92 nsew signal input
rlabel metal3 s 0 71120 400 71176 6 itasegm[148]
port 93 nsew signal input
rlabel metal3 s 0 71400 400 71456 6 itasegm[149]
port 94 nsew signal input
rlabel metal3 s 0 35840 400 35896 6 itasegm[14]
port 95 nsew signal input
rlabel metal3 s 0 71680 400 71736 6 itasegm[150]
port 96 nsew signal input
rlabel metal3 s 0 71960 400 72016 6 itasegm[151]
port 97 nsew signal input
rlabel metal3 s 0 72240 400 72296 6 itasegm[152]
port 98 nsew signal input
rlabel metal3 s 0 72520 400 72576 6 itasegm[153]
port 99 nsew signal input
rlabel metal3 s 0 72800 400 72856 6 itasegm[154]
port 100 nsew signal input
rlabel metal3 s 0 73080 400 73136 6 itasegm[155]
port 101 nsew signal input
rlabel metal3 s 0 73360 400 73416 6 itasegm[156]
port 102 nsew signal input
rlabel metal3 s 0 73640 400 73696 6 itasegm[157]
port 103 nsew signal input
rlabel metal3 s 0 73920 400 73976 6 itasegm[158]
port 104 nsew signal input
rlabel metal3 s 0 74200 400 74256 6 itasegm[159]
port 105 nsew signal input
rlabel metal3 s 0 36120 400 36176 6 itasegm[15]
port 106 nsew signal input
rlabel metal3 s 0 74480 400 74536 6 itasegm[160]
port 107 nsew signal input
rlabel metal3 s 0 74760 400 74816 6 itasegm[161]
port 108 nsew signal input
rlabel metal3 s 0 75040 400 75096 6 itasegm[162]
port 109 nsew signal input
rlabel metal3 s 0 75320 400 75376 6 itasegm[163]
port 110 nsew signal input
rlabel metal3 s 0 75600 400 75656 6 itasegm[164]
port 111 nsew signal input
rlabel metal3 s 0 75880 400 75936 6 itasegm[165]
port 112 nsew signal input
rlabel metal3 s 0 76160 400 76216 6 itasegm[166]
port 113 nsew signal input
rlabel metal3 s 0 76440 400 76496 6 itasegm[167]
port 114 nsew signal input
rlabel metal3 s 31600 61040 32000 61096 6 itasegm[168]
port 115 nsew signal input
rlabel metal3 s 31600 61320 32000 61376 6 itasegm[169]
port 116 nsew signal input
rlabel metal3 s 0 36400 400 36456 6 itasegm[16]
port 117 nsew signal input
rlabel metal3 s 31600 61600 32000 61656 6 itasegm[170]
port 118 nsew signal input
rlabel metal3 s 31600 61880 32000 61936 6 itasegm[171]
port 119 nsew signal input
rlabel metal3 s 31600 62160 32000 62216 6 itasegm[172]
port 120 nsew signal input
rlabel metal3 s 31600 62440 32000 62496 6 itasegm[173]
port 121 nsew signal input
rlabel metal3 s 31600 62720 32000 62776 6 itasegm[174]
port 122 nsew signal input
rlabel metal3 s 31600 63000 32000 63056 6 itasegm[175]
port 123 nsew signal input
rlabel metal3 s 31600 63280 32000 63336 6 itasegm[176]
port 124 nsew signal input
rlabel metal3 s 31600 63560 32000 63616 6 itasegm[177]
port 125 nsew signal input
rlabel metal3 s 31600 63840 32000 63896 6 itasegm[178]
port 126 nsew signal input
rlabel metal3 s 31600 64120 32000 64176 6 itasegm[179]
port 127 nsew signal input
rlabel metal3 s 0 36680 400 36736 6 itasegm[17]
port 128 nsew signal input
rlabel metal3 s 31600 64400 32000 64456 6 itasegm[180]
port 129 nsew signal input
rlabel metal3 s 31600 64680 32000 64736 6 itasegm[181]
port 130 nsew signal input
rlabel metal3 s 31600 64960 32000 65016 6 itasegm[182]
port 131 nsew signal input
rlabel metal3 s 31600 65240 32000 65296 6 itasegm[183]
port 132 nsew signal input
rlabel metal3 s 31600 65520 32000 65576 6 itasegm[184]
port 133 nsew signal input
rlabel metal3 s 31600 65800 32000 65856 6 itasegm[185]
port 134 nsew signal input
rlabel metal3 s 31600 66080 32000 66136 6 itasegm[186]
port 135 nsew signal input
rlabel metal3 s 31600 66360 32000 66416 6 itasegm[187]
port 136 nsew signal input
rlabel metal3 s 31600 66640 32000 66696 6 itasegm[188]
port 137 nsew signal input
rlabel metal3 s 31600 66920 32000 66976 6 itasegm[189]
port 138 nsew signal input
rlabel metal3 s 0 36960 400 37016 6 itasegm[18]
port 139 nsew signal input
rlabel metal3 s 31600 67200 32000 67256 6 itasegm[190]
port 140 nsew signal input
rlabel metal3 s 31600 67480 32000 67536 6 itasegm[191]
port 141 nsew signal input
rlabel metal3 s 31600 67760 32000 67816 6 itasegm[192]
port 142 nsew signal input
rlabel metal3 s 31600 68040 32000 68096 6 itasegm[193]
port 143 nsew signal input
rlabel metal3 s 31600 68320 32000 68376 6 itasegm[194]
port 144 nsew signal input
rlabel metal3 s 31600 68600 32000 68656 6 itasegm[195]
port 145 nsew signal input
rlabel metal3 s 31600 68880 32000 68936 6 itasegm[196]
port 146 nsew signal input
rlabel metal3 s 31600 69160 32000 69216 6 itasegm[197]
port 147 nsew signal input
rlabel metal3 s 31600 69440 32000 69496 6 itasegm[198]
port 148 nsew signal input
rlabel metal3 s 31600 69720 32000 69776 6 itasegm[199]
port 149 nsew signal input
rlabel metal3 s 0 37240 400 37296 6 itasegm[19]
port 150 nsew signal input
rlabel metal3 s 0 32200 400 32256 6 itasegm[1]
port 151 nsew signal input
rlabel metal3 s 31600 70000 32000 70056 6 itasegm[200]
port 152 nsew signal input
rlabel metal3 s 31600 70280 32000 70336 6 itasegm[201]
port 153 nsew signal input
rlabel metal3 s 31600 70560 32000 70616 6 itasegm[202]
port 154 nsew signal input
rlabel metal3 s 31600 70840 32000 70896 6 itasegm[203]
port 155 nsew signal input
rlabel metal3 s 31600 71120 32000 71176 6 itasegm[204]
port 156 nsew signal input
rlabel metal3 s 31600 71400 32000 71456 6 itasegm[205]
port 157 nsew signal input
rlabel metal3 s 31600 71680 32000 71736 6 itasegm[206]
port 158 nsew signal input
rlabel metal3 s 31600 71960 32000 72016 6 itasegm[207]
port 159 nsew signal input
rlabel metal3 s 31600 72240 32000 72296 6 itasegm[208]
port 160 nsew signal input
rlabel metal3 s 31600 72520 32000 72576 6 itasegm[209]
port 161 nsew signal input
rlabel metal3 s 0 37520 400 37576 6 itasegm[20]
port 162 nsew signal input
rlabel metal3 s 31600 72800 32000 72856 6 itasegm[210]
port 163 nsew signal input
rlabel metal3 s 31600 73080 32000 73136 6 itasegm[211]
port 164 nsew signal input
rlabel metal3 s 31600 73360 32000 73416 6 itasegm[212]
port 165 nsew signal input
rlabel metal3 s 31600 73640 32000 73696 6 itasegm[213]
port 166 nsew signal input
rlabel metal3 s 31600 73920 32000 73976 6 itasegm[214]
port 167 nsew signal input
rlabel metal3 s 31600 74200 32000 74256 6 itasegm[215]
port 168 nsew signal input
rlabel metal3 s 31600 74480 32000 74536 6 itasegm[216]
port 169 nsew signal input
rlabel metal3 s 31600 74760 32000 74816 6 itasegm[217]
port 170 nsew signal input
rlabel metal3 s 31600 75040 32000 75096 6 itasegm[218]
port 171 nsew signal input
rlabel metal3 s 31600 75320 32000 75376 6 itasegm[219]
port 172 nsew signal input
rlabel metal3 s 0 37800 400 37856 6 itasegm[21]
port 173 nsew signal input
rlabel metal3 s 31600 75600 32000 75656 6 itasegm[220]
port 174 nsew signal input
rlabel metal3 s 31600 75880 32000 75936 6 itasegm[221]
port 175 nsew signal input
rlabel metal3 s 31600 76160 32000 76216 6 itasegm[222]
port 176 nsew signal input
rlabel metal3 s 31600 76440 32000 76496 6 itasegm[223]
port 177 nsew signal input
rlabel metal3 s 0 90160 400 90216 6 itasegm[224]
port 178 nsew signal input
rlabel metal3 s 0 90440 400 90496 6 itasegm[225]
port 179 nsew signal input
rlabel metal3 s 0 90720 400 90776 6 itasegm[226]
port 180 nsew signal input
rlabel metal3 s 0 91000 400 91056 6 itasegm[227]
port 181 nsew signal input
rlabel metal3 s 0 91280 400 91336 6 itasegm[228]
port 182 nsew signal input
rlabel metal3 s 0 91560 400 91616 6 itasegm[229]
port 183 nsew signal input
rlabel metal3 s 0 38080 400 38136 6 itasegm[22]
port 184 nsew signal input
rlabel metal3 s 0 91840 400 91896 6 itasegm[230]
port 185 nsew signal input
rlabel metal3 s 0 92120 400 92176 6 itasegm[231]
port 186 nsew signal input
rlabel metal3 s 0 92400 400 92456 6 itasegm[232]
port 187 nsew signal input
rlabel metal3 s 0 92680 400 92736 6 itasegm[233]
port 188 nsew signal input
rlabel metal3 s 0 92960 400 93016 6 itasegm[234]
port 189 nsew signal input
rlabel metal3 s 0 93240 400 93296 6 itasegm[235]
port 190 nsew signal input
rlabel metal3 s 0 93520 400 93576 6 itasegm[236]
port 191 nsew signal input
rlabel metal3 s 0 93800 400 93856 6 itasegm[237]
port 192 nsew signal input
rlabel metal3 s 0 94080 400 94136 6 itasegm[238]
port 193 nsew signal input
rlabel metal3 s 0 94360 400 94416 6 itasegm[239]
port 194 nsew signal input
rlabel metal3 s 0 38360 400 38416 6 itasegm[23]
port 195 nsew signal input
rlabel metal3 s 0 94640 400 94696 6 itasegm[240]
port 196 nsew signal input
rlabel metal3 s 0 94920 400 94976 6 itasegm[241]
port 197 nsew signal input
rlabel metal3 s 0 95200 400 95256 6 itasegm[242]
port 198 nsew signal input
rlabel metal3 s 0 95480 400 95536 6 itasegm[243]
port 199 nsew signal input
rlabel metal3 s 0 95760 400 95816 6 itasegm[244]
port 200 nsew signal input
rlabel metal3 s 0 96040 400 96096 6 itasegm[245]
port 201 nsew signal input
rlabel metal3 s 0 96320 400 96376 6 itasegm[246]
port 202 nsew signal input
rlabel metal3 s 0 96600 400 96656 6 itasegm[247]
port 203 nsew signal input
rlabel metal3 s 0 96880 400 96936 6 itasegm[248]
port 204 nsew signal input
rlabel metal3 s 0 97160 400 97216 6 itasegm[249]
port 205 nsew signal input
rlabel metal3 s 0 38640 400 38696 6 itasegm[24]
port 206 nsew signal input
rlabel metal3 s 0 97440 400 97496 6 itasegm[250]
port 207 nsew signal input
rlabel metal3 s 0 97720 400 97776 6 itasegm[251]
port 208 nsew signal input
rlabel metal3 s 0 98000 400 98056 6 itasegm[252]
port 209 nsew signal input
rlabel metal3 s 0 98280 400 98336 6 itasegm[253]
port 210 nsew signal input
rlabel metal3 s 0 98560 400 98616 6 itasegm[254]
port 211 nsew signal input
rlabel metal3 s 0 98840 400 98896 6 itasegm[255]
port 212 nsew signal input
rlabel metal3 s 0 99120 400 99176 6 itasegm[256]
port 213 nsew signal input
rlabel metal3 s 0 99400 400 99456 6 itasegm[257]
port 214 nsew signal input
rlabel metal3 s 0 99680 400 99736 6 itasegm[258]
port 215 nsew signal input
rlabel metal3 s 0 99960 400 100016 6 itasegm[259]
port 216 nsew signal input
rlabel metal3 s 0 38920 400 38976 6 itasegm[25]
port 217 nsew signal input
rlabel metal3 s 0 100240 400 100296 6 itasegm[260]
port 218 nsew signal input
rlabel metal3 s 0 100520 400 100576 6 itasegm[261]
port 219 nsew signal input
rlabel metal3 s 0 100800 400 100856 6 itasegm[262]
port 220 nsew signal input
rlabel metal3 s 0 101080 400 101136 6 itasegm[263]
port 221 nsew signal input
rlabel metal3 s 0 101360 400 101416 6 itasegm[264]
port 222 nsew signal input
rlabel metal3 s 0 101640 400 101696 6 itasegm[265]
port 223 nsew signal input
rlabel metal3 s 0 101920 400 101976 6 itasegm[266]
port 224 nsew signal input
rlabel metal3 s 0 102200 400 102256 6 itasegm[267]
port 225 nsew signal input
rlabel metal3 s 0 102480 400 102536 6 itasegm[268]
port 226 nsew signal input
rlabel metal3 s 0 102760 400 102816 6 itasegm[269]
port 227 nsew signal input
rlabel metal3 s 0 39200 400 39256 6 itasegm[26]
port 228 nsew signal input
rlabel metal3 s 0 103040 400 103096 6 itasegm[270]
port 229 nsew signal input
rlabel metal3 s 0 103320 400 103376 6 itasegm[271]
port 230 nsew signal input
rlabel metal3 s 0 103600 400 103656 6 itasegm[272]
port 231 nsew signal input
rlabel metal3 s 0 103880 400 103936 6 itasegm[273]
port 232 nsew signal input
rlabel metal3 s 0 104160 400 104216 6 itasegm[274]
port 233 nsew signal input
rlabel metal3 s 0 104440 400 104496 6 itasegm[275]
port 234 nsew signal input
rlabel metal3 s 0 104720 400 104776 6 itasegm[276]
port 235 nsew signal input
rlabel metal3 s 0 105000 400 105056 6 itasegm[277]
port 236 nsew signal input
rlabel metal3 s 0 105280 400 105336 6 itasegm[278]
port 237 nsew signal input
rlabel metal3 s 0 105560 400 105616 6 itasegm[279]
port 238 nsew signal input
rlabel metal3 s 0 39480 400 39536 6 itasegm[27]
port 239 nsew signal input
rlabel metal3 s 31600 90160 32000 90216 6 itasegm[280]
port 240 nsew signal input
rlabel metal3 s 31600 90440 32000 90496 6 itasegm[281]
port 241 nsew signal input
rlabel metal3 s 31600 90720 32000 90776 6 itasegm[282]
port 242 nsew signal input
rlabel metal3 s 31600 91000 32000 91056 6 itasegm[283]
port 243 nsew signal input
rlabel metal3 s 31600 91280 32000 91336 6 itasegm[284]
port 244 nsew signal input
rlabel metal3 s 31600 91560 32000 91616 6 itasegm[285]
port 245 nsew signal input
rlabel metal3 s 31600 91840 32000 91896 6 itasegm[286]
port 246 nsew signal input
rlabel metal3 s 31600 92120 32000 92176 6 itasegm[287]
port 247 nsew signal input
rlabel metal3 s 31600 92400 32000 92456 6 itasegm[288]
port 248 nsew signal input
rlabel metal3 s 31600 92680 32000 92736 6 itasegm[289]
port 249 nsew signal input
rlabel metal3 s 0 39760 400 39816 6 itasegm[28]
port 250 nsew signal input
rlabel metal3 s 31600 92960 32000 93016 6 itasegm[290]
port 251 nsew signal input
rlabel metal3 s 31600 93240 32000 93296 6 itasegm[291]
port 252 nsew signal input
rlabel metal3 s 31600 93520 32000 93576 6 itasegm[292]
port 253 nsew signal input
rlabel metal3 s 31600 93800 32000 93856 6 itasegm[293]
port 254 nsew signal input
rlabel metal3 s 31600 94080 32000 94136 6 itasegm[294]
port 255 nsew signal input
rlabel metal3 s 31600 94360 32000 94416 6 itasegm[295]
port 256 nsew signal input
rlabel metal3 s 31600 94640 32000 94696 6 itasegm[296]
port 257 nsew signal input
rlabel metal3 s 31600 94920 32000 94976 6 itasegm[297]
port 258 nsew signal input
rlabel metal3 s 31600 95200 32000 95256 6 itasegm[298]
port 259 nsew signal input
rlabel metal3 s 31600 95480 32000 95536 6 itasegm[299]
port 260 nsew signal input
rlabel metal3 s 0 40040 400 40096 6 itasegm[29]
port 261 nsew signal input
rlabel metal3 s 0 32480 400 32536 6 itasegm[2]
port 262 nsew signal input
rlabel metal3 s 31600 95760 32000 95816 6 itasegm[300]
port 263 nsew signal input
rlabel metal3 s 31600 96040 32000 96096 6 itasegm[301]
port 264 nsew signal input
rlabel metal3 s 31600 96320 32000 96376 6 itasegm[302]
port 265 nsew signal input
rlabel metal3 s 31600 96600 32000 96656 6 itasegm[303]
port 266 nsew signal input
rlabel metal3 s 31600 96880 32000 96936 6 itasegm[304]
port 267 nsew signal input
rlabel metal3 s 31600 97160 32000 97216 6 itasegm[305]
port 268 nsew signal input
rlabel metal3 s 31600 97440 32000 97496 6 itasegm[306]
port 269 nsew signal input
rlabel metal3 s 31600 97720 32000 97776 6 itasegm[307]
port 270 nsew signal input
rlabel metal3 s 31600 98000 32000 98056 6 itasegm[308]
port 271 nsew signal input
rlabel metal3 s 31600 98280 32000 98336 6 itasegm[309]
port 272 nsew signal input
rlabel metal3 s 0 40320 400 40376 6 itasegm[30]
port 273 nsew signal input
rlabel metal3 s 31600 98560 32000 98616 6 itasegm[310]
port 274 nsew signal input
rlabel metal3 s 31600 98840 32000 98896 6 itasegm[311]
port 275 nsew signal input
rlabel metal3 s 31600 99120 32000 99176 6 itasegm[312]
port 276 nsew signal input
rlabel metal3 s 31600 99400 32000 99456 6 itasegm[313]
port 277 nsew signal input
rlabel metal3 s 31600 99680 32000 99736 6 itasegm[314]
port 278 nsew signal input
rlabel metal3 s 31600 99960 32000 100016 6 itasegm[315]
port 279 nsew signal input
rlabel metal3 s 31600 100240 32000 100296 6 itasegm[316]
port 280 nsew signal input
rlabel metal3 s 31600 100520 32000 100576 6 itasegm[317]
port 281 nsew signal input
rlabel metal3 s 31600 100800 32000 100856 6 itasegm[318]
port 282 nsew signal input
rlabel metal3 s 31600 101080 32000 101136 6 itasegm[319]
port 283 nsew signal input
rlabel metal3 s 0 40600 400 40656 6 itasegm[31]
port 284 nsew signal input
rlabel metal3 s 31600 101360 32000 101416 6 itasegm[320]
port 285 nsew signal input
rlabel metal3 s 31600 101640 32000 101696 6 itasegm[321]
port 286 nsew signal input
rlabel metal3 s 31600 101920 32000 101976 6 itasegm[322]
port 287 nsew signal input
rlabel metal3 s 31600 102200 32000 102256 6 itasegm[323]
port 288 nsew signal input
rlabel metal3 s 31600 102480 32000 102536 6 itasegm[324]
port 289 nsew signal input
rlabel metal3 s 31600 102760 32000 102816 6 itasegm[325]
port 290 nsew signal input
rlabel metal3 s 31600 103040 32000 103096 6 itasegm[326]
port 291 nsew signal input
rlabel metal3 s 31600 103320 32000 103376 6 itasegm[327]
port 292 nsew signal input
rlabel metal3 s 31600 103600 32000 103656 6 itasegm[328]
port 293 nsew signal input
rlabel metal3 s 31600 103880 32000 103936 6 itasegm[329]
port 294 nsew signal input
rlabel metal3 s 0 40880 400 40936 6 itasegm[32]
port 295 nsew signal input
rlabel metal3 s 31600 104160 32000 104216 6 itasegm[330]
port 296 nsew signal input
rlabel metal3 s 31600 104440 32000 104496 6 itasegm[331]
port 297 nsew signal input
rlabel metal3 s 31600 104720 32000 104776 6 itasegm[332]
port 298 nsew signal input
rlabel metal3 s 31600 105000 32000 105056 6 itasegm[333]
port 299 nsew signal input
rlabel metal3 s 31600 105280 32000 105336 6 itasegm[334]
port 300 nsew signal input
rlabel metal3 s 31600 105560 32000 105616 6 itasegm[335]
port 301 nsew signal input
rlabel metal3 s 0 119280 400 119336 6 itasegm[336]
port 302 nsew signal input
rlabel metal3 s 0 119560 400 119616 6 itasegm[337]
port 303 nsew signal input
rlabel metal3 s 0 119840 400 119896 6 itasegm[338]
port 304 nsew signal input
rlabel metal3 s 0 120120 400 120176 6 itasegm[339]
port 305 nsew signal input
rlabel metal3 s 0 41160 400 41216 6 itasegm[33]
port 306 nsew signal input
rlabel metal3 s 0 120400 400 120456 6 itasegm[340]
port 307 nsew signal input
rlabel metal3 s 0 120680 400 120736 6 itasegm[341]
port 308 nsew signal input
rlabel metal3 s 0 120960 400 121016 6 itasegm[342]
port 309 nsew signal input
rlabel metal3 s 0 121240 400 121296 6 itasegm[343]
port 310 nsew signal input
rlabel metal3 s 0 121520 400 121576 6 itasegm[344]
port 311 nsew signal input
rlabel metal3 s 0 121800 400 121856 6 itasegm[345]
port 312 nsew signal input
rlabel metal3 s 0 122080 400 122136 6 itasegm[346]
port 313 nsew signal input
rlabel metal3 s 0 122360 400 122416 6 itasegm[347]
port 314 nsew signal input
rlabel metal3 s 0 122640 400 122696 6 itasegm[348]
port 315 nsew signal input
rlabel metal3 s 0 122920 400 122976 6 itasegm[349]
port 316 nsew signal input
rlabel metal3 s 0 41440 400 41496 6 itasegm[34]
port 317 nsew signal input
rlabel metal3 s 0 123200 400 123256 6 itasegm[350]
port 318 nsew signal input
rlabel metal3 s 0 123480 400 123536 6 itasegm[351]
port 319 nsew signal input
rlabel metal3 s 0 123760 400 123816 6 itasegm[352]
port 320 nsew signal input
rlabel metal3 s 0 124040 400 124096 6 itasegm[353]
port 321 nsew signal input
rlabel metal3 s 0 124320 400 124376 6 itasegm[354]
port 322 nsew signal input
rlabel metal3 s 0 124600 400 124656 6 itasegm[355]
port 323 nsew signal input
rlabel metal3 s 0 124880 400 124936 6 itasegm[356]
port 324 nsew signal input
rlabel metal3 s 0 125160 400 125216 6 itasegm[357]
port 325 nsew signal input
rlabel metal3 s 0 125440 400 125496 6 itasegm[358]
port 326 nsew signal input
rlabel metal3 s 0 125720 400 125776 6 itasegm[359]
port 327 nsew signal input
rlabel metal3 s 0 41720 400 41776 6 itasegm[35]
port 328 nsew signal input
rlabel metal3 s 0 126000 400 126056 6 itasegm[360]
port 329 nsew signal input
rlabel metal3 s 0 126280 400 126336 6 itasegm[361]
port 330 nsew signal input
rlabel metal3 s 0 126560 400 126616 6 itasegm[362]
port 331 nsew signal input
rlabel metal3 s 0 126840 400 126896 6 itasegm[363]
port 332 nsew signal input
rlabel metal3 s 0 127120 400 127176 6 itasegm[364]
port 333 nsew signal input
rlabel metal3 s 0 127400 400 127456 6 itasegm[365]
port 334 nsew signal input
rlabel metal3 s 0 127680 400 127736 6 itasegm[366]
port 335 nsew signal input
rlabel metal3 s 0 127960 400 128016 6 itasegm[367]
port 336 nsew signal input
rlabel metal3 s 0 128240 400 128296 6 itasegm[368]
port 337 nsew signal input
rlabel metal3 s 0 128520 400 128576 6 itasegm[369]
port 338 nsew signal input
rlabel metal3 s 0 42000 400 42056 6 itasegm[36]
port 339 nsew signal input
rlabel metal3 s 0 128800 400 128856 6 itasegm[370]
port 340 nsew signal input
rlabel metal3 s 0 129080 400 129136 6 itasegm[371]
port 341 nsew signal input
rlabel metal3 s 0 129360 400 129416 6 itasegm[372]
port 342 nsew signal input
rlabel metal3 s 0 129640 400 129696 6 itasegm[373]
port 343 nsew signal input
rlabel metal3 s 0 129920 400 129976 6 itasegm[374]
port 344 nsew signal input
rlabel metal3 s 0 130200 400 130256 6 itasegm[375]
port 345 nsew signal input
rlabel metal3 s 0 130480 400 130536 6 itasegm[376]
port 346 nsew signal input
rlabel metal3 s 0 130760 400 130816 6 itasegm[377]
port 347 nsew signal input
rlabel metal3 s 0 131040 400 131096 6 itasegm[378]
port 348 nsew signal input
rlabel metal3 s 0 131320 400 131376 6 itasegm[379]
port 349 nsew signal input
rlabel metal3 s 0 42280 400 42336 6 itasegm[37]
port 350 nsew signal input
rlabel metal3 s 0 131600 400 131656 6 itasegm[380]
port 351 nsew signal input
rlabel metal3 s 0 131880 400 131936 6 itasegm[381]
port 352 nsew signal input
rlabel metal3 s 0 132160 400 132216 6 itasegm[382]
port 353 nsew signal input
rlabel metal3 s 0 132440 400 132496 6 itasegm[383]
port 354 nsew signal input
rlabel metal3 s 0 132720 400 132776 6 itasegm[384]
port 355 nsew signal input
rlabel metal3 s 0 133000 400 133056 6 itasegm[385]
port 356 nsew signal input
rlabel metal3 s 0 133280 400 133336 6 itasegm[386]
port 357 nsew signal input
rlabel metal3 s 0 133560 400 133616 6 itasegm[387]
port 358 nsew signal input
rlabel metal3 s 0 133840 400 133896 6 itasegm[388]
port 359 nsew signal input
rlabel metal3 s 0 134120 400 134176 6 itasegm[389]
port 360 nsew signal input
rlabel metal3 s 0 42560 400 42616 6 itasegm[38]
port 361 nsew signal input
rlabel metal3 s 0 134400 400 134456 6 itasegm[390]
port 362 nsew signal input
rlabel metal3 s 0 134680 400 134736 6 itasegm[391]
port 363 nsew signal input
rlabel metal3 s 31600 119280 32000 119336 6 itasegm[392]
port 364 nsew signal input
rlabel metal3 s 31600 119560 32000 119616 6 itasegm[393]
port 365 nsew signal input
rlabel metal3 s 31600 119840 32000 119896 6 itasegm[394]
port 366 nsew signal input
rlabel metal3 s 31600 120120 32000 120176 6 itasegm[395]
port 367 nsew signal input
rlabel metal3 s 31600 120400 32000 120456 6 itasegm[396]
port 368 nsew signal input
rlabel metal3 s 31600 120680 32000 120736 6 itasegm[397]
port 369 nsew signal input
rlabel metal3 s 31600 120960 32000 121016 6 itasegm[398]
port 370 nsew signal input
rlabel metal3 s 31600 121240 32000 121296 6 itasegm[399]
port 371 nsew signal input
rlabel metal3 s 0 42840 400 42896 6 itasegm[39]
port 372 nsew signal input
rlabel metal3 s 0 32760 400 32816 6 itasegm[3]
port 373 nsew signal input
rlabel metal3 s 31600 121520 32000 121576 6 itasegm[400]
port 374 nsew signal input
rlabel metal3 s 31600 121800 32000 121856 6 itasegm[401]
port 375 nsew signal input
rlabel metal3 s 31600 122080 32000 122136 6 itasegm[402]
port 376 nsew signal input
rlabel metal3 s 31600 122360 32000 122416 6 itasegm[403]
port 377 nsew signal input
rlabel metal3 s 31600 122640 32000 122696 6 itasegm[404]
port 378 nsew signal input
rlabel metal3 s 31600 122920 32000 122976 6 itasegm[405]
port 379 nsew signal input
rlabel metal3 s 31600 123200 32000 123256 6 itasegm[406]
port 380 nsew signal input
rlabel metal3 s 31600 123480 32000 123536 6 itasegm[407]
port 381 nsew signal input
rlabel metal3 s 31600 123760 32000 123816 6 itasegm[408]
port 382 nsew signal input
rlabel metal3 s 31600 124040 32000 124096 6 itasegm[409]
port 383 nsew signal input
rlabel metal3 s 0 43120 400 43176 6 itasegm[40]
port 384 nsew signal input
rlabel metal3 s 31600 124320 32000 124376 6 itasegm[410]
port 385 nsew signal input
rlabel metal3 s 31600 124600 32000 124656 6 itasegm[411]
port 386 nsew signal input
rlabel metal3 s 31600 124880 32000 124936 6 itasegm[412]
port 387 nsew signal input
rlabel metal3 s 31600 125160 32000 125216 6 itasegm[413]
port 388 nsew signal input
rlabel metal3 s 31600 125440 32000 125496 6 itasegm[414]
port 389 nsew signal input
rlabel metal3 s 31600 125720 32000 125776 6 itasegm[415]
port 390 nsew signal input
rlabel metal3 s 31600 126000 32000 126056 6 itasegm[416]
port 391 nsew signal input
rlabel metal3 s 31600 126280 32000 126336 6 itasegm[417]
port 392 nsew signal input
rlabel metal3 s 31600 126560 32000 126616 6 itasegm[418]
port 393 nsew signal input
rlabel metal3 s 31600 126840 32000 126896 6 itasegm[419]
port 394 nsew signal input
rlabel metal3 s 0 43400 400 43456 6 itasegm[41]
port 395 nsew signal input
rlabel metal3 s 31600 127120 32000 127176 6 itasegm[420]
port 396 nsew signal input
rlabel metal3 s 31600 127400 32000 127456 6 itasegm[421]
port 397 nsew signal input
rlabel metal3 s 31600 127680 32000 127736 6 itasegm[422]
port 398 nsew signal input
rlabel metal3 s 31600 127960 32000 128016 6 itasegm[423]
port 399 nsew signal input
rlabel metal3 s 31600 128240 32000 128296 6 itasegm[424]
port 400 nsew signal input
rlabel metal3 s 31600 128520 32000 128576 6 itasegm[425]
port 401 nsew signal input
rlabel metal3 s 31600 128800 32000 128856 6 itasegm[426]
port 402 nsew signal input
rlabel metal3 s 31600 129080 32000 129136 6 itasegm[427]
port 403 nsew signal input
rlabel metal3 s 31600 129360 32000 129416 6 itasegm[428]
port 404 nsew signal input
rlabel metal3 s 31600 129640 32000 129696 6 itasegm[429]
port 405 nsew signal input
rlabel metal3 s 0 43680 400 43736 6 itasegm[42]
port 406 nsew signal input
rlabel metal3 s 31600 129920 32000 129976 6 itasegm[430]
port 407 nsew signal input
rlabel metal3 s 31600 130200 32000 130256 6 itasegm[431]
port 408 nsew signal input
rlabel metal3 s 31600 130480 32000 130536 6 itasegm[432]
port 409 nsew signal input
rlabel metal3 s 31600 130760 32000 130816 6 itasegm[433]
port 410 nsew signal input
rlabel metal3 s 31600 131040 32000 131096 6 itasegm[434]
port 411 nsew signal input
rlabel metal3 s 31600 131320 32000 131376 6 itasegm[435]
port 412 nsew signal input
rlabel metal3 s 31600 131600 32000 131656 6 itasegm[436]
port 413 nsew signal input
rlabel metal3 s 31600 131880 32000 131936 6 itasegm[437]
port 414 nsew signal input
rlabel metal3 s 31600 132160 32000 132216 6 itasegm[438]
port 415 nsew signal input
rlabel metal3 s 31600 132440 32000 132496 6 itasegm[439]
port 416 nsew signal input
rlabel metal3 s 0 43960 400 44016 6 itasegm[43]
port 417 nsew signal input
rlabel metal3 s 31600 132720 32000 132776 6 itasegm[440]
port 418 nsew signal input
rlabel metal3 s 31600 133000 32000 133056 6 itasegm[441]
port 419 nsew signal input
rlabel metal3 s 31600 133280 32000 133336 6 itasegm[442]
port 420 nsew signal input
rlabel metal3 s 31600 133560 32000 133616 6 itasegm[443]
port 421 nsew signal input
rlabel metal3 s 31600 133840 32000 133896 6 itasegm[444]
port 422 nsew signal input
rlabel metal3 s 31600 134120 32000 134176 6 itasegm[445]
port 423 nsew signal input
rlabel metal3 s 31600 134400 32000 134456 6 itasegm[446]
port 424 nsew signal input
rlabel metal3 s 31600 134680 32000 134736 6 itasegm[447]
port 425 nsew signal input
rlabel metal3 s 0 148400 400 148456 6 itasegm[448]
port 426 nsew signal input
rlabel metal3 s 0 148680 400 148736 6 itasegm[449]
port 427 nsew signal input
rlabel metal3 s 0 44240 400 44296 6 itasegm[44]
port 428 nsew signal input
rlabel metal3 s 0 148960 400 149016 6 itasegm[450]
port 429 nsew signal input
rlabel metal3 s 0 149240 400 149296 6 itasegm[451]
port 430 nsew signal input
rlabel metal3 s 0 149520 400 149576 6 itasegm[452]
port 431 nsew signal input
rlabel metal3 s 0 149800 400 149856 6 itasegm[453]
port 432 nsew signal input
rlabel metal3 s 0 150080 400 150136 6 itasegm[454]
port 433 nsew signal input
rlabel metal3 s 0 150360 400 150416 6 itasegm[455]
port 434 nsew signal input
rlabel metal3 s 0 150640 400 150696 6 itasegm[456]
port 435 nsew signal input
rlabel metal3 s 0 150920 400 150976 6 itasegm[457]
port 436 nsew signal input
rlabel metal3 s 0 151200 400 151256 6 itasegm[458]
port 437 nsew signal input
rlabel metal3 s 0 151480 400 151536 6 itasegm[459]
port 438 nsew signal input
rlabel metal3 s 0 44520 400 44576 6 itasegm[45]
port 439 nsew signal input
rlabel metal3 s 0 151760 400 151816 6 itasegm[460]
port 440 nsew signal input
rlabel metal3 s 0 152040 400 152096 6 itasegm[461]
port 441 nsew signal input
rlabel metal3 s 0 152320 400 152376 6 itasegm[462]
port 442 nsew signal input
rlabel metal3 s 0 152600 400 152656 6 itasegm[463]
port 443 nsew signal input
rlabel metal3 s 0 152880 400 152936 6 itasegm[464]
port 444 nsew signal input
rlabel metal3 s 0 153160 400 153216 6 itasegm[465]
port 445 nsew signal input
rlabel metal3 s 0 153440 400 153496 6 itasegm[466]
port 446 nsew signal input
rlabel metal3 s 0 153720 400 153776 6 itasegm[467]
port 447 nsew signal input
rlabel metal3 s 0 154000 400 154056 6 itasegm[468]
port 448 nsew signal input
rlabel metal3 s 0 154280 400 154336 6 itasegm[469]
port 449 nsew signal input
rlabel metal3 s 0 44800 400 44856 6 itasegm[46]
port 450 nsew signal input
rlabel metal3 s 0 154560 400 154616 6 itasegm[470]
port 451 nsew signal input
rlabel metal3 s 0 154840 400 154896 6 itasegm[471]
port 452 nsew signal input
rlabel metal3 s 0 155120 400 155176 6 itasegm[472]
port 453 nsew signal input
rlabel metal3 s 0 155400 400 155456 6 itasegm[473]
port 454 nsew signal input
rlabel metal3 s 0 155680 400 155736 6 itasegm[474]
port 455 nsew signal input
rlabel metal3 s 0 155960 400 156016 6 itasegm[475]
port 456 nsew signal input
rlabel metal3 s 0 156240 400 156296 6 itasegm[476]
port 457 nsew signal input
rlabel metal3 s 0 156520 400 156576 6 itasegm[477]
port 458 nsew signal input
rlabel metal3 s 0 156800 400 156856 6 itasegm[478]
port 459 nsew signal input
rlabel metal3 s 0 157080 400 157136 6 itasegm[479]
port 460 nsew signal input
rlabel metal3 s 0 45080 400 45136 6 itasegm[47]
port 461 nsew signal input
rlabel metal3 s 0 157360 400 157416 6 itasegm[480]
port 462 nsew signal input
rlabel metal3 s 0 157640 400 157696 6 itasegm[481]
port 463 nsew signal input
rlabel metal3 s 0 157920 400 157976 6 itasegm[482]
port 464 nsew signal input
rlabel metal3 s 0 158200 400 158256 6 itasegm[483]
port 465 nsew signal input
rlabel metal3 s 0 158480 400 158536 6 itasegm[484]
port 466 nsew signal input
rlabel metal3 s 0 158760 400 158816 6 itasegm[485]
port 467 nsew signal input
rlabel metal3 s 0 159040 400 159096 6 itasegm[486]
port 468 nsew signal input
rlabel metal3 s 0 159320 400 159376 6 itasegm[487]
port 469 nsew signal input
rlabel metal3 s 0 159600 400 159656 6 itasegm[488]
port 470 nsew signal input
rlabel metal3 s 0 159880 400 159936 6 itasegm[489]
port 471 nsew signal input
rlabel metal3 s 0 45360 400 45416 6 itasegm[48]
port 472 nsew signal input
rlabel metal3 s 0 160160 400 160216 6 itasegm[490]
port 473 nsew signal input
rlabel metal3 s 0 160440 400 160496 6 itasegm[491]
port 474 nsew signal input
rlabel metal3 s 0 160720 400 160776 6 itasegm[492]
port 475 nsew signal input
rlabel metal3 s 0 161000 400 161056 6 itasegm[493]
port 476 nsew signal input
rlabel metal3 s 0 161280 400 161336 6 itasegm[494]
port 477 nsew signal input
rlabel metal3 s 0 161560 400 161616 6 itasegm[495]
port 478 nsew signal input
rlabel metal3 s 0 161840 400 161896 6 itasegm[496]
port 479 nsew signal input
rlabel metal3 s 0 162120 400 162176 6 itasegm[497]
port 480 nsew signal input
rlabel metal3 s 0 162400 400 162456 6 itasegm[498]
port 481 nsew signal input
rlabel metal3 s 0 162680 400 162736 6 itasegm[499]
port 482 nsew signal input
rlabel metal3 s 0 45640 400 45696 6 itasegm[49]
port 483 nsew signal input
rlabel metal3 s 0 33040 400 33096 6 itasegm[4]
port 484 nsew signal input
rlabel metal3 s 0 162960 400 163016 6 itasegm[500]
port 485 nsew signal input
rlabel metal3 s 0 163240 400 163296 6 itasegm[501]
port 486 nsew signal input
rlabel metal3 s 0 163520 400 163576 6 itasegm[502]
port 487 nsew signal input
rlabel metal3 s 0 163800 400 163856 6 itasegm[503]
port 488 nsew signal input
rlabel metal3 s 31600 148400 32000 148456 6 itasegm[504]
port 489 nsew signal input
rlabel metal3 s 31600 148680 32000 148736 6 itasegm[505]
port 490 nsew signal input
rlabel metal3 s 31600 148960 32000 149016 6 itasegm[506]
port 491 nsew signal input
rlabel metal3 s 31600 149240 32000 149296 6 itasegm[507]
port 492 nsew signal input
rlabel metal3 s 31600 149520 32000 149576 6 itasegm[508]
port 493 nsew signal input
rlabel metal3 s 31600 149800 32000 149856 6 itasegm[509]
port 494 nsew signal input
rlabel metal3 s 0 45920 400 45976 6 itasegm[50]
port 495 nsew signal input
rlabel metal3 s 31600 150080 32000 150136 6 itasegm[510]
port 496 nsew signal input
rlabel metal3 s 31600 150360 32000 150416 6 itasegm[511]
port 497 nsew signal input
rlabel metal3 s 31600 150640 32000 150696 6 itasegm[512]
port 498 nsew signal input
rlabel metal3 s 31600 150920 32000 150976 6 itasegm[513]
port 499 nsew signal input
rlabel metal3 s 31600 151200 32000 151256 6 itasegm[514]
port 500 nsew signal input
rlabel metal3 s 31600 151480 32000 151536 6 itasegm[515]
port 501 nsew signal input
rlabel metal3 s 31600 151760 32000 151816 6 itasegm[516]
port 502 nsew signal input
rlabel metal3 s 31600 152040 32000 152096 6 itasegm[517]
port 503 nsew signal input
rlabel metal3 s 31600 152320 32000 152376 6 itasegm[518]
port 504 nsew signal input
rlabel metal3 s 31600 152600 32000 152656 6 itasegm[519]
port 505 nsew signal input
rlabel metal3 s 0 46200 400 46256 6 itasegm[51]
port 506 nsew signal input
rlabel metal3 s 31600 152880 32000 152936 6 itasegm[520]
port 507 nsew signal input
rlabel metal3 s 31600 153160 32000 153216 6 itasegm[521]
port 508 nsew signal input
rlabel metal3 s 31600 153440 32000 153496 6 itasegm[522]
port 509 nsew signal input
rlabel metal3 s 31600 153720 32000 153776 6 itasegm[523]
port 510 nsew signal input
rlabel metal3 s 31600 154000 32000 154056 6 itasegm[524]
port 511 nsew signal input
rlabel metal3 s 31600 154280 32000 154336 6 itasegm[525]
port 512 nsew signal input
rlabel metal3 s 31600 154560 32000 154616 6 itasegm[526]
port 513 nsew signal input
rlabel metal3 s 31600 154840 32000 154896 6 itasegm[527]
port 514 nsew signal input
rlabel metal3 s 31600 155120 32000 155176 6 itasegm[528]
port 515 nsew signal input
rlabel metal3 s 31600 155400 32000 155456 6 itasegm[529]
port 516 nsew signal input
rlabel metal3 s 0 46480 400 46536 6 itasegm[52]
port 517 nsew signal input
rlabel metal3 s 31600 155680 32000 155736 6 itasegm[530]
port 518 nsew signal input
rlabel metal3 s 31600 155960 32000 156016 6 itasegm[531]
port 519 nsew signal input
rlabel metal3 s 31600 156240 32000 156296 6 itasegm[532]
port 520 nsew signal input
rlabel metal3 s 31600 156520 32000 156576 6 itasegm[533]
port 521 nsew signal input
rlabel metal3 s 31600 156800 32000 156856 6 itasegm[534]
port 522 nsew signal input
rlabel metal3 s 31600 157080 32000 157136 6 itasegm[535]
port 523 nsew signal input
rlabel metal3 s 31600 157360 32000 157416 6 itasegm[536]
port 524 nsew signal input
rlabel metal3 s 31600 157640 32000 157696 6 itasegm[537]
port 525 nsew signal input
rlabel metal3 s 31600 157920 32000 157976 6 itasegm[538]
port 526 nsew signal input
rlabel metal3 s 31600 158200 32000 158256 6 itasegm[539]
port 527 nsew signal input
rlabel metal3 s 0 46760 400 46816 6 itasegm[53]
port 528 nsew signal input
rlabel metal3 s 31600 158480 32000 158536 6 itasegm[540]
port 529 nsew signal input
rlabel metal3 s 31600 158760 32000 158816 6 itasegm[541]
port 530 nsew signal input
rlabel metal3 s 31600 159040 32000 159096 6 itasegm[542]
port 531 nsew signal input
rlabel metal3 s 31600 159320 32000 159376 6 itasegm[543]
port 532 nsew signal input
rlabel metal3 s 31600 159600 32000 159656 6 itasegm[544]
port 533 nsew signal input
rlabel metal3 s 31600 159880 32000 159936 6 itasegm[545]
port 534 nsew signal input
rlabel metal3 s 31600 160160 32000 160216 6 itasegm[546]
port 535 nsew signal input
rlabel metal3 s 31600 160440 32000 160496 6 itasegm[547]
port 536 nsew signal input
rlabel metal3 s 31600 160720 32000 160776 6 itasegm[548]
port 537 nsew signal input
rlabel metal3 s 31600 161000 32000 161056 6 itasegm[549]
port 538 nsew signal input
rlabel metal3 s 0 47040 400 47096 6 itasegm[54]
port 539 nsew signal input
rlabel metal3 s 31600 161280 32000 161336 6 itasegm[550]
port 540 nsew signal input
rlabel metal3 s 31600 161560 32000 161616 6 itasegm[551]
port 541 nsew signal input
rlabel metal3 s 31600 161840 32000 161896 6 itasegm[552]
port 542 nsew signal input
rlabel metal3 s 31600 162120 32000 162176 6 itasegm[553]
port 543 nsew signal input
rlabel metal3 s 31600 162400 32000 162456 6 itasegm[554]
port 544 nsew signal input
rlabel metal3 s 31600 162680 32000 162736 6 itasegm[555]
port 545 nsew signal input
rlabel metal3 s 31600 162960 32000 163016 6 itasegm[556]
port 546 nsew signal input
rlabel metal3 s 31600 163240 32000 163296 6 itasegm[557]
port 547 nsew signal input
rlabel metal3 s 31600 163520 32000 163576 6 itasegm[558]
port 548 nsew signal input
rlabel metal3 s 31600 163800 32000 163856 6 itasegm[559]
port 549 nsew signal input
rlabel metal3 s 0 47320 400 47376 6 itasegm[55]
port 550 nsew signal input
rlabel metal3 s 0 177520 400 177576 6 itasegm[560]
port 551 nsew signal input
rlabel metal3 s 0 177800 400 177856 6 itasegm[561]
port 552 nsew signal input
rlabel metal3 s 0 178080 400 178136 6 itasegm[562]
port 553 nsew signal input
rlabel metal3 s 0 178360 400 178416 6 itasegm[563]
port 554 nsew signal input
rlabel metal3 s 0 178640 400 178696 6 itasegm[564]
port 555 nsew signal input
rlabel metal3 s 0 178920 400 178976 6 itasegm[565]
port 556 nsew signal input
rlabel metal3 s 0 179200 400 179256 6 itasegm[566]
port 557 nsew signal input
rlabel metal3 s 0 179480 400 179536 6 itasegm[567]
port 558 nsew signal input
rlabel metal3 s 0 179760 400 179816 6 itasegm[568]
port 559 nsew signal input
rlabel metal3 s 0 180040 400 180096 6 itasegm[569]
port 560 nsew signal input
rlabel metal3 s 31600 31920 32000 31976 6 itasegm[56]
port 561 nsew signal input
rlabel metal3 s 0 180320 400 180376 6 itasegm[570]
port 562 nsew signal input
rlabel metal3 s 0 180600 400 180656 6 itasegm[571]
port 563 nsew signal input
rlabel metal3 s 0 180880 400 180936 6 itasegm[572]
port 564 nsew signal input
rlabel metal3 s 0 181160 400 181216 6 itasegm[573]
port 565 nsew signal input
rlabel metal3 s 0 181440 400 181496 6 itasegm[574]
port 566 nsew signal input
rlabel metal3 s 0 181720 400 181776 6 itasegm[575]
port 567 nsew signal input
rlabel metal3 s 0 182000 400 182056 6 itasegm[576]
port 568 nsew signal input
rlabel metal3 s 0 182280 400 182336 6 itasegm[577]
port 569 nsew signal input
rlabel metal3 s 0 182560 400 182616 6 itasegm[578]
port 570 nsew signal input
rlabel metal3 s 0 182840 400 182896 6 itasegm[579]
port 571 nsew signal input
rlabel metal3 s 31600 32200 32000 32256 6 itasegm[57]
port 572 nsew signal input
rlabel metal3 s 0 183120 400 183176 6 itasegm[580]
port 573 nsew signal input
rlabel metal3 s 0 183400 400 183456 6 itasegm[581]
port 574 nsew signal input
rlabel metal3 s 0 183680 400 183736 6 itasegm[582]
port 575 nsew signal input
rlabel metal3 s 0 183960 400 184016 6 itasegm[583]
port 576 nsew signal input
rlabel metal3 s 0 184240 400 184296 6 itasegm[584]
port 577 nsew signal input
rlabel metal3 s 0 184520 400 184576 6 itasegm[585]
port 578 nsew signal input
rlabel metal3 s 0 184800 400 184856 6 itasegm[586]
port 579 nsew signal input
rlabel metal3 s 0 185080 400 185136 6 itasegm[587]
port 580 nsew signal input
rlabel metal3 s 0 185360 400 185416 6 itasegm[588]
port 581 nsew signal input
rlabel metal3 s 0 185640 400 185696 6 itasegm[589]
port 582 nsew signal input
rlabel metal3 s 31600 32480 32000 32536 6 itasegm[58]
port 583 nsew signal input
rlabel metal3 s 0 185920 400 185976 6 itasegm[590]
port 584 nsew signal input
rlabel metal3 s 0 186200 400 186256 6 itasegm[591]
port 585 nsew signal input
rlabel metal3 s 0 186480 400 186536 6 itasegm[592]
port 586 nsew signal input
rlabel metal3 s 0 186760 400 186816 6 itasegm[593]
port 587 nsew signal input
rlabel metal3 s 0 187040 400 187096 6 itasegm[594]
port 588 nsew signal input
rlabel metal3 s 0 187320 400 187376 6 itasegm[595]
port 589 nsew signal input
rlabel metal3 s 0 187600 400 187656 6 itasegm[596]
port 590 nsew signal input
rlabel metal3 s 0 187880 400 187936 6 itasegm[597]
port 591 nsew signal input
rlabel metal3 s 0 188160 400 188216 6 itasegm[598]
port 592 nsew signal input
rlabel metal3 s 0 188440 400 188496 6 itasegm[599]
port 593 nsew signal input
rlabel metal3 s 31600 32760 32000 32816 6 itasegm[59]
port 594 nsew signal input
rlabel metal3 s 0 33320 400 33376 6 itasegm[5]
port 595 nsew signal input
rlabel metal3 s 0 188720 400 188776 6 itasegm[600]
port 596 nsew signal input
rlabel metal3 s 0 189000 400 189056 6 itasegm[601]
port 597 nsew signal input
rlabel metal3 s 0 189280 400 189336 6 itasegm[602]
port 598 nsew signal input
rlabel metal3 s 0 189560 400 189616 6 itasegm[603]
port 599 nsew signal input
rlabel metal3 s 0 189840 400 189896 6 itasegm[604]
port 600 nsew signal input
rlabel metal3 s 0 190120 400 190176 6 itasegm[605]
port 601 nsew signal input
rlabel metal3 s 0 190400 400 190456 6 itasegm[606]
port 602 nsew signal input
rlabel metal3 s 0 190680 400 190736 6 itasegm[607]
port 603 nsew signal input
rlabel metal3 s 0 190960 400 191016 6 itasegm[608]
port 604 nsew signal input
rlabel metal3 s 0 191240 400 191296 6 itasegm[609]
port 605 nsew signal input
rlabel metal3 s 31600 33040 32000 33096 6 itasegm[60]
port 606 nsew signal input
rlabel metal3 s 0 191520 400 191576 6 itasegm[610]
port 607 nsew signal input
rlabel metal3 s 0 191800 400 191856 6 itasegm[611]
port 608 nsew signal input
rlabel metal3 s 0 192080 400 192136 6 itasegm[612]
port 609 nsew signal input
rlabel metal3 s 0 192360 400 192416 6 itasegm[613]
port 610 nsew signal input
rlabel metal3 s 0 192640 400 192696 6 itasegm[614]
port 611 nsew signal input
rlabel metal3 s 0 192920 400 192976 6 itasegm[615]
port 612 nsew signal input
rlabel metal3 s 31600 177520 32000 177576 6 itasegm[616]
port 613 nsew signal input
rlabel metal3 s 31600 177800 32000 177856 6 itasegm[617]
port 614 nsew signal input
rlabel metal3 s 31600 178080 32000 178136 6 itasegm[618]
port 615 nsew signal input
rlabel metal3 s 31600 178360 32000 178416 6 itasegm[619]
port 616 nsew signal input
rlabel metal3 s 31600 33320 32000 33376 6 itasegm[61]
port 617 nsew signal input
rlabel metal3 s 31600 178640 32000 178696 6 itasegm[620]
port 618 nsew signal input
rlabel metal3 s 31600 178920 32000 178976 6 itasegm[621]
port 619 nsew signal input
rlabel metal3 s 31600 179200 32000 179256 6 itasegm[622]
port 620 nsew signal input
rlabel metal3 s 31600 179480 32000 179536 6 itasegm[623]
port 621 nsew signal input
rlabel metal3 s 31600 179760 32000 179816 6 itasegm[624]
port 622 nsew signal input
rlabel metal3 s 31600 180040 32000 180096 6 itasegm[625]
port 623 nsew signal input
rlabel metal3 s 31600 180320 32000 180376 6 itasegm[626]
port 624 nsew signal input
rlabel metal3 s 31600 180600 32000 180656 6 itasegm[627]
port 625 nsew signal input
rlabel metal3 s 31600 180880 32000 180936 6 itasegm[628]
port 626 nsew signal input
rlabel metal3 s 31600 181160 32000 181216 6 itasegm[629]
port 627 nsew signal input
rlabel metal3 s 31600 33600 32000 33656 6 itasegm[62]
port 628 nsew signal input
rlabel metal3 s 31600 181440 32000 181496 6 itasegm[630]
port 629 nsew signal input
rlabel metal3 s 31600 181720 32000 181776 6 itasegm[631]
port 630 nsew signal input
rlabel metal3 s 31600 182000 32000 182056 6 itasegm[632]
port 631 nsew signal input
rlabel metal3 s 31600 182280 32000 182336 6 itasegm[633]
port 632 nsew signal input
rlabel metal3 s 31600 182560 32000 182616 6 itasegm[634]
port 633 nsew signal input
rlabel metal3 s 31600 182840 32000 182896 6 itasegm[635]
port 634 nsew signal input
rlabel metal3 s 31600 183120 32000 183176 6 itasegm[636]
port 635 nsew signal input
rlabel metal3 s 31600 183400 32000 183456 6 itasegm[637]
port 636 nsew signal input
rlabel metal3 s 31600 183680 32000 183736 6 itasegm[638]
port 637 nsew signal input
rlabel metal3 s 31600 183960 32000 184016 6 itasegm[639]
port 638 nsew signal input
rlabel metal3 s 31600 33880 32000 33936 6 itasegm[63]
port 639 nsew signal input
rlabel metal3 s 31600 184240 32000 184296 6 itasegm[640]
port 640 nsew signal input
rlabel metal3 s 31600 184520 32000 184576 6 itasegm[641]
port 641 nsew signal input
rlabel metal3 s 31600 184800 32000 184856 6 itasegm[642]
port 642 nsew signal input
rlabel metal3 s 31600 185080 32000 185136 6 itasegm[643]
port 643 nsew signal input
rlabel metal3 s 31600 185360 32000 185416 6 itasegm[644]
port 644 nsew signal input
rlabel metal3 s 31600 185640 32000 185696 6 itasegm[645]
port 645 nsew signal input
rlabel metal3 s 31600 185920 32000 185976 6 itasegm[646]
port 646 nsew signal input
rlabel metal3 s 31600 186200 32000 186256 6 itasegm[647]
port 647 nsew signal input
rlabel metal3 s 31600 186480 32000 186536 6 itasegm[648]
port 648 nsew signal input
rlabel metal3 s 31600 186760 32000 186816 6 itasegm[649]
port 649 nsew signal input
rlabel metal3 s 31600 34160 32000 34216 6 itasegm[64]
port 650 nsew signal input
rlabel metal3 s 31600 187040 32000 187096 6 itasegm[650]
port 651 nsew signal input
rlabel metal3 s 31600 187320 32000 187376 6 itasegm[651]
port 652 nsew signal input
rlabel metal3 s 31600 187600 32000 187656 6 itasegm[652]
port 653 nsew signal input
rlabel metal3 s 31600 187880 32000 187936 6 itasegm[653]
port 654 nsew signal input
rlabel metal3 s 31600 188160 32000 188216 6 itasegm[654]
port 655 nsew signal input
rlabel metal3 s 31600 188440 32000 188496 6 itasegm[655]
port 656 nsew signal input
rlabel metal3 s 31600 188720 32000 188776 6 itasegm[656]
port 657 nsew signal input
rlabel metal3 s 31600 189000 32000 189056 6 itasegm[657]
port 658 nsew signal input
rlabel metal3 s 31600 189280 32000 189336 6 itasegm[658]
port 659 nsew signal input
rlabel metal3 s 31600 189560 32000 189616 6 itasegm[659]
port 660 nsew signal input
rlabel metal3 s 31600 34440 32000 34496 6 itasegm[65]
port 661 nsew signal input
rlabel metal3 s 31600 189840 32000 189896 6 itasegm[660]
port 662 nsew signal input
rlabel metal3 s 31600 190120 32000 190176 6 itasegm[661]
port 663 nsew signal input
rlabel metal3 s 31600 190400 32000 190456 6 itasegm[662]
port 664 nsew signal input
rlabel metal3 s 31600 190680 32000 190736 6 itasegm[663]
port 665 nsew signal input
rlabel metal3 s 31600 190960 32000 191016 6 itasegm[664]
port 666 nsew signal input
rlabel metal3 s 31600 191240 32000 191296 6 itasegm[665]
port 667 nsew signal input
rlabel metal3 s 31600 191520 32000 191576 6 itasegm[666]
port 668 nsew signal input
rlabel metal3 s 31600 191800 32000 191856 6 itasegm[667]
port 669 nsew signal input
rlabel metal3 s 31600 192080 32000 192136 6 itasegm[668]
port 670 nsew signal input
rlabel metal3 s 31600 192360 32000 192416 6 itasegm[669]
port 671 nsew signal input
rlabel metal3 s 31600 34720 32000 34776 6 itasegm[66]
port 672 nsew signal input
rlabel metal3 s 31600 192640 32000 192696 6 itasegm[670]
port 673 nsew signal input
rlabel metal3 s 31600 192920 32000 192976 6 itasegm[671]
port 674 nsew signal input
rlabel metal3 s 0 206640 400 206696 6 itasegm[672]
port 675 nsew signal input
rlabel metal3 s 0 206920 400 206976 6 itasegm[673]
port 676 nsew signal input
rlabel metal3 s 0 207200 400 207256 6 itasegm[674]
port 677 nsew signal input
rlabel metal3 s 0 207480 400 207536 6 itasegm[675]
port 678 nsew signal input
rlabel metal3 s 0 207760 400 207816 6 itasegm[676]
port 679 nsew signal input
rlabel metal3 s 0 208040 400 208096 6 itasegm[677]
port 680 nsew signal input
rlabel metal3 s 0 208320 400 208376 6 itasegm[678]
port 681 nsew signal input
rlabel metal3 s 0 208600 400 208656 6 itasegm[679]
port 682 nsew signal input
rlabel metal3 s 31600 35000 32000 35056 6 itasegm[67]
port 683 nsew signal input
rlabel metal3 s 0 208880 400 208936 6 itasegm[680]
port 684 nsew signal input
rlabel metal3 s 0 209160 400 209216 6 itasegm[681]
port 685 nsew signal input
rlabel metal3 s 0 209440 400 209496 6 itasegm[682]
port 686 nsew signal input
rlabel metal3 s 0 209720 400 209776 6 itasegm[683]
port 687 nsew signal input
rlabel metal3 s 0 210000 400 210056 6 itasegm[684]
port 688 nsew signal input
rlabel metal3 s 0 210280 400 210336 6 itasegm[685]
port 689 nsew signal input
rlabel metal3 s 0 210560 400 210616 6 itasegm[686]
port 690 nsew signal input
rlabel metal3 s 0 210840 400 210896 6 itasegm[687]
port 691 nsew signal input
rlabel metal3 s 0 211120 400 211176 6 itasegm[688]
port 692 nsew signal input
rlabel metal3 s 0 211400 400 211456 6 itasegm[689]
port 693 nsew signal input
rlabel metal3 s 31600 35280 32000 35336 6 itasegm[68]
port 694 nsew signal input
rlabel metal3 s 0 211680 400 211736 6 itasegm[690]
port 695 nsew signal input
rlabel metal3 s 0 211960 400 212016 6 itasegm[691]
port 696 nsew signal input
rlabel metal3 s 0 212240 400 212296 6 itasegm[692]
port 697 nsew signal input
rlabel metal3 s 0 212520 400 212576 6 itasegm[693]
port 698 nsew signal input
rlabel metal3 s 0 212800 400 212856 6 itasegm[694]
port 699 nsew signal input
rlabel metal3 s 0 213080 400 213136 6 itasegm[695]
port 700 nsew signal input
rlabel metal3 s 0 213360 400 213416 6 itasegm[696]
port 701 nsew signal input
rlabel metal3 s 0 213640 400 213696 6 itasegm[697]
port 702 nsew signal input
rlabel metal3 s 0 213920 400 213976 6 itasegm[698]
port 703 nsew signal input
rlabel metal3 s 0 214200 400 214256 6 itasegm[699]
port 704 nsew signal input
rlabel metal3 s 31600 35560 32000 35616 6 itasegm[69]
port 705 nsew signal input
rlabel metal3 s 0 33600 400 33656 6 itasegm[6]
port 706 nsew signal input
rlabel metal3 s 0 214480 400 214536 6 itasegm[700]
port 707 nsew signal input
rlabel metal3 s 0 214760 400 214816 6 itasegm[701]
port 708 nsew signal input
rlabel metal3 s 0 215040 400 215096 6 itasegm[702]
port 709 nsew signal input
rlabel metal3 s 0 215320 400 215376 6 itasegm[703]
port 710 nsew signal input
rlabel metal3 s 0 215600 400 215656 6 itasegm[704]
port 711 nsew signal input
rlabel metal3 s 0 215880 400 215936 6 itasegm[705]
port 712 nsew signal input
rlabel metal3 s 0 216160 400 216216 6 itasegm[706]
port 713 nsew signal input
rlabel metal3 s 0 216440 400 216496 6 itasegm[707]
port 714 nsew signal input
rlabel metal3 s 0 216720 400 216776 6 itasegm[708]
port 715 nsew signal input
rlabel metal3 s 0 217000 400 217056 6 itasegm[709]
port 716 nsew signal input
rlabel metal3 s 31600 35840 32000 35896 6 itasegm[70]
port 717 nsew signal input
rlabel metal3 s 0 217280 400 217336 6 itasegm[710]
port 718 nsew signal input
rlabel metal3 s 0 217560 400 217616 6 itasegm[711]
port 719 nsew signal input
rlabel metal3 s 0 217840 400 217896 6 itasegm[712]
port 720 nsew signal input
rlabel metal3 s 0 218120 400 218176 6 itasegm[713]
port 721 nsew signal input
rlabel metal3 s 0 218400 400 218456 6 itasegm[714]
port 722 nsew signal input
rlabel metal3 s 0 218680 400 218736 6 itasegm[715]
port 723 nsew signal input
rlabel metal3 s 0 218960 400 219016 6 itasegm[716]
port 724 nsew signal input
rlabel metal3 s 0 219240 400 219296 6 itasegm[717]
port 725 nsew signal input
rlabel metal3 s 0 219520 400 219576 6 itasegm[718]
port 726 nsew signal input
rlabel metal3 s 0 219800 400 219856 6 itasegm[719]
port 727 nsew signal input
rlabel metal3 s 31600 36120 32000 36176 6 itasegm[71]
port 728 nsew signal input
rlabel metal3 s 0 220080 400 220136 6 itasegm[720]
port 729 nsew signal input
rlabel metal3 s 0 220360 400 220416 6 itasegm[721]
port 730 nsew signal input
rlabel metal3 s 0 220640 400 220696 6 itasegm[722]
port 731 nsew signal input
rlabel metal3 s 0 220920 400 220976 6 itasegm[723]
port 732 nsew signal input
rlabel metal3 s 0 221200 400 221256 6 itasegm[724]
port 733 nsew signal input
rlabel metal3 s 0 221480 400 221536 6 itasegm[725]
port 734 nsew signal input
rlabel metal3 s 0 221760 400 221816 6 itasegm[726]
port 735 nsew signal input
rlabel metal3 s 0 222040 400 222096 6 itasegm[727]
port 736 nsew signal input
rlabel metal3 s 31600 206640 32000 206696 6 itasegm[728]
port 737 nsew signal input
rlabel metal3 s 31600 206920 32000 206976 6 itasegm[729]
port 738 nsew signal input
rlabel metal3 s 31600 36400 32000 36456 6 itasegm[72]
port 739 nsew signal input
rlabel metal3 s 31600 207200 32000 207256 6 itasegm[730]
port 740 nsew signal input
rlabel metal3 s 31600 207480 32000 207536 6 itasegm[731]
port 741 nsew signal input
rlabel metal3 s 31600 207760 32000 207816 6 itasegm[732]
port 742 nsew signal input
rlabel metal3 s 31600 208040 32000 208096 6 itasegm[733]
port 743 nsew signal input
rlabel metal3 s 31600 208320 32000 208376 6 itasegm[734]
port 744 nsew signal input
rlabel metal3 s 31600 208600 32000 208656 6 itasegm[735]
port 745 nsew signal input
rlabel metal3 s 31600 208880 32000 208936 6 itasegm[736]
port 746 nsew signal input
rlabel metal3 s 31600 209160 32000 209216 6 itasegm[737]
port 747 nsew signal input
rlabel metal3 s 31600 209440 32000 209496 6 itasegm[738]
port 748 nsew signal input
rlabel metal3 s 31600 209720 32000 209776 6 itasegm[739]
port 749 nsew signal input
rlabel metal3 s 31600 36680 32000 36736 6 itasegm[73]
port 750 nsew signal input
rlabel metal3 s 31600 210000 32000 210056 6 itasegm[740]
port 751 nsew signal input
rlabel metal3 s 31600 210280 32000 210336 6 itasegm[741]
port 752 nsew signal input
rlabel metal3 s 31600 210560 32000 210616 6 itasegm[742]
port 753 nsew signal input
rlabel metal3 s 31600 210840 32000 210896 6 itasegm[743]
port 754 nsew signal input
rlabel metal3 s 31600 211120 32000 211176 6 itasegm[744]
port 755 nsew signal input
rlabel metal3 s 31600 211400 32000 211456 6 itasegm[745]
port 756 nsew signal input
rlabel metal3 s 31600 211680 32000 211736 6 itasegm[746]
port 757 nsew signal input
rlabel metal3 s 31600 211960 32000 212016 6 itasegm[747]
port 758 nsew signal input
rlabel metal3 s 31600 212240 32000 212296 6 itasegm[748]
port 759 nsew signal input
rlabel metal3 s 31600 212520 32000 212576 6 itasegm[749]
port 760 nsew signal input
rlabel metal3 s 31600 36960 32000 37016 6 itasegm[74]
port 761 nsew signal input
rlabel metal3 s 31600 212800 32000 212856 6 itasegm[750]
port 762 nsew signal input
rlabel metal3 s 31600 213080 32000 213136 6 itasegm[751]
port 763 nsew signal input
rlabel metal3 s 31600 213360 32000 213416 6 itasegm[752]
port 764 nsew signal input
rlabel metal3 s 31600 213640 32000 213696 6 itasegm[753]
port 765 nsew signal input
rlabel metal3 s 31600 213920 32000 213976 6 itasegm[754]
port 766 nsew signal input
rlabel metal3 s 31600 214200 32000 214256 6 itasegm[755]
port 767 nsew signal input
rlabel metal3 s 31600 214480 32000 214536 6 itasegm[756]
port 768 nsew signal input
rlabel metal3 s 31600 214760 32000 214816 6 itasegm[757]
port 769 nsew signal input
rlabel metal3 s 31600 215040 32000 215096 6 itasegm[758]
port 770 nsew signal input
rlabel metal3 s 31600 215320 32000 215376 6 itasegm[759]
port 771 nsew signal input
rlabel metal3 s 31600 37240 32000 37296 6 itasegm[75]
port 772 nsew signal input
rlabel metal3 s 31600 215600 32000 215656 6 itasegm[760]
port 773 nsew signal input
rlabel metal3 s 31600 215880 32000 215936 6 itasegm[761]
port 774 nsew signal input
rlabel metal3 s 31600 216160 32000 216216 6 itasegm[762]
port 775 nsew signal input
rlabel metal3 s 31600 216440 32000 216496 6 itasegm[763]
port 776 nsew signal input
rlabel metal3 s 31600 216720 32000 216776 6 itasegm[764]
port 777 nsew signal input
rlabel metal3 s 31600 217000 32000 217056 6 itasegm[765]
port 778 nsew signal input
rlabel metal3 s 31600 217280 32000 217336 6 itasegm[766]
port 779 nsew signal input
rlabel metal3 s 31600 217560 32000 217616 6 itasegm[767]
port 780 nsew signal input
rlabel metal3 s 31600 217840 32000 217896 6 itasegm[768]
port 781 nsew signal input
rlabel metal3 s 31600 218120 32000 218176 6 itasegm[769]
port 782 nsew signal input
rlabel metal3 s 31600 37520 32000 37576 6 itasegm[76]
port 783 nsew signal input
rlabel metal3 s 31600 218400 32000 218456 6 itasegm[770]
port 784 nsew signal input
rlabel metal3 s 31600 218680 32000 218736 6 itasegm[771]
port 785 nsew signal input
rlabel metal3 s 31600 218960 32000 219016 6 itasegm[772]
port 786 nsew signal input
rlabel metal3 s 31600 219240 32000 219296 6 itasegm[773]
port 787 nsew signal input
rlabel metal3 s 31600 219520 32000 219576 6 itasegm[774]
port 788 nsew signal input
rlabel metal3 s 31600 219800 32000 219856 6 itasegm[775]
port 789 nsew signal input
rlabel metal3 s 31600 220080 32000 220136 6 itasegm[776]
port 790 nsew signal input
rlabel metal3 s 31600 220360 32000 220416 6 itasegm[777]
port 791 nsew signal input
rlabel metal3 s 31600 220640 32000 220696 6 itasegm[778]
port 792 nsew signal input
rlabel metal3 s 31600 220920 32000 220976 6 itasegm[779]
port 793 nsew signal input
rlabel metal3 s 31600 37800 32000 37856 6 itasegm[77]
port 794 nsew signal input
rlabel metal3 s 31600 221200 32000 221256 6 itasegm[780]
port 795 nsew signal input
rlabel metal3 s 31600 221480 32000 221536 6 itasegm[781]
port 796 nsew signal input
rlabel metal3 s 31600 221760 32000 221816 6 itasegm[782]
port 797 nsew signal input
rlabel metal3 s 31600 222040 32000 222096 6 itasegm[783]
port 798 nsew signal input
rlabel metal3 s 0 235760 400 235816 6 itasegm[784]
port 799 nsew signal input
rlabel metal3 s 0 236040 400 236096 6 itasegm[785]
port 800 nsew signal input
rlabel metal3 s 0 236320 400 236376 6 itasegm[786]
port 801 nsew signal input
rlabel metal3 s 0 236600 400 236656 6 itasegm[787]
port 802 nsew signal input
rlabel metal3 s 0 236880 400 236936 6 itasegm[788]
port 803 nsew signal input
rlabel metal3 s 0 237160 400 237216 6 itasegm[789]
port 804 nsew signal input
rlabel metal3 s 31600 38080 32000 38136 6 itasegm[78]
port 805 nsew signal input
rlabel metal3 s 0 237440 400 237496 6 itasegm[790]
port 806 nsew signal input
rlabel metal3 s 0 237720 400 237776 6 itasegm[791]
port 807 nsew signal input
rlabel metal3 s 0 238000 400 238056 6 itasegm[792]
port 808 nsew signal input
rlabel metal3 s 0 238280 400 238336 6 itasegm[793]
port 809 nsew signal input
rlabel metal3 s 0 238560 400 238616 6 itasegm[794]
port 810 nsew signal input
rlabel metal3 s 0 238840 400 238896 6 itasegm[795]
port 811 nsew signal input
rlabel metal3 s 0 239120 400 239176 6 itasegm[796]
port 812 nsew signal input
rlabel metal3 s 0 239400 400 239456 6 itasegm[797]
port 813 nsew signal input
rlabel metal3 s 0 239680 400 239736 6 itasegm[798]
port 814 nsew signal input
rlabel metal3 s 0 239960 400 240016 6 itasegm[799]
port 815 nsew signal input
rlabel metal3 s 31600 38360 32000 38416 6 itasegm[79]
port 816 nsew signal input
rlabel metal3 s 0 33880 400 33936 6 itasegm[7]
port 817 nsew signal input
rlabel metal3 s 0 240240 400 240296 6 itasegm[800]
port 818 nsew signal input
rlabel metal3 s 0 240520 400 240576 6 itasegm[801]
port 819 nsew signal input
rlabel metal3 s 0 240800 400 240856 6 itasegm[802]
port 820 nsew signal input
rlabel metal3 s 0 241080 400 241136 6 itasegm[803]
port 821 nsew signal input
rlabel metal3 s 0 241360 400 241416 6 itasegm[804]
port 822 nsew signal input
rlabel metal3 s 0 241640 400 241696 6 itasegm[805]
port 823 nsew signal input
rlabel metal3 s 0 241920 400 241976 6 itasegm[806]
port 824 nsew signal input
rlabel metal3 s 0 242200 400 242256 6 itasegm[807]
port 825 nsew signal input
rlabel metal3 s 0 242480 400 242536 6 itasegm[808]
port 826 nsew signal input
rlabel metal3 s 0 242760 400 242816 6 itasegm[809]
port 827 nsew signal input
rlabel metal3 s 31600 38640 32000 38696 6 itasegm[80]
port 828 nsew signal input
rlabel metal3 s 0 243040 400 243096 6 itasegm[810]
port 829 nsew signal input
rlabel metal3 s 0 243320 400 243376 6 itasegm[811]
port 830 nsew signal input
rlabel metal3 s 0 243600 400 243656 6 itasegm[812]
port 831 nsew signal input
rlabel metal3 s 0 243880 400 243936 6 itasegm[813]
port 832 nsew signal input
rlabel metal3 s 0 244160 400 244216 6 itasegm[814]
port 833 nsew signal input
rlabel metal3 s 0 244440 400 244496 6 itasegm[815]
port 834 nsew signal input
rlabel metal3 s 0 244720 400 244776 6 itasegm[816]
port 835 nsew signal input
rlabel metal3 s 0 245000 400 245056 6 itasegm[817]
port 836 nsew signal input
rlabel metal3 s 0 245280 400 245336 6 itasegm[818]
port 837 nsew signal input
rlabel metal3 s 0 245560 400 245616 6 itasegm[819]
port 838 nsew signal input
rlabel metal3 s 31600 38920 32000 38976 6 itasegm[81]
port 839 nsew signal input
rlabel metal3 s 0 245840 400 245896 6 itasegm[820]
port 840 nsew signal input
rlabel metal3 s 0 246120 400 246176 6 itasegm[821]
port 841 nsew signal input
rlabel metal3 s 0 246400 400 246456 6 itasegm[822]
port 842 nsew signal input
rlabel metal3 s 0 246680 400 246736 6 itasegm[823]
port 843 nsew signal input
rlabel metal3 s 0 246960 400 247016 6 itasegm[824]
port 844 nsew signal input
rlabel metal3 s 0 247240 400 247296 6 itasegm[825]
port 845 nsew signal input
rlabel metal3 s 0 247520 400 247576 6 itasegm[826]
port 846 nsew signal input
rlabel metal3 s 0 247800 400 247856 6 itasegm[827]
port 847 nsew signal input
rlabel metal3 s 0 248080 400 248136 6 itasegm[828]
port 848 nsew signal input
rlabel metal3 s 0 248360 400 248416 6 itasegm[829]
port 849 nsew signal input
rlabel metal3 s 31600 39200 32000 39256 6 itasegm[82]
port 850 nsew signal input
rlabel metal3 s 0 248640 400 248696 6 itasegm[830]
port 851 nsew signal input
rlabel metal3 s 0 248920 400 248976 6 itasegm[831]
port 852 nsew signal input
rlabel metal3 s 0 249200 400 249256 6 itasegm[832]
port 853 nsew signal input
rlabel metal3 s 0 249480 400 249536 6 itasegm[833]
port 854 nsew signal input
rlabel metal3 s 0 249760 400 249816 6 itasegm[834]
port 855 nsew signal input
rlabel metal3 s 0 250040 400 250096 6 itasegm[835]
port 856 nsew signal input
rlabel metal3 s 0 250320 400 250376 6 itasegm[836]
port 857 nsew signal input
rlabel metal3 s 0 250600 400 250656 6 itasegm[837]
port 858 nsew signal input
rlabel metal3 s 0 250880 400 250936 6 itasegm[838]
port 859 nsew signal input
rlabel metal3 s 0 251160 400 251216 6 itasegm[839]
port 860 nsew signal input
rlabel metal3 s 31600 39480 32000 39536 6 itasegm[83]
port 861 nsew signal input
rlabel metal3 s 31600 235760 32000 235816 6 itasegm[840]
port 862 nsew signal input
rlabel metal3 s 31600 236040 32000 236096 6 itasegm[841]
port 863 nsew signal input
rlabel metal3 s 31600 236320 32000 236376 6 itasegm[842]
port 864 nsew signal input
rlabel metal3 s 31600 236600 32000 236656 6 itasegm[843]
port 865 nsew signal input
rlabel metal3 s 31600 236880 32000 236936 6 itasegm[844]
port 866 nsew signal input
rlabel metal3 s 31600 237160 32000 237216 6 itasegm[845]
port 867 nsew signal input
rlabel metal3 s 31600 237440 32000 237496 6 itasegm[846]
port 868 nsew signal input
rlabel metal3 s 31600 237720 32000 237776 6 itasegm[847]
port 869 nsew signal input
rlabel metal3 s 31600 238000 32000 238056 6 itasegm[848]
port 870 nsew signal input
rlabel metal3 s 31600 238280 32000 238336 6 itasegm[849]
port 871 nsew signal input
rlabel metal3 s 31600 39760 32000 39816 6 itasegm[84]
port 872 nsew signal input
rlabel metal3 s 31600 238560 32000 238616 6 itasegm[850]
port 873 nsew signal input
rlabel metal3 s 31600 238840 32000 238896 6 itasegm[851]
port 874 nsew signal input
rlabel metal3 s 31600 239120 32000 239176 6 itasegm[852]
port 875 nsew signal input
rlabel metal3 s 31600 239400 32000 239456 6 itasegm[853]
port 876 nsew signal input
rlabel metal3 s 31600 239680 32000 239736 6 itasegm[854]
port 877 nsew signal input
rlabel metal3 s 31600 239960 32000 240016 6 itasegm[855]
port 878 nsew signal input
rlabel metal3 s 31600 240240 32000 240296 6 itasegm[856]
port 879 nsew signal input
rlabel metal3 s 31600 240520 32000 240576 6 itasegm[857]
port 880 nsew signal input
rlabel metal3 s 31600 240800 32000 240856 6 itasegm[858]
port 881 nsew signal input
rlabel metal3 s 31600 241080 32000 241136 6 itasegm[859]
port 882 nsew signal input
rlabel metal3 s 31600 40040 32000 40096 6 itasegm[85]
port 883 nsew signal input
rlabel metal3 s 31600 241360 32000 241416 6 itasegm[860]
port 884 nsew signal input
rlabel metal3 s 31600 241640 32000 241696 6 itasegm[861]
port 885 nsew signal input
rlabel metal3 s 31600 241920 32000 241976 6 itasegm[862]
port 886 nsew signal input
rlabel metal3 s 31600 242200 32000 242256 6 itasegm[863]
port 887 nsew signal input
rlabel metal3 s 31600 242480 32000 242536 6 itasegm[864]
port 888 nsew signal input
rlabel metal3 s 31600 242760 32000 242816 6 itasegm[865]
port 889 nsew signal input
rlabel metal3 s 31600 243040 32000 243096 6 itasegm[866]
port 890 nsew signal input
rlabel metal3 s 31600 243320 32000 243376 6 itasegm[867]
port 891 nsew signal input
rlabel metal3 s 31600 243600 32000 243656 6 itasegm[868]
port 892 nsew signal input
rlabel metal3 s 31600 243880 32000 243936 6 itasegm[869]
port 893 nsew signal input
rlabel metal3 s 31600 40320 32000 40376 6 itasegm[86]
port 894 nsew signal input
rlabel metal3 s 31600 244160 32000 244216 6 itasegm[870]
port 895 nsew signal input
rlabel metal3 s 31600 244440 32000 244496 6 itasegm[871]
port 896 nsew signal input
rlabel metal3 s 31600 244720 32000 244776 6 itasegm[872]
port 897 nsew signal input
rlabel metal3 s 31600 245000 32000 245056 6 itasegm[873]
port 898 nsew signal input
rlabel metal3 s 31600 245280 32000 245336 6 itasegm[874]
port 899 nsew signal input
rlabel metal3 s 31600 245560 32000 245616 6 itasegm[875]
port 900 nsew signal input
rlabel metal3 s 31600 245840 32000 245896 6 itasegm[876]
port 901 nsew signal input
rlabel metal3 s 31600 246120 32000 246176 6 itasegm[877]
port 902 nsew signal input
rlabel metal3 s 31600 246400 32000 246456 6 itasegm[878]
port 903 nsew signal input
rlabel metal3 s 31600 246680 32000 246736 6 itasegm[879]
port 904 nsew signal input
rlabel metal3 s 31600 40600 32000 40656 6 itasegm[87]
port 905 nsew signal input
rlabel metal3 s 31600 246960 32000 247016 6 itasegm[880]
port 906 nsew signal input
rlabel metal3 s 31600 247240 32000 247296 6 itasegm[881]
port 907 nsew signal input
rlabel metal3 s 31600 247520 32000 247576 6 itasegm[882]
port 908 nsew signal input
rlabel metal3 s 31600 247800 32000 247856 6 itasegm[883]
port 909 nsew signal input
rlabel metal3 s 31600 248080 32000 248136 6 itasegm[884]
port 910 nsew signal input
rlabel metal3 s 31600 248360 32000 248416 6 itasegm[885]
port 911 nsew signal input
rlabel metal3 s 31600 248640 32000 248696 6 itasegm[886]
port 912 nsew signal input
rlabel metal3 s 31600 248920 32000 248976 6 itasegm[887]
port 913 nsew signal input
rlabel metal3 s 31600 249200 32000 249256 6 itasegm[888]
port 914 nsew signal input
rlabel metal3 s 31600 249480 32000 249536 6 itasegm[889]
port 915 nsew signal input
rlabel metal3 s 31600 40880 32000 40936 6 itasegm[88]
port 916 nsew signal input
rlabel metal3 s 31600 249760 32000 249816 6 itasegm[890]
port 917 nsew signal input
rlabel metal3 s 31600 250040 32000 250096 6 itasegm[891]
port 918 nsew signal input
rlabel metal3 s 31600 250320 32000 250376 6 itasegm[892]
port 919 nsew signal input
rlabel metal3 s 31600 250600 32000 250656 6 itasegm[893]
port 920 nsew signal input
rlabel metal3 s 31600 250880 32000 250936 6 itasegm[894]
port 921 nsew signal input
rlabel metal3 s 31600 251160 32000 251216 6 itasegm[895]
port 922 nsew signal input
rlabel metal3 s 31600 41160 32000 41216 6 itasegm[89]
port 923 nsew signal input
rlabel metal3 s 0 34160 400 34216 6 itasegm[8]
port 924 nsew signal input
rlabel metal3 s 31600 41440 32000 41496 6 itasegm[90]
port 925 nsew signal input
rlabel metal3 s 31600 41720 32000 41776 6 itasegm[91]
port 926 nsew signal input
rlabel metal3 s 31600 42000 32000 42056 6 itasegm[92]
port 927 nsew signal input
rlabel metal3 s 31600 42280 32000 42336 6 itasegm[93]
port 928 nsew signal input
rlabel metal3 s 31600 42560 32000 42616 6 itasegm[94]
port 929 nsew signal input
rlabel metal3 s 31600 42840 32000 42896 6 itasegm[95]
port 930 nsew signal input
rlabel metal3 s 31600 43120 32000 43176 6 itasegm[96]
port 931 nsew signal input
rlabel metal3 s 31600 43400 32000 43456 6 itasegm[97]
port 932 nsew signal input
rlabel metal3 s 31600 43680 32000 43736 6 itasegm[98]
port 933 nsew signal input
rlabel metal3 s 31600 43960 32000 44016 6 itasegm[99]
port 934 nsew signal input
rlabel metal3 s 0 34440 400 34496 6 itasegm[9]
port 935 nsew signal input
rlabel metal3 s 0 18480 400 18536 6 itasel[0]
port 936 nsew signal input
rlabel metal3 s 0 48720 400 48776 6 itasel[100]
port 937 nsew signal input
rlabel metal3 s 0 49000 400 49056 6 itasel[101]
port 938 nsew signal input
rlabel metal3 s 0 49280 400 49336 6 itasel[102]
port 939 nsew signal input
rlabel metal3 s 0 49560 400 49616 6 itasel[103]
port 940 nsew signal input
rlabel metal3 s 0 49840 400 49896 6 itasel[104]
port 941 nsew signal input
rlabel metal3 s 0 50120 400 50176 6 itasel[105]
port 942 nsew signal input
rlabel metal3 s 0 50400 400 50456 6 itasel[106]
port 943 nsew signal input
rlabel metal3 s 0 50680 400 50736 6 itasel[107]
port 944 nsew signal input
rlabel metal3 s 0 50960 400 51016 6 itasel[108]
port 945 nsew signal input
rlabel metal3 s 0 51240 400 51296 6 itasel[109]
port 946 nsew signal input
rlabel metal3 s 0 21280 400 21336 6 itasel[10]
port 947 nsew signal input
rlabel metal3 s 0 51520 400 51576 6 itasel[110]
port 948 nsew signal input
rlabel metal3 s 0 51800 400 51856 6 itasel[111]
port 949 nsew signal input
rlabel metal3 s 0 52080 400 52136 6 itasel[112]
port 950 nsew signal input
rlabel metal3 s 0 52360 400 52416 6 itasel[113]
port 951 nsew signal input
rlabel metal3 s 0 52640 400 52696 6 itasel[114]
port 952 nsew signal input
rlabel metal3 s 0 52920 400 52976 6 itasel[115]
port 953 nsew signal input
rlabel metal3 s 0 53200 400 53256 6 itasel[116]
port 954 nsew signal input
rlabel metal3 s 0 53480 400 53536 6 itasel[117]
port 955 nsew signal input
rlabel metal3 s 0 53760 400 53816 6 itasel[118]
port 956 nsew signal input
rlabel metal3 s 0 54040 400 54096 6 itasel[119]
port 957 nsew signal input
rlabel metal3 s 0 21560 400 21616 6 itasel[11]
port 958 nsew signal input
rlabel metal3 s 0 54320 400 54376 6 itasel[120]
port 959 nsew signal input
rlabel metal3 s 0 54600 400 54656 6 itasel[121]
port 960 nsew signal input
rlabel metal3 s 0 54880 400 54936 6 itasel[122]
port 961 nsew signal input
rlabel metal3 s 0 55160 400 55216 6 itasel[123]
port 962 nsew signal input
rlabel metal3 s 0 55440 400 55496 6 itasel[124]
port 963 nsew signal input
rlabel metal3 s 0 55720 400 55776 6 itasel[125]
port 964 nsew signal input
rlabel metal3 s 0 56000 400 56056 6 itasel[126]
port 965 nsew signal input
rlabel metal3 s 0 56280 400 56336 6 itasel[127]
port 966 nsew signal input
rlabel metal3 s 0 56560 400 56616 6 itasel[128]
port 967 nsew signal input
rlabel metal3 s 0 56840 400 56896 6 itasel[129]
port 968 nsew signal input
rlabel metal3 s 0 21840 400 21896 6 itasel[12]
port 969 nsew signal input
rlabel metal3 s 0 57120 400 57176 6 itasel[130]
port 970 nsew signal input
rlabel metal3 s 0 57400 400 57456 6 itasel[131]
port 971 nsew signal input
rlabel metal3 s 0 57680 400 57736 6 itasel[132]
port 972 nsew signal input
rlabel metal3 s 0 57960 400 58016 6 itasel[133]
port 973 nsew signal input
rlabel metal3 s 0 58240 400 58296 6 itasel[134]
port 974 nsew signal input
rlabel metal3 s 0 58520 400 58576 6 itasel[135]
port 975 nsew signal input
rlabel metal3 s 0 58800 400 58856 6 itasel[136]
port 976 nsew signal input
rlabel metal3 s 0 59080 400 59136 6 itasel[137]
port 977 nsew signal input
rlabel metal3 s 0 59360 400 59416 6 itasel[138]
port 978 nsew signal input
rlabel metal3 s 0 59640 400 59696 6 itasel[139]
port 979 nsew signal input
rlabel metal3 s 0 22120 400 22176 6 itasel[13]
port 980 nsew signal input
rlabel metal3 s 0 59920 400 59976 6 itasel[140]
port 981 nsew signal input
rlabel metal3 s 0 60200 400 60256 6 itasel[141]
port 982 nsew signal input
rlabel metal3 s 0 60480 400 60536 6 itasel[142]
port 983 nsew signal input
rlabel metal3 s 0 60760 400 60816 6 itasel[143]
port 984 nsew signal input
rlabel metal3 s 31600 47600 32000 47656 6 itasel[144]
port 985 nsew signal input
rlabel metal3 s 31600 47880 32000 47936 6 itasel[145]
port 986 nsew signal input
rlabel metal3 s 31600 48160 32000 48216 6 itasel[146]
port 987 nsew signal input
rlabel metal3 s 31600 48440 32000 48496 6 itasel[147]
port 988 nsew signal input
rlabel metal3 s 31600 48720 32000 48776 6 itasel[148]
port 989 nsew signal input
rlabel metal3 s 31600 49000 32000 49056 6 itasel[149]
port 990 nsew signal input
rlabel metal3 s 0 22400 400 22456 6 itasel[14]
port 991 nsew signal input
rlabel metal3 s 31600 49280 32000 49336 6 itasel[150]
port 992 nsew signal input
rlabel metal3 s 31600 49560 32000 49616 6 itasel[151]
port 993 nsew signal input
rlabel metal3 s 31600 49840 32000 49896 6 itasel[152]
port 994 nsew signal input
rlabel metal3 s 31600 50120 32000 50176 6 itasel[153]
port 995 nsew signal input
rlabel metal3 s 31600 50400 32000 50456 6 itasel[154]
port 996 nsew signal input
rlabel metal3 s 31600 50680 32000 50736 6 itasel[155]
port 997 nsew signal input
rlabel metal3 s 31600 50960 32000 51016 6 itasel[156]
port 998 nsew signal input
rlabel metal3 s 31600 51240 32000 51296 6 itasel[157]
port 999 nsew signal input
rlabel metal3 s 31600 51520 32000 51576 6 itasel[158]
port 1000 nsew signal input
rlabel metal3 s 31600 51800 32000 51856 6 itasel[159]
port 1001 nsew signal input
rlabel metal3 s 0 22680 400 22736 6 itasel[15]
port 1002 nsew signal input
rlabel metal3 s 31600 52080 32000 52136 6 itasel[160]
port 1003 nsew signal input
rlabel metal3 s 31600 52360 32000 52416 6 itasel[161]
port 1004 nsew signal input
rlabel metal3 s 31600 52640 32000 52696 6 itasel[162]
port 1005 nsew signal input
rlabel metal3 s 31600 52920 32000 52976 6 itasel[163]
port 1006 nsew signal input
rlabel metal3 s 31600 53200 32000 53256 6 itasel[164]
port 1007 nsew signal input
rlabel metal3 s 31600 53480 32000 53536 6 itasel[165]
port 1008 nsew signal input
rlabel metal3 s 31600 53760 32000 53816 6 itasel[166]
port 1009 nsew signal input
rlabel metal3 s 31600 54040 32000 54096 6 itasel[167]
port 1010 nsew signal input
rlabel metal3 s 31600 54320 32000 54376 6 itasel[168]
port 1011 nsew signal input
rlabel metal3 s 31600 54600 32000 54656 6 itasel[169]
port 1012 nsew signal input
rlabel metal3 s 0 22960 400 23016 6 itasel[16]
port 1013 nsew signal input
rlabel metal3 s 31600 54880 32000 54936 6 itasel[170]
port 1014 nsew signal input
rlabel metal3 s 31600 55160 32000 55216 6 itasel[171]
port 1015 nsew signal input
rlabel metal3 s 31600 55440 32000 55496 6 itasel[172]
port 1016 nsew signal input
rlabel metal3 s 31600 55720 32000 55776 6 itasel[173]
port 1017 nsew signal input
rlabel metal3 s 31600 56000 32000 56056 6 itasel[174]
port 1018 nsew signal input
rlabel metal3 s 31600 56280 32000 56336 6 itasel[175]
port 1019 nsew signal input
rlabel metal3 s 31600 56560 32000 56616 6 itasel[176]
port 1020 nsew signal input
rlabel metal3 s 31600 56840 32000 56896 6 itasel[177]
port 1021 nsew signal input
rlabel metal3 s 31600 57120 32000 57176 6 itasel[178]
port 1022 nsew signal input
rlabel metal3 s 31600 57400 32000 57456 6 itasel[179]
port 1023 nsew signal input
rlabel metal3 s 0 23240 400 23296 6 itasel[17]
port 1024 nsew signal input
rlabel metal3 s 31600 57680 32000 57736 6 itasel[180]
port 1025 nsew signal input
rlabel metal3 s 31600 57960 32000 58016 6 itasel[181]
port 1026 nsew signal input
rlabel metal3 s 31600 58240 32000 58296 6 itasel[182]
port 1027 nsew signal input
rlabel metal3 s 31600 58520 32000 58576 6 itasel[183]
port 1028 nsew signal input
rlabel metal3 s 31600 58800 32000 58856 6 itasel[184]
port 1029 nsew signal input
rlabel metal3 s 31600 59080 32000 59136 6 itasel[185]
port 1030 nsew signal input
rlabel metal3 s 31600 59360 32000 59416 6 itasel[186]
port 1031 nsew signal input
rlabel metal3 s 31600 59640 32000 59696 6 itasel[187]
port 1032 nsew signal input
rlabel metal3 s 31600 59920 32000 59976 6 itasel[188]
port 1033 nsew signal input
rlabel metal3 s 31600 60200 32000 60256 6 itasel[189]
port 1034 nsew signal input
rlabel metal3 s 0 23520 400 23576 6 itasel[18]
port 1035 nsew signal input
rlabel metal3 s 31600 60480 32000 60536 6 itasel[190]
port 1036 nsew signal input
rlabel metal3 s 31600 60760 32000 60816 6 itasel[191]
port 1037 nsew signal input
rlabel metal3 s 0 76720 400 76776 6 itasel[192]
port 1038 nsew signal input
rlabel metal3 s 0 77000 400 77056 6 itasel[193]
port 1039 nsew signal input
rlabel metal3 s 0 77280 400 77336 6 itasel[194]
port 1040 nsew signal input
rlabel metal3 s 0 77560 400 77616 6 itasel[195]
port 1041 nsew signal input
rlabel metal3 s 0 77840 400 77896 6 itasel[196]
port 1042 nsew signal input
rlabel metal3 s 0 78120 400 78176 6 itasel[197]
port 1043 nsew signal input
rlabel metal3 s 0 78400 400 78456 6 itasel[198]
port 1044 nsew signal input
rlabel metal3 s 0 78680 400 78736 6 itasel[199]
port 1045 nsew signal input
rlabel metal3 s 0 23800 400 23856 6 itasel[19]
port 1046 nsew signal input
rlabel metal3 s 0 18760 400 18816 6 itasel[1]
port 1047 nsew signal input
rlabel metal3 s 0 78960 400 79016 6 itasel[200]
port 1048 nsew signal input
rlabel metal3 s 0 79240 400 79296 6 itasel[201]
port 1049 nsew signal input
rlabel metal3 s 0 79520 400 79576 6 itasel[202]
port 1050 nsew signal input
rlabel metal3 s 0 79800 400 79856 6 itasel[203]
port 1051 nsew signal input
rlabel metal3 s 0 80080 400 80136 6 itasel[204]
port 1052 nsew signal input
rlabel metal3 s 0 80360 400 80416 6 itasel[205]
port 1053 nsew signal input
rlabel metal3 s 0 80640 400 80696 6 itasel[206]
port 1054 nsew signal input
rlabel metal3 s 0 80920 400 80976 6 itasel[207]
port 1055 nsew signal input
rlabel metal3 s 0 81200 400 81256 6 itasel[208]
port 1056 nsew signal input
rlabel metal3 s 0 81480 400 81536 6 itasel[209]
port 1057 nsew signal input
rlabel metal3 s 0 24080 400 24136 6 itasel[20]
port 1058 nsew signal input
rlabel metal3 s 0 81760 400 81816 6 itasel[210]
port 1059 nsew signal input
rlabel metal3 s 0 82040 400 82096 6 itasel[211]
port 1060 nsew signal input
rlabel metal3 s 0 82320 400 82376 6 itasel[212]
port 1061 nsew signal input
rlabel metal3 s 0 82600 400 82656 6 itasel[213]
port 1062 nsew signal input
rlabel metal3 s 0 82880 400 82936 6 itasel[214]
port 1063 nsew signal input
rlabel metal3 s 0 83160 400 83216 6 itasel[215]
port 1064 nsew signal input
rlabel metal3 s 0 83440 400 83496 6 itasel[216]
port 1065 nsew signal input
rlabel metal3 s 0 83720 400 83776 6 itasel[217]
port 1066 nsew signal input
rlabel metal3 s 0 84000 400 84056 6 itasel[218]
port 1067 nsew signal input
rlabel metal3 s 0 84280 400 84336 6 itasel[219]
port 1068 nsew signal input
rlabel metal3 s 0 24360 400 24416 6 itasel[21]
port 1069 nsew signal input
rlabel metal3 s 0 84560 400 84616 6 itasel[220]
port 1070 nsew signal input
rlabel metal3 s 0 84840 400 84896 6 itasel[221]
port 1071 nsew signal input
rlabel metal3 s 0 85120 400 85176 6 itasel[222]
port 1072 nsew signal input
rlabel metal3 s 0 85400 400 85456 6 itasel[223]
port 1073 nsew signal input
rlabel metal3 s 0 85680 400 85736 6 itasel[224]
port 1074 nsew signal input
rlabel metal3 s 0 85960 400 86016 6 itasel[225]
port 1075 nsew signal input
rlabel metal3 s 0 86240 400 86296 6 itasel[226]
port 1076 nsew signal input
rlabel metal3 s 0 86520 400 86576 6 itasel[227]
port 1077 nsew signal input
rlabel metal3 s 0 86800 400 86856 6 itasel[228]
port 1078 nsew signal input
rlabel metal3 s 0 87080 400 87136 6 itasel[229]
port 1079 nsew signal input
rlabel metal3 s 0 24640 400 24696 6 itasel[22]
port 1080 nsew signal input
rlabel metal3 s 0 87360 400 87416 6 itasel[230]
port 1081 nsew signal input
rlabel metal3 s 0 87640 400 87696 6 itasel[231]
port 1082 nsew signal input
rlabel metal3 s 0 87920 400 87976 6 itasel[232]
port 1083 nsew signal input
rlabel metal3 s 0 88200 400 88256 6 itasel[233]
port 1084 nsew signal input
rlabel metal3 s 0 88480 400 88536 6 itasel[234]
port 1085 nsew signal input
rlabel metal3 s 0 88760 400 88816 6 itasel[235]
port 1086 nsew signal input
rlabel metal3 s 0 89040 400 89096 6 itasel[236]
port 1087 nsew signal input
rlabel metal3 s 0 89320 400 89376 6 itasel[237]
port 1088 nsew signal input
rlabel metal3 s 0 89600 400 89656 6 itasel[238]
port 1089 nsew signal input
rlabel metal3 s 0 89880 400 89936 6 itasel[239]
port 1090 nsew signal input
rlabel metal3 s 0 24920 400 24976 6 itasel[23]
port 1091 nsew signal input
rlabel metal3 s 31600 76720 32000 76776 6 itasel[240]
port 1092 nsew signal input
rlabel metal3 s 31600 77000 32000 77056 6 itasel[241]
port 1093 nsew signal input
rlabel metal3 s 31600 77280 32000 77336 6 itasel[242]
port 1094 nsew signal input
rlabel metal3 s 31600 77560 32000 77616 6 itasel[243]
port 1095 nsew signal input
rlabel metal3 s 31600 77840 32000 77896 6 itasel[244]
port 1096 nsew signal input
rlabel metal3 s 31600 78120 32000 78176 6 itasel[245]
port 1097 nsew signal input
rlabel metal3 s 31600 78400 32000 78456 6 itasel[246]
port 1098 nsew signal input
rlabel metal3 s 31600 78680 32000 78736 6 itasel[247]
port 1099 nsew signal input
rlabel metal3 s 31600 78960 32000 79016 6 itasel[248]
port 1100 nsew signal input
rlabel metal3 s 31600 79240 32000 79296 6 itasel[249]
port 1101 nsew signal input
rlabel metal3 s 0 25200 400 25256 6 itasel[24]
port 1102 nsew signal input
rlabel metal3 s 31600 79520 32000 79576 6 itasel[250]
port 1103 nsew signal input
rlabel metal3 s 31600 79800 32000 79856 6 itasel[251]
port 1104 nsew signal input
rlabel metal3 s 31600 80080 32000 80136 6 itasel[252]
port 1105 nsew signal input
rlabel metal3 s 31600 80360 32000 80416 6 itasel[253]
port 1106 nsew signal input
rlabel metal3 s 31600 80640 32000 80696 6 itasel[254]
port 1107 nsew signal input
rlabel metal3 s 31600 80920 32000 80976 6 itasel[255]
port 1108 nsew signal input
rlabel metal3 s 31600 81200 32000 81256 6 itasel[256]
port 1109 nsew signal input
rlabel metal3 s 31600 81480 32000 81536 6 itasel[257]
port 1110 nsew signal input
rlabel metal3 s 31600 81760 32000 81816 6 itasel[258]
port 1111 nsew signal input
rlabel metal3 s 31600 82040 32000 82096 6 itasel[259]
port 1112 nsew signal input
rlabel metal3 s 0 25480 400 25536 6 itasel[25]
port 1113 nsew signal input
rlabel metal3 s 31600 82320 32000 82376 6 itasel[260]
port 1114 nsew signal input
rlabel metal3 s 31600 82600 32000 82656 6 itasel[261]
port 1115 nsew signal input
rlabel metal3 s 31600 82880 32000 82936 6 itasel[262]
port 1116 nsew signal input
rlabel metal3 s 31600 83160 32000 83216 6 itasel[263]
port 1117 nsew signal input
rlabel metal3 s 31600 83440 32000 83496 6 itasel[264]
port 1118 nsew signal input
rlabel metal3 s 31600 83720 32000 83776 6 itasel[265]
port 1119 nsew signal input
rlabel metal3 s 31600 84000 32000 84056 6 itasel[266]
port 1120 nsew signal input
rlabel metal3 s 31600 84280 32000 84336 6 itasel[267]
port 1121 nsew signal input
rlabel metal3 s 31600 84560 32000 84616 6 itasel[268]
port 1122 nsew signal input
rlabel metal3 s 31600 84840 32000 84896 6 itasel[269]
port 1123 nsew signal input
rlabel metal3 s 0 25760 400 25816 6 itasel[26]
port 1124 nsew signal input
rlabel metal3 s 31600 85120 32000 85176 6 itasel[270]
port 1125 nsew signal input
rlabel metal3 s 31600 85400 32000 85456 6 itasel[271]
port 1126 nsew signal input
rlabel metal3 s 31600 85680 32000 85736 6 itasel[272]
port 1127 nsew signal input
rlabel metal3 s 31600 85960 32000 86016 6 itasel[273]
port 1128 nsew signal input
rlabel metal3 s 31600 86240 32000 86296 6 itasel[274]
port 1129 nsew signal input
rlabel metal3 s 31600 86520 32000 86576 6 itasel[275]
port 1130 nsew signal input
rlabel metal3 s 31600 86800 32000 86856 6 itasel[276]
port 1131 nsew signal input
rlabel metal3 s 31600 87080 32000 87136 6 itasel[277]
port 1132 nsew signal input
rlabel metal3 s 31600 87360 32000 87416 6 itasel[278]
port 1133 nsew signal input
rlabel metal3 s 31600 87640 32000 87696 6 itasel[279]
port 1134 nsew signal input
rlabel metal3 s 0 26040 400 26096 6 itasel[27]
port 1135 nsew signal input
rlabel metal3 s 31600 87920 32000 87976 6 itasel[280]
port 1136 nsew signal input
rlabel metal3 s 31600 88200 32000 88256 6 itasel[281]
port 1137 nsew signal input
rlabel metal3 s 31600 88480 32000 88536 6 itasel[282]
port 1138 nsew signal input
rlabel metal3 s 31600 88760 32000 88816 6 itasel[283]
port 1139 nsew signal input
rlabel metal3 s 31600 89040 32000 89096 6 itasel[284]
port 1140 nsew signal input
rlabel metal3 s 31600 89320 32000 89376 6 itasel[285]
port 1141 nsew signal input
rlabel metal3 s 31600 89600 32000 89656 6 itasel[286]
port 1142 nsew signal input
rlabel metal3 s 31600 89880 32000 89936 6 itasel[287]
port 1143 nsew signal input
rlabel metal3 s 0 105840 400 105896 6 itasel[288]
port 1144 nsew signal input
rlabel metal3 s 0 106120 400 106176 6 itasel[289]
port 1145 nsew signal input
rlabel metal3 s 0 26320 400 26376 6 itasel[28]
port 1146 nsew signal input
rlabel metal3 s 0 106400 400 106456 6 itasel[290]
port 1147 nsew signal input
rlabel metal3 s 0 106680 400 106736 6 itasel[291]
port 1148 nsew signal input
rlabel metal3 s 0 106960 400 107016 6 itasel[292]
port 1149 nsew signal input
rlabel metal3 s 0 107240 400 107296 6 itasel[293]
port 1150 nsew signal input
rlabel metal3 s 0 107520 400 107576 6 itasel[294]
port 1151 nsew signal input
rlabel metal3 s 0 107800 400 107856 6 itasel[295]
port 1152 nsew signal input
rlabel metal3 s 0 108080 400 108136 6 itasel[296]
port 1153 nsew signal input
rlabel metal3 s 0 108360 400 108416 6 itasel[297]
port 1154 nsew signal input
rlabel metal3 s 0 108640 400 108696 6 itasel[298]
port 1155 nsew signal input
rlabel metal3 s 0 108920 400 108976 6 itasel[299]
port 1156 nsew signal input
rlabel metal3 s 0 26600 400 26656 6 itasel[29]
port 1157 nsew signal input
rlabel metal3 s 0 19040 400 19096 6 itasel[2]
port 1158 nsew signal input
rlabel metal3 s 0 109200 400 109256 6 itasel[300]
port 1159 nsew signal input
rlabel metal3 s 0 109480 400 109536 6 itasel[301]
port 1160 nsew signal input
rlabel metal3 s 0 109760 400 109816 6 itasel[302]
port 1161 nsew signal input
rlabel metal3 s 0 110040 400 110096 6 itasel[303]
port 1162 nsew signal input
rlabel metal3 s 0 110320 400 110376 6 itasel[304]
port 1163 nsew signal input
rlabel metal3 s 0 110600 400 110656 6 itasel[305]
port 1164 nsew signal input
rlabel metal3 s 0 110880 400 110936 6 itasel[306]
port 1165 nsew signal input
rlabel metal3 s 0 111160 400 111216 6 itasel[307]
port 1166 nsew signal input
rlabel metal3 s 0 111440 400 111496 6 itasel[308]
port 1167 nsew signal input
rlabel metal3 s 0 111720 400 111776 6 itasel[309]
port 1168 nsew signal input
rlabel metal3 s 0 26880 400 26936 6 itasel[30]
port 1169 nsew signal input
rlabel metal3 s 0 112000 400 112056 6 itasel[310]
port 1170 nsew signal input
rlabel metal3 s 0 112280 400 112336 6 itasel[311]
port 1171 nsew signal input
rlabel metal3 s 0 112560 400 112616 6 itasel[312]
port 1172 nsew signal input
rlabel metal3 s 0 112840 400 112896 6 itasel[313]
port 1173 nsew signal input
rlabel metal3 s 0 113120 400 113176 6 itasel[314]
port 1174 nsew signal input
rlabel metal3 s 0 113400 400 113456 6 itasel[315]
port 1175 nsew signal input
rlabel metal3 s 0 113680 400 113736 6 itasel[316]
port 1176 nsew signal input
rlabel metal3 s 0 113960 400 114016 6 itasel[317]
port 1177 nsew signal input
rlabel metal3 s 0 114240 400 114296 6 itasel[318]
port 1178 nsew signal input
rlabel metal3 s 0 114520 400 114576 6 itasel[319]
port 1179 nsew signal input
rlabel metal3 s 0 27160 400 27216 6 itasel[31]
port 1180 nsew signal input
rlabel metal3 s 0 114800 400 114856 6 itasel[320]
port 1181 nsew signal input
rlabel metal3 s 0 115080 400 115136 6 itasel[321]
port 1182 nsew signal input
rlabel metal3 s 0 115360 400 115416 6 itasel[322]
port 1183 nsew signal input
rlabel metal3 s 0 115640 400 115696 6 itasel[323]
port 1184 nsew signal input
rlabel metal3 s 0 115920 400 115976 6 itasel[324]
port 1185 nsew signal input
rlabel metal3 s 0 116200 400 116256 6 itasel[325]
port 1186 nsew signal input
rlabel metal3 s 0 116480 400 116536 6 itasel[326]
port 1187 nsew signal input
rlabel metal3 s 0 116760 400 116816 6 itasel[327]
port 1188 nsew signal input
rlabel metal3 s 0 117040 400 117096 6 itasel[328]
port 1189 nsew signal input
rlabel metal3 s 0 117320 400 117376 6 itasel[329]
port 1190 nsew signal input
rlabel metal3 s 0 27440 400 27496 6 itasel[32]
port 1191 nsew signal input
rlabel metal3 s 0 117600 400 117656 6 itasel[330]
port 1192 nsew signal input
rlabel metal3 s 0 117880 400 117936 6 itasel[331]
port 1193 nsew signal input
rlabel metal3 s 0 118160 400 118216 6 itasel[332]
port 1194 nsew signal input
rlabel metal3 s 0 118440 400 118496 6 itasel[333]
port 1195 nsew signal input
rlabel metal3 s 0 118720 400 118776 6 itasel[334]
port 1196 nsew signal input
rlabel metal3 s 0 119000 400 119056 6 itasel[335]
port 1197 nsew signal input
rlabel metal3 s 31600 105840 32000 105896 6 itasel[336]
port 1198 nsew signal input
rlabel metal3 s 31600 106120 32000 106176 6 itasel[337]
port 1199 nsew signal input
rlabel metal3 s 31600 106400 32000 106456 6 itasel[338]
port 1200 nsew signal input
rlabel metal3 s 31600 106680 32000 106736 6 itasel[339]
port 1201 nsew signal input
rlabel metal3 s 0 27720 400 27776 6 itasel[33]
port 1202 nsew signal input
rlabel metal3 s 31600 106960 32000 107016 6 itasel[340]
port 1203 nsew signal input
rlabel metal3 s 31600 107240 32000 107296 6 itasel[341]
port 1204 nsew signal input
rlabel metal3 s 31600 107520 32000 107576 6 itasel[342]
port 1205 nsew signal input
rlabel metal3 s 31600 107800 32000 107856 6 itasel[343]
port 1206 nsew signal input
rlabel metal3 s 31600 108080 32000 108136 6 itasel[344]
port 1207 nsew signal input
rlabel metal3 s 31600 108360 32000 108416 6 itasel[345]
port 1208 nsew signal input
rlabel metal3 s 31600 108640 32000 108696 6 itasel[346]
port 1209 nsew signal input
rlabel metal3 s 31600 108920 32000 108976 6 itasel[347]
port 1210 nsew signal input
rlabel metal3 s 31600 109200 32000 109256 6 itasel[348]
port 1211 nsew signal input
rlabel metal3 s 31600 109480 32000 109536 6 itasel[349]
port 1212 nsew signal input
rlabel metal3 s 0 28000 400 28056 6 itasel[34]
port 1213 nsew signal input
rlabel metal3 s 31600 109760 32000 109816 6 itasel[350]
port 1214 nsew signal input
rlabel metal3 s 31600 110040 32000 110096 6 itasel[351]
port 1215 nsew signal input
rlabel metal3 s 31600 110320 32000 110376 6 itasel[352]
port 1216 nsew signal input
rlabel metal3 s 31600 110600 32000 110656 6 itasel[353]
port 1217 nsew signal input
rlabel metal3 s 31600 110880 32000 110936 6 itasel[354]
port 1218 nsew signal input
rlabel metal3 s 31600 111160 32000 111216 6 itasel[355]
port 1219 nsew signal input
rlabel metal3 s 31600 111440 32000 111496 6 itasel[356]
port 1220 nsew signal input
rlabel metal3 s 31600 111720 32000 111776 6 itasel[357]
port 1221 nsew signal input
rlabel metal3 s 31600 112000 32000 112056 6 itasel[358]
port 1222 nsew signal input
rlabel metal3 s 31600 112280 32000 112336 6 itasel[359]
port 1223 nsew signal input
rlabel metal3 s 0 28280 400 28336 6 itasel[35]
port 1224 nsew signal input
rlabel metal3 s 31600 112560 32000 112616 6 itasel[360]
port 1225 nsew signal input
rlabel metal3 s 31600 112840 32000 112896 6 itasel[361]
port 1226 nsew signal input
rlabel metal3 s 31600 113120 32000 113176 6 itasel[362]
port 1227 nsew signal input
rlabel metal3 s 31600 113400 32000 113456 6 itasel[363]
port 1228 nsew signal input
rlabel metal3 s 31600 113680 32000 113736 6 itasel[364]
port 1229 nsew signal input
rlabel metal3 s 31600 113960 32000 114016 6 itasel[365]
port 1230 nsew signal input
rlabel metal3 s 31600 114240 32000 114296 6 itasel[366]
port 1231 nsew signal input
rlabel metal3 s 31600 114520 32000 114576 6 itasel[367]
port 1232 nsew signal input
rlabel metal3 s 31600 114800 32000 114856 6 itasel[368]
port 1233 nsew signal input
rlabel metal3 s 31600 115080 32000 115136 6 itasel[369]
port 1234 nsew signal input
rlabel metal3 s 0 28560 400 28616 6 itasel[36]
port 1235 nsew signal input
rlabel metal3 s 31600 115360 32000 115416 6 itasel[370]
port 1236 nsew signal input
rlabel metal3 s 31600 115640 32000 115696 6 itasel[371]
port 1237 nsew signal input
rlabel metal3 s 31600 115920 32000 115976 6 itasel[372]
port 1238 nsew signal input
rlabel metal3 s 31600 116200 32000 116256 6 itasel[373]
port 1239 nsew signal input
rlabel metal3 s 31600 116480 32000 116536 6 itasel[374]
port 1240 nsew signal input
rlabel metal3 s 31600 116760 32000 116816 6 itasel[375]
port 1241 nsew signal input
rlabel metal3 s 31600 117040 32000 117096 6 itasel[376]
port 1242 nsew signal input
rlabel metal3 s 31600 117320 32000 117376 6 itasel[377]
port 1243 nsew signal input
rlabel metal3 s 31600 117600 32000 117656 6 itasel[378]
port 1244 nsew signal input
rlabel metal3 s 31600 117880 32000 117936 6 itasel[379]
port 1245 nsew signal input
rlabel metal3 s 0 28840 400 28896 6 itasel[37]
port 1246 nsew signal input
rlabel metal3 s 31600 118160 32000 118216 6 itasel[380]
port 1247 nsew signal input
rlabel metal3 s 31600 118440 32000 118496 6 itasel[381]
port 1248 nsew signal input
rlabel metal3 s 31600 118720 32000 118776 6 itasel[382]
port 1249 nsew signal input
rlabel metal3 s 31600 119000 32000 119056 6 itasel[383]
port 1250 nsew signal input
rlabel metal3 s 0 134960 400 135016 6 itasel[384]
port 1251 nsew signal input
rlabel metal3 s 0 135240 400 135296 6 itasel[385]
port 1252 nsew signal input
rlabel metal3 s 0 135520 400 135576 6 itasel[386]
port 1253 nsew signal input
rlabel metal3 s 0 135800 400 135856 6 itasel[387]
port 1254 nsew signal input
rlabel metal3 s 0 136080 400 136136 6 itasel[388]
port 1255 nsew signal input
rlabel metal3 s 0 136360 400 136416 6 itasel[389]
port 1256 nsew signal input
rlabel metal3 s 0 29120 400 29176 6 itasel[38]
port 1257 nsew signal input
rlabel metal3 s 0 136640 400 136696 6 itasel[390]
port 1258 nsew signal input
rlabel metal3 s 0 136920 400 136976 6 itasel[391]
port 1259 nsew signal input
rlabel metal3 s 0 137200 400 137256 6 itasel[392]
port 1260 nsew signal input
rlabel metal3 s 0 137480 400 137536 6 itasel[393]
port 1261 nsew signal input
rlabel metal3 s 0 137760 400 137816 6 itasel[394]
port 1262 nsew signal input
rlabel metal3 s 0 138040 400 138096 6 itasel[395]
port 1263 nsew signal input
rlabel metal3 s 0 138320 400 138376 6 itasel[396]
port 1264 nsew signal input
rlabel metal3 s 0 138600 400 138656 6 itasel[397]
port 1265 nsew signal input
rlabel metal3 s 0 138880 400 138936 6 itasel[398]
port 1266 nsew signal input
rlabel metal3 s 0 139160 400 139216 6 itasel[399]
port 1267 nsew signal input
rlabel metal3 s 0 29400 400 29456 6 itasel[39]
port 1268 nsew signal input
rlabel metal3 s 0 19320 400 19376 6 itasel[3]
port 1269 nsew signal input
rlabel metal3 s 0 139440 400 139496 6 itasel[400]
port 1270 nsew signal input
rlabel metal3 s 0 139720 400 139776 6 itasel[401]
port 1271 nsew signal input
rlabel metal3 s 0 140000 400 140056 6 itasel[402]
port 1272 nsew signal input
rlabel metal3 s 0 140280 400 140336 6 itasel[403]
port 1273 nsew signal input
rlabel metal3 s 0 140560 400 140616 6 itasel[404]
port 1274 nsew signal input
rlabel metal3 s 0 140840 400 140896 6 itasel[405]
port 1275 nsew signal input
rlabel metal3 s 0 141120 400 141176 6 itasel[406]
port 1276 nsew signal input
rlabel metal3 s 0 141400 400 141456 6 itasel[407]
port 1277 nsew signal input
rlabel metal3 s 0 141680 400 141736 6 itasel[408]
port 1278 nsew signal input
rlabel metal3 s 0 141960 400 142016 6 itasel[409]
port 1279 nsew signal input
rlabel metal3 s 0 29680 400 29736 6 itasel[40]
port 1280 nsew signal input
rlabel metal3 s 0 142240 400 142296 6 itasel[410]
port 1281 nsew signal input
rlabel metal3 s 0 142520 400 142576 6 itasel[411]
port 1282 nsew signal input
rlabel metal3 s 0 142800 400 142856 6 itasel[412]
port 1283 nsew signal input
rlabel metal3 s 0 143080 400 143136 6 itasel[413]
port 1284 nsew signal input
rlabel metal3 s 0 143360 400 143416 6 itasel[414]
port 1285 nsew signal input
rlabel metal3 s 0 143640 400 143696 6 itasel[415]
port 1286 nsew signal input
rlabel metal3 s 0 143920 400 143976 6 itasel[416]
port 1287 nsew signal input
rlabel metal3 s 0 144200 400 144256 6 itasel[417]
port 1288 nsew signal input
rlabel metal3 s 0 144480 400 144536 6 itasel[418]
port 1289 nsew signal input
rlabel metal3 s 0 144760 400 144816 6 itasel[419]
port 1290 nsew signal input
rlabel metal3 s 0 29960 400 30016 6 itasel[41]
port 1291 nsew signal input
rlabel metal3 s 0 145040 400 145096 6 itasel[420]
port 1292 nsew signal input
rlabel metal3 s 0 145320 400 145376 6 itasel[421]
port 1293 nsew signal input
rlabel metal3 s 0 145600 400 145656 6 itasel[422]
port 1294 nsew signal input
rlabel metal3 s 0 145880 400 145936 6 itasel[423]
port 1295 nsew signal input
rlabel metal3 s 0 146160 400 146216 6 itasel[424]
port 1296 nsew signal input
rlabel metal3 s 0 146440 400 146496 6 itasel[425]
port 1297 nsew signal input
rlabel metal3 s 0 146720 400 146776 6 itasel[426]
port 1298 nsew signal input
rlabel metal3 s 0 147000 400 147056 6 itasel[427]
port 1299 nsew signal input
rlabel metal3 s 0 147280 400 147336 6 itasel[428]
port 1300 nsew signal input
rlabel metal3 s 0 147560 400 147616 6 itasel[429]
port 1301 nsew signal input
rlabel metal3 s 0 30240 400 30296 6 itasel[42]
port 1302 nsew signal input
rlabel metal3 s 0 147840 400 147896 6 itasel[430]
port 1303 nsew signal input
rlabel metal3 s 0 148120 400 148176 6 itasel[431]
port 1304 nsew signal input
rlabel metal3 s 31600 134960 32000 135016 6 itasel[432]
port 1305 nsew signal input
rlabel metal3 s 31600 135240 32000 135296 6 itasel[433]
port 1306 nsew signal input
rlabel metal3 s 31600 135520 32000 135576 6 itasel[434]
port 1307 nsew signal input
rlabel metal3 s 31600 135800 32000 135856 6 itasel[435]
port 1308 nsew signal input
rlabel metal3 s 31600 136080 32000 136136 6 itasel[436]
port 1309 nsew signal input
rlabel metal3 s 31600 136360 32000 136416 6 itasel[437]
port 1310 nsew signal input
rlabel metal3 s 31600 136640 32000 136696 6 itasel[438]
port 1311 nsew signal input
rlabel metal3 s 31600 136920 32000 136976 6 itasel[439]
port 1312 nsew signal input
rlabel metal3 s 0 30520 400 30576 6 itasel[43]
port 1313 nsew signal input
rlabel metal3 s 31600 137200 32000 137256 6 itasel[440]
port 1314 nsew signal input
rlabel metal3 s 31600 137480 32000 137536 6 itasel[441]
port 1315 nsew signal input
rlabel metal3 s 31600 137760 32000 137816 6 itasel[442]
port 1316 nsew signal input
rlabel metal3 s 31600 138040 32000 138096 6 itasel[443]
port 1317 nsew signal input
rlabel metal3 s 31600 138320 32000 138376 6 itasel[444]
port 1318 nsew signal input
rlabel metal3 s 31600 138600 32000 138656 6 itasel[445]
port 1319 nsew signal input
rlabel metal3 s 31600 138880 32000 138936 6 itasel[446]
port 1320 nsew signal input
rlabel metal3 s 31600 139160 32000 139216 6 itasel[447]
port 1321 nsew signal input
rlabel metal3 s 31600 139440 32000 139496 6 itasel[448]
port 1322 nsew signal input
rlabel metal3 s 31600 139720 32000 139776 6 itasel[449]
port 1323 nsew signal input
rlabel metal3 s 0 30800 400 30856 6 itasel[44]
port 1324 nsew signal input
rlabel metal3 s 31600 140000 32000 140056 6 itasel[450]
port 1325 nsew signal input
rlabel metal3 s 31600 140280 32000 140336 6 itasel[451]
port 1326 nsew signal input
rlabel metal3 s 31600 140560 32000 140616 6 itasel[452]
port 1327 nsew signal input
rlabel metal3 s 31600 140840 32000 140896 6 itasel[453]
port 1328 nsew signal input
rlabel metal3 s 31600 141120 32000 141176 6 itasel[454]
port 1329 nsew signal input
rlabel metal3 s 31600 141400 32000 141456 6 itasel[455]
port 1330 nsew signal input
rlabel metal3 s 31600 141680 32000 141736 6 itasel[456]
port 1331 nsew signal input
rlabel metal3 s 31600 141960 32000 142016 6 itasel[457]
port 1332 nsew signal input
rlabel metal3 s 31600 142240 32000 142296 6 itasel[458]
port 1333 nsew signal input
rlabel metal3 s 31600 142520 32000 142576 6 itasel[459]
port 1334 nsew signal input
rlabel metal3 s 0 31080 400 31136 6 itasel[45]
port 1335 nsew signal input
rlabel metal3 s 31600 142800 32000 142856 6 itasel[460]
port 1336 nsew signal input
rlabel metal3 s 31600 143080 32000 143136 6 itasel[461]
port 1337 nsew signal input
rlabel metal3 s 31600 143360 32000 143416 6 itasel[462]
port 1338 nsew signal input
rlabel metal3 s 31600 143640 32000 143696 6 itasel[463]
port 1339 nsew signal input
rlabel metal3 s 31600 143920 32000 143976 6 itasel[464]
port 1340 nsew signal input
rlabel metal3 s 31600 144200 32000 144256 6 itasel[465]
port 1341 nsew signal input
rlabel metal3 s 31600 144480 32000 144536 6 itasel[466]
port 1342 nsew signal input
rlabel metal3 s 31600 144760 32000 144816 6 itasel[467]
port 1343 nsew signal input
rlabel metal3 s 31600 145040 32000 145096 6 itasel[468]
port 1344 nsew signal input
rlabel metal3 s 31600 145320 32000 145376 6 itasel[469]
port 1345 nsew signal input
rlabel metal3 s 0 31360 400 31416 6 itasel[46]
port 1346 nsew signal input
rlabel metal3 s 31600 145600 32000 145656 6 itasel[470]
port 1347 nsew signal input
rlabel metal3 s 31600 145880 32000 145936 6 itasel[471]
port 1348 nsew signal input
rlabel metal3 s 31600 146160 32000 146216 6 itasel[472]
port 1349 nsew signal input
rlabel metal3 s 31600 146440 32000 146496 6 itasel[473]
port 1350 nsew signal input
rlabel metal3 s 31600 146720 32000 146776 6 itasel[474]
port 1351 nsew signal input
rlabel metal3 s 31600 147000 32000 147056 6 itasel[475]
port 1352 nsew signal input
rlabel metal3 s 31600 147280 32000 147336 6 itasel[476]
port 1353 nsew signal input
rlabel metal3 s 31600 147560 32000 147616 6 itasel[477]
port 1354 nsew signal input
rlabel metal3 s 31600 147840 32000 147896 6 itasel[478]
port 1355 nsew signal input
rlabel metal3 s 31600 148120 32000 148176 6 itasel[479]
port 1356 nsew signal input
rlabel metal3 s 0 31640 400 31696 6 itasel[47]
port 1357 nsew signal input
rlabel metal3 s 0 164080 400 164136 6 itasel[480]
port 1358 nsew signal input
rlabel metal3 s 0 164360 400 164416 6 itasel[481]
port 1359 nsew signal input
rlabel metal3 s 0 164640 400 164696 6 itasel[482]
port 1360 nsew signal input
rlabel metal3 s 0 164920 400 164976 6 itasel[483]
port 1361 nsew signal input
rlabel metal3 s 0 165200 400 165256 6 itasel[484]
port 1362 nsew signal input
rlabel metal3 s 0 165480 400 165536 6 itasel[485]
port 1363 nsew signal input
rlabel metal3 s 0 165760 400 165816 6 itasel[486]
port 1364 nsew signal input
rlabel metal3 s 0 166040 400 166096 6 itasel[487]
port 1365 nsew signal input
rlabel metal3 s 0 166320 400 166376 6 itasel[488]
port 1366 nsew signal input
rlabel metal3 s 0 166600 400 166656 6 itasel[489]
port 1367 nsew signal input
rlabel metal3 s 31600 18480 32000 18536 6 itasel[48]
port 1368 nsew signal input
rlabel metal3 s 0 166880 400 166936 6 itasel[490]
port 1369 nsew signal input
rlabel metal3 s 0 167160 400 167216 6 itasel[491]
port 1370 nsew signal input
rlabel metal3 s 0 167440 400 167496 6 itasel[492]
port 1371 nsew signal input
rlabel metal3 s 0 167720 400 167776 6 itasel[493]
port 1372 nsew signal input
rlabel metal3 s 0 168000 400 168056 6 itasel[494]
port 1373 nsew signal input
rlabel metal3 s 0 168280 400 168336 6 itasel[495]
port 1374 nsew signal input
rlabel metal3 s 0 168560 400 168616 6 itasel[496]
port 1375 nsew signal input
rlabel metal3 s 0 168840 400 168896 6 itasel[497]
port 1376 nsew signal input
rlabel metal3 s 0 169120 400 169176 6 itasel[498]
port 1377 nsew signal input
rlabel metal3 s 0 169400 400 169456 6 itasel[499]
port 1378 nsew signal input
rlabel metal3 s 31600 18760 32000 18816 6 itasel[49]
port 1379 nsew signal input
rlabel metal3 s 0 19600 400 19656 6 itasel[4]
port 1380 nsew signal input
rlabel metal3 s 0 169680 400 169736 6 itasel[500]
port 1381 nsew signal input
rlabel metal3 s 0 169960 400 170016 6 itasel[501]
port 1382 nsew signal input
rlabel metal3 s 0 170240 400 170296 6 itasel[502]
port 1383 nsew signal input
rlabel metal3 s 0 170520 400 170576 6 itasel[503]
port 1384 nsew signal input
rlabel metal3 s 0 170800 400 170856 6 itasel[504]
port 1385 nsew signal input
rlabel metal3 s 0 171080 400 171136 6 itasel[505]
port 1386 nsew signal input
rlabel metal3 s 0 171360 400 171416 6 itasel[506]
port 1387 nsew signal input
rlabel metal3 s 0 171640 400 171696 6 itasel[507]
port 1388 nsew signal input
rlabel metal3 s 0 171920 400 171976 6 itasel[508]
port 1389 nsew signal input
rlabel metal3 s 0 172200 400 172256 6 itasel[509]
port 1390 nsew signal input
rlabel metal3 s 31600 19040 32000 19096 6 itasel[50]
port 1391 nsew signal input
rlabel metal3 s 0 172480 400 172536 6 itasel[510]
port 1392 nsew signal input
rlabel metal3 s 0 172760 400 172816 6 itasel[511]
port 1393 nsew signal input
rlabel metal3 s 0 173040 400 173096 6 itasel[512]
port 1394 nsew signal input
rlabel metal3 s 0 173320 400 173376 6 itasel[513]
port 1395 nsew signal input
rlabel metal3 s 0 173600 400 173656 6 itasel[514]
port 1396 nsew signal input
rlabel metal3 s 0 173880 400 173936 6 itasel[515]
port 1397 nsew signal input
rlabel metal3 s 0 174160 400 174216 6 itasel[516]
port 1398 nsew signal input
rlabel metal3 s 0 174440 400 174496 6 itasel[517]
port 1399 nsew signal input
rlabel metal3 s 0 174720 400 174776 6 itasel[518]
port 1400 nsew signal input
rlabel metal3 s 0 175000 400 175056 6 itasel[519]
port 1401 nsew signal input
rlabel metal3 s 31600 19320 32000 19376 6 itasel[51]
port 1402 nsew signal input
rlabel metal3 s 0 175280 400 175336 6 itasel[520]
port 1403 nsew signal input
rlabel metal3 s 0 175560 400 175616 6 itasel[521]
port 1404 nsew signal input
rlabel metal3 s 0 175840 400 175896 6 itasel[522]
port 1405 nsew signal input
rlabel metal3 s 0 176120 400 176176 6 itasel[523]
port 1406 nsew signal input
rlabel metal3 s 0 176400 400 176456 6 itasel[524]
port 1407 nsew signal input
rlabel metal3 s 0 176680 400 176736 6 itasel[525]
port 1408 nsew signal input
rlabel metal3 s 0 176960 400 177016 6 itasel[526]
port 1409 nsew signal input
rlabel metal3 s 0 177240 400 177296 6 itasel[527]
port 1410 nsew signal input
rlabel metal3 s 31600 164080 32000 164136 6 itasel[528]
port 1411 nsew signal input
rlabel metal3 s 31600 164360 32000 164416 6 itasel[529]
port 1412 nsew signal input
rlabel metal3 s 31600 19600 32000 19656 6 itasel[52]
port 1413 nsew signal input
rlabel metal3 s 31600 164640 32000 164696 6 itasel[530]
port 1414 nsew signal input
rlabel metal3 s 31600 164920 32000 164976 6 itasel[531]
port 1415 nsew signal input
rlabel metal3 s 31600 165200 32000 165256 6 itasel[532]
port 1416 nsew signal input
rlabel metal3 s 31600 165480 32000 165536 6 itasel[533]
port 1417 nsew signal input
rlabel metal3 s 31600 165760 32000 165816 6 itasel[534]
port 1418 nsew signal input
rlabel metal3 s 31600 166040 32000 166096 6 itasel[535]
port 1419 nsew signal input
rlabel metal3 s 31600 166320 32000 166376 6 itasel[536]
port 1420 nsew signal input
rlabel metal3 s 31600 166600 32000 166656 6 itasel[537]
port 1421 nsew signal input
rlabel metal3 s 31600 166880 32000 166936 6 itasel[538]
port 1422 nsew signal input
rlabel metal3 s 31600 167160 32000 167216 6 itasel[539]
port 1423 nsew signal input
rlabel metal3 s 31600 19880 32000 19936 6 itasel[53]
port 1424 nsew signal input
rlabel metal3 s 31600 167440 32000 167496 6 itasel[540]
port 1425 nsew signal input
rlabel metal3 s 31600 167720 32000 167776 6 itasel[541]
port 1426 nsew signal input
rlabel metal3 s 31600 168000 32000 168056 6 itasel[542]
port 1427 nsew signal input
rlabel metal3 s 31600 168280 32000 168336 6 itasel[543]
port 1428 nsew signal input
rlabel metal3 s 31600 168560 32000 168616 6 itasel[544]
port 1429 nsew signal input
rlabel metal3 s 31600 168840 32000 168896 6 itasel[545]
port 1430 nsew signal input
rlabel metal3 s 31600 169120 32000 169176 6 itasel[546]
port 1431 nsew signal input
rlabel metal3 s 31600 169400 32000 169456 6 itasel[547]
port 1432 nsew signal input
rlabel metal3 s 31600 169680 32000 169736 6 itasel[548]
port 1433 nsew signal input
rlabel metal3 s 31600 169960 32000 170016 6 itasel[549]
port 1434 nsew signal input
rlabel metal3 s 31600 20160 32000 20216 6 itasel[54]
port 1435 nsew signal input
rlabel metal3 s 31600 170240 32000 170296 6 itasel[550]
port 1436 nsew signal input
rlabel metal3 s 31600 170520 32000 170576 6 itasel[551]
port 1437 nsew signal input
rlabel metal3 s 31600 170800 32000 170856 6 itasel[552]
port 1438 nsew signal input
rlabel metal3 s 31600 171080 32000 171136 6 itasel[553]
port 1439 nsew signal input
rlabel metal3 s 31600 171360 32000 171416 6 itasel[554]
port 1440 nsew signal input
rlabel metal3 s 31600 171640 32000 171696 6 itasel[555]
port 1441 nsew signal input
rlabel metal3 s 31600 171920 32000 171976 6 itasel[556]
port 1442 nsew signal input
rlabel metal3 s 31600 172200 32000 172256 6 itasel[557]
port 1443 nsew signal input
rlabel metal3 s 31600 172480 32000 172536 6 itasel[558]
port 1444 nsew signal input
rlabel metal3 s 31600 172760 32000 172816 6 itasel[559]
port 1445 nsew signal input
rlabel metal3 s 31600 20440 32000 20496 6 itasel[55]
port 1446 nsew signal input
rlabel metal3 s 31600 173040 32000 173096 6 itasel[560]
port 1447 nsew signal input
rlabel metal3 s 31600 173320 32000 173376 6 itasel[561]
port 1448 nsew signal input
rlabel metal3 s 31600 173600 32000 173656 6 itasel[562]
port 1449 nsew signal input
rlabel metal3 s 31600 173880 32000 173936 6 itasel[563]
port 1450 nsew signal input
rlabel metal3 s 31600 174160 32000 174216 6 itasel[564]
port 1451 nsew signal input
rlabel metal3 s 31600 174440 32000 174496 6 itasel[565]
port 1452 nsew signal input
rlabel metal3 s 31600 174720 32000 174776 6 itasel[566]
port 1453 nsew signal input
rlabel metal3 s 31600 175000 32000 175056 6 itasel[567]
port 1454 nsew signal input
rlabel metal3 s 31600 175280 32000 175336 6 itasel[568]
port 1455 nsew signal input
rlabel metal3 s 31600 175560 32000 175616 6 itasel[569]
port 1456 nsew signal input
rlabel metal3 s 31600 20720 32000 20776 6 itasel[56]
port 1457 nsew signal input
rlabel metal3 s 31600 175840 32000 175896 6 itasel[570]
port 1458 nsew signal input
rlabel metal3 s 31600 176120 32000 176176 6 itasel[571]
port 1459 nsew signal input
rlabel metal3 s 31600 176400 32000 176456 6 itasel[572]
port 1460 nsew signal input
rlabel metal3 s 31600 176680 32000 176736 6 itasel[573]
port 1461 nsew signal input
rlabel metal3 s 31600 176960 32000 177016 6 itasel[574]
port 1462 nsew signal input
rlabel metal3 s 31600 177240 32000 177296 6 itasel[575]
port 1463 nsew signal input
rlabel metal3 s 0 193200 400 193256 6 itasel[576]
port 1464 nsew signal input
rlabel metal3 s 0 193480 400 193536 6 itasel[577]
port 1465 nsew signal input
rlabel metal3 s 0 193760 400 193816 6 itasel[578]
port 1466 nsew signal input
rlabel metal3 s 0 194040 400 194096 6 itasel[579]
port 1467 nsew signal input
rlabel metal3 s 31600 21000 32000 21056 6 itasel[57]
port 1468 nsew signal input
rlabel metal3 s 0 194320 400 194376 6 itasel[580]
port 1469 nsew signal input
rlabel metal3 s 0 194600 400 194656 6 itasel[581]
port 1470 nsew signal input
rlabel metal3 s 0 194880 400 194936 6 itasel[582]
port 1471 nsew signal input
rlabel metal3 s 0 195160 400 195216 6 itasel[583]
port 1472 nsew signal input
rlabel metal3 s 0 195440 400 195496 6 itasel[584]
port 1473 nsew signal input
rlabel metal3 s 0 195720 400 195776 6 itasel[585]
port 1474 nsew signal input
rlabel metal3 s 0 196000 400 196056 6 itasel[586]
port 1475 nsew signal input
rlabel metal3 s 0 196280 400 196336 6 itasel[587]
port 1476 nsew signal input
rlabel metal3 s 0 196560 400 196616 6 itasel[588]
port 1477 nsew signal input
rlabel metal3 s 0 196840 400 196896 6 itasel[589]
port 1478 nsew signal input
rlabel metal3 s 31600 21280 32000 21336 6 itasel[58]
port 1479 nsew signal input
rlabel metal3 s 0 197120 400 197176 6 itasel[590]
port 1480 nsew signal input
rlabel metal3 s 0 197400 400 197456 6 itasel[591]
port 1481 nsew signal input
rlabel metal3 s 0 197680 400 197736 6 itasel[592]
port 1482 nsew signal input
rlabel metal3 s 0 197960 400 198016 6 itasel[593]
port 1483 nsew signal input
rlabel metal3 s 0 198240 400 198296 6 itasel[594]
port 1484 nsew signal input
rlabel metal3 s 0 198520 400 198576 6 itasel[595]
port 1485 nsew signal input
rlabel metal3 s 0 198800 400 198856 6 itasel[596]
port 1486 nsew signal input
rlabel metal3 s 0 199080 400 199136 6 itasel[597]
port 1487 nsew signal input
rlabel metal3 s 0 199360 400 199416 6 itasel[598]
port 1488 nsew signal input
rlabel metal3 s 0 199640 400 199696 6 itasel[599]
port 1489 nsew signal input
rlabel metal3 s 31600 21560 32000 21616 6 itasel[59]
port 1490 nsew signal input
rlabel metal3 s 0 19880 400 19936 6 itasel[5]
port 1491 nsew signal input
rlabel metal3 s 0 199920 400 199976 6 itasel[600]
port 1492 nsew signal input
rlabel metal3 s 0 200200 400 200256 6 itasel[601]
port 1493 nsew signal input
rlabel metal3 s 0 200480 400 200536 6 itasel[602]
port 1494 nsew signal input
rlabel metal3 s 0 200760 400 200816 6 itasel[603]
port 1495 nsew signal input
rlabel metal3 s 0 201040 400 201096 6 itasel[604]
port 1496 nsew signal input
rlabel metal3 s 0 201320 400 201376 6 itasel[605]
port 1497 nsew signal input
rlabel metal3 s 0 201600 400 201656 6 itasel[606]
port 1498 nsew signal input
rlabel metal3 s 0 201880 400 201936 6 itasel[607]
port 1499 nsew signal input
rlabel metal3 s 0 202160 400 202216 6 itasel[608]
port 1500 nsew signal input
rlabel metal3 s 0 202440 400 202496 6 itasel[609]
port 1501 nsew signal input
rlabel metal3 s 31600 21840 32000 21896 6 itasel[60]
port 1502 nsew signal input
rlabel metal3 s 0 202720 400 202776 6 itasel[610]
port 1503 nsew signal input
rlabel metal3 s 0 203000 400 203056 6 itasel[611]
port 1504 nsew signal input
rlabel metal3 s 0 203280 400 203336 6 itasel[612]
port 1505 nsew signal input
rlabel metal3 s 0 203560 400 203616 6 itasel[613]
port 1506 nsew signal input
rlabel metal3 s 0 203840 400 203896 6 itasel[614]
port 1507 nsew signal input
rlabel metal3 s 0 204120 400 204176 6 itasel[615]
port 1508 nsew signal input
rlabel metal3 s 0 204400 400 204456 6 itasel[616]
port 1509 nsew signal input
rlabel metal3 s 0 204680 400 204736 6 itasel[617]
port 1510 nsew signal input
rlabel metal3 s 0 204960 400 205016 6 itasel[618]
port 1511 nsew signal input
rlabel metal3 s 0 205240 400 205296 6 itasel[619]
port 1512 nsew signal input
rlabel metal3 s 31600 22120 32000 22176 6 itasel[61]
port 1513 nsew signal input
rlabel metal3 s 0 205520 400 205576 6 itasel[620]
port 1514 nsew signal input
rlabel metal3 s 0 205800 400 205856 6 itasel[621]
port 1515 nsew signal input
rlabel metal3 s 0 206080 400 206136 6 itasel[622]
port 1516 nsew signal input
rlabel metal3 s 0 206360 400 206416 6 itasel[623]
port 1517 nsew signal input
rlabel metal3 s 31600 193200 32000 193256 6 itasel[624]
port 1518 nsew signal input
rlabel metal3 s 31600 193480 32000 193536 6 itasel[625]
port 1519 nsew signal input
rlabel metal3 s 31600 193760 32000 193816 6 itasel[626]
port 1520 nsew signal input
rlabel metal3 s 31600 194040 32000 194096 6 itasel[627]
port 1521 nsew signal input
rlabel metal3 s 31600 194320 32000 194376 6 itasel[628]
port 1522 nsew signal input
rlabel metal3 s 31600 194600 32000 194656 6 itasel[629]
port 1523 nsew signal input
rlabel metal3 s 31600 22400 32000 22456 6 itasel[62]
port 1524 nsew signal input
rlabel metal3 s 31600 194880 32000 194936 6 itasel[630]
port 1525 nsew signal input
rlabel metal3 s 31600 195160 32000 195216 6 itasel[631]
port 1526 nsew signal input
rlabel metal3 s 31600 195440 32000 195496 6 itasel[632]
port 1527 nsew signal input
rlabel metal3 s 31600 195720 32000 195776 6 itasel[633]
port 1528 nsew signal input
rlabel metal3 s 31600 196000 32000 196056 6 itasel[634]
port 1529 nsew signal input
rlabel metal3 s 31600 196280 32000 196336 6 itasel[635]
port 1530 nsew signal input
rlabel metal3 s 31600 196560 32000 196616 6 itasel[636]
port 1531 nsew signal input
rlabel metal3 s 31600 196840 32000 196896 6 itasel[637]
port 1532 nsew signal input
rlabel metal3 s 31600 197120 32000 197176 6 itasel[638]
port 1533 nsew signal input
rlabel metal3 s 31600 197400 32000 197456 6 itasel[639]
port 1534 nsew signal input
rlabel metal3 s 31600 22680 32000 22736 6 itasel[63]
port 1535 nsew signal input
rlabel metal3 s 31600 197680 32000 197736 6 itasel[640]
port 1536 nsew signal input
rlabel metal3 s 31600 197960 32000 198016 6 itasel[641]
port 1537 nsew signal input
rlabel metal3 s 31600 198240 32000 198296 6 itasel[642]
port 1538 nsew signal input
rlabel metal3 s 31600 198520 32000 198576 6 itasel[643]
port 1539 nsew signal input
rlabel metal3 s 31600 198800 32000 198856 6 itasel[644]
port 1540 nsew signal input
rlabel metal3 s 31600 199080 32000 199136 6 itasel[645]
port 1541 nsew signal input
rlabel metal3 s 31600 199360 32000 199416 6 itasel[646]
port 1542 nsew signal input
rlabel metal3 s 31600 199640 32000 199696 6 itasel[647]
port 1543 nsew signal input
rlabel metal3 s 31600 199920 32000 199976 6 itasel[648]
port 1544 nsew signal input
rlabel metal3 s 31600 200200 32000 200256 6 itasel[649]
port 1545 nsew signal input
rlabel metal3 s 31600 22960 32000 23016 6 itasel[64]
port 1546 nsew signal input
rlabel metal3 s 31600 200480 32000 200536 6 itasel[650]
port 1547 nsew signal input
rlabel metal3 s 31600 200760 32000 200816 6 itasel[651]
port 1548 nsew signal input
rlabel metal3 s 31600 201040 32000 201096 6 itasel[652]
port 1549 nsew signal input
rlabel metal3 s 31600 201320 32000 201376 6 itasel[653]
port 1550 nsew signal input
rlabel metal3 s 31600 201600 32000 201656 6 itasel[654]
port 1551 nsew signal input
rlabel metal3 s 31600 201880 32000 201936 6 itasel[655]
port 1552 nsew signal input
rlabel metal3 s 31600 202160 32000 202216 6 itasel[656]
port 1553 nsew signal input
rlabel metal3 s 31600 202440 32000 202496 6 itasel[657]
port 1554 nsew signal input
rlabel metal3 s 31600 202720 32000 202776 6 itasel[658]
port 1555 nsew signal input
rlabel metal3 s 31600 203000 32000 203056 6 itasel[659]
port 1556 nsew signal input
rlabel metal3 s 31600 23240 32000 23296 6 itasel[65]
port 1557 nsew signal input
rlabel metal3 s 31600 203280 32000 203336 6 itasel[660]
port 1558 nsew signal input
rlabel metal3 s 31600 203560 32000 203616 6 itasel[661]
port 1559 nsew signal input
rlabel metal3 s 31600 203840 32000 203896 6 itasel[662]
port 1560 nsew signal input
rlabel metal3 s 31600 204120 32000 204176 6 itasel[663]
port 1561 nsew signal input
rlabel metal3 s 31600 204400 32000 204456 6 itasel[664]
port 1562 nsew signal input
rlabel metal3 s 31600 204680 32000 204736 6 itasel[665]
port 1563 nsew signal input
rlabel metal3 s 31600 204960 32000 205016 6 itasel[666]
port 1564 nsew signal input
rlabel metal3 s 31600 205240 32000 205296 6 itasel[667]
port 1565 nsew signal input
rlabel metal3 s 31600 205520 32000 205576 6 itasel[668]
port 1566 nsew signal input
rlabel metal3 s 31600 205800 32000 205856 6 itasel[669]
port 1567 nsew signal input
rlabel metal3 s 31600 23520 32000 23576 6 itasel[66]
port 1568 nsew signal input
rlabel metal3 s 31600 206080 32000 206136 6 itasel[670]
port 1569 nsew signal input
rlabel metal3 s 31600 206360 32000 206416 6 itasel[671]
port 1570 nsew signal input
rlabel metal3 s 0 222320 400 222376 6 itasel[672]
port 1571 nsew signal input
rlabel metal3 s 0 222600 400 222656 6 itasel[673]
port 1572 nsew signal input
rlabel metal3 s 0 222880 400 222936 6 itasel[674]
port 1573 nsew signal input
rlabel metal3 s 0 223160 400 223216 6 itasel[675]
port 1574 nsew signal input
rlabel metal3 s 0 223440 400 223496 6 itasel[676]
port 1575 nsew signal input
rlabel metal3 s 0 223720 400 223776 6 itasel[677]
port 1576 nsew signal input
rlabel metal3 s 0 224000 400 224056 6 itasel[678]
port 1577 nsew signal input
rlabel metal3 s 0 224280 400 224336 6 itasel[679]
port 1578 nsew signal input
rlabel metal3 s 31600 23800 32000 23856 6 itasel[67]
port 1579 nsew signal input
rlabel metal3 s 0 224560 400 224616 6 itasel[680]
port 1580 nsew signal input
rlabel metal3 s 0 224840 400 224896 6 itasel[681]
port 1581 nsew signal input
rlabel metal3 s 0 225120 400 225176 6 itasel[682]
port 1582 nsew signal input
rlabel metal3 s 0 225400 400 225456 6 itasel[683]
port 1583 nsew signal input
rlabel metal3 s 0 225680 400 225736 6 itasel[684]
port 1584 nsew signal input
rlabel metal3 s 0 225960 400 226016 6 itasel[685]
port 1585 nsew signal input
rlabel metal3 s 0 226240 400 226296 6 itasel[686]
port 1586 nsew signal input
rlabel metal3 s 0 226520 400 226576 6 itasel[687]
port 1587 nsew signal input
rlabel metal3 s 0 226800 400 226856 6 itasel[688]
port 1588 nsew signal input
rlabel metal3 s 0 227080 400 227136 6 itasel[689]
port 1589 nsew signal input
rlabel metal3 s 31600 24080 32000 24136 6 itasel[68]
port 1590 nsew signal input
rlabel metal3 s 0 227360 400 227416 6 itasel[690]
port 1591 nsew signal input
rlabel metal3 s 0 227640 400 227696 6 itasel[691]
port 1592 nsew signal input
rlabel metal3 s 0 227920 400 227976 6 itasel[692]
port 1593 nsew signal input
rlabel metal3 s 0 228200 400 228256 6 itasel[693]
port 1594 nsew signal input
rlabel metal3 s 0 228480 400 228536 6 itasel[694]
port 1595 nsew signal input
rlabel metal3 s 0 228760 400 228816 6 itasel[695]
port 1596 nsew signal input
rlabel metal3 s 0 229040 400 229096 6 itasel[696]
port 1597 nsew signal input
rlabel metal3 s 0 229320 400 229376 6 itasel[697]
port 1598 nsew signal input
rlabel metal3 s 0 229600 400 229656 6 itasel[698]
port 1599 nsew signal input
rlabel metal3 s 0 229880 400 229936 6 itasel[699]
port 1600 nsew signal input
rlabel metal3 s 31600 24360 32000 24416 6 itasel[69]
port 1601 nsew signal input
rlabel metal3 s 0 20160 400 20216 6 itasel[6]
port 1602 nsew signal input
rlabel metal3 s 0 230160 400 230216 6 itasel[700]
port 1603 nsew signal input
rlabel metal3 s 0 230440 400 230496 6 itasel[701]
port 1604 nsew signal input
rlabel metal3 s 0 230720 400 230776 6 itasel[702]
port 1605 nsew signal input
rlabel metal3 s 0 231000 400 231056 6 itasel[703]
port 1606 nsew signal input
rlabel metal3 s 0 231280 400 231336 6 itasel[704]
port 1607 nsew signal input
rlabel metal3 s 0 231560 400 231616 6 itasel[705]
port 1608 nsew signal input
rlabel metal3 s 0 231840 400 231896 6 itasel[706]
port 1609 nsew signal input
rlabel metal3 s 0 232120 400 232176 6 itasel[707]
port 1610 nsew signal input
rlabel metal3 s 0 232400 400 232456 6 itasel[708]
port 1611 nsew signal input
rlabel metal3 s 0 232680 400 232736 6 itasel[709]
port 1612 nsew signal input
rlabel metal3 s 31600 24640 32000 24696 6 itasel[70]
port 1613 nsew signal input
rlabel metal3 s 0 232960 400 233016 6 itasel[710]
port 1614 nsew signal input
rlabel metal3 s 0 233240 400 233296 6 itasel[711]
port 1615 nsew signal input
rlabel metal3 s 0 233520 400 233576 6 itasel[712]
port 1616 nsew signal input
rlabel metal3 s 0 233800 400 233856 6 itasel[713]
port 1617 nsew signal input
rlabel metal3 s 0 234080 400 234136 6 itasel[714]
port 1618 nsew signal input
rlabel metal3 s 0 234360 400 234416 6 itasel[715]
port 1619 nsew signal input
rlabel metal3 s 0 234640 400 234696 6 itasel[716]
port 1620 nsew signal input
rlabel metal3 s 0 234920 400 234976 6 itasel[717]
port 1621 nsew signal input
rlabel metal3 s 0 235200 400 235256 6 itasel[718]
port 1622 nsew signal input
rlabel metal3 s 0 235480 400 235536 6 itasel[719]
port 1623 nsew signal input
rlabel metal3 s 31600 24920 32000 24976 6 itasel[71]
port 1624 nsew signal input
rlabel metal3 s 31600 222320 32000 222376 6 itasel[720]
port 1625 nsew signal input
rlabel metal3 s 31600 222600 32000 222656 6 itasel[721]
port 1626 nsew signal input
rlabel metal3 s 31600 222880 32000 222936 6 itasel[722]
port 1627 nsew signal input
rlabel metal3 s 31600 223160 32000 223216 6 itasel[723]
port 1628 nsew signal input
rlabel metal3 s 31600 223440 32000 223496 6 itasel[724]
port 1629 nsew signal input
rlabel metal3 s 31600 223720 32000 223776 6 itasel[725]
port 1630 nsew signal input
rlabel metal3 s 31600 224000 32000 224056 6 itasel[726]
port 1631 nsew signal input
rlabel metal3 s 31600 224280 32000 224336 6 itasel[727]
port 1632 nsew signal input
rlabel metal3 s 31600 224560 32000 224616 6 itasel[728]
port 1633 nsew signal input
rlabel metal3 s 31600 224840 32000 224896 6 itasel[729]
port 1634 nsew signal input
rlabel metal3 s 31600 25200 32000 25256 6 itasel[72]
port 1635 nsew signal input
rlabel metal3 s 31600 225120 32000 225176 6 itasel[730]
port 1636 nsew signal input
rlabel metal3 s 31600 225400 32000 225456 6 itasel[731]
port 1637 nsew signal input
rlabel metal3 s 31600 225680 32000 225736 6 itasel[732]
port 1638 nsew signal input
rlabel metal3 s 31600 225960 32000 226016 6 itasel[733]
port 1639 nsew signal input
rlabel metal3 s 31600 226240 32000 226296 6 itasel[734]
port 1640 nsew signal input
rlabel metal3 s 31600 226520 32000 226576 6 itasel[735]
port 1641 nsew signal input
rlabel metal3 s 31600 226800 32000 226856 6 itasel[736]
port 1642 nsew signal input
rlabel metal3 s 31600 227080 32000 227136 6 itasel[737]
port 1643 nsew signal input
rlabel metal3 s 31600 227360 32000 227416 6 itasel[738]
port 1644 nsew signal input
rlabel metal3 s 31600 227640 32000 227696 6 itasel[739]
port 1645 nsew signal input
rlabel metal3 s 31600 25480 32000 25536 6 itasel[73]
port 1646 nsew signal input
rlabel metal3 s 31600 227920 32000 227976 6 itasel[740]
port 1647 nsew signal input
rlabel metal3 s 31600 228200 32000 228256 6 itasel[741]
port 1648 nsew signal input
rlabel metal3 s 31600 228480 32000 228536 6 itasel[742]
port 1649 nsew signal input
rlabel metal3 s 31600 228760 32000 228816 6 itasel[743]
port 1650 nsew signal input
rlabel metal3 s 31600 229040 32000 229096 6 itasel[744]
port 1651 nsew signal input
rlabel metal3 s 31600 229320 32000 229376 6 itasel[745]
port 1652 nsew signal input
rlabel metal3 s 31600 229600 32000 229656 6 itasel[746]
port 1653 nsew signal input
rlabel metal3 s 31600 229880 32000 229936 6 itasel[747]
port 1654 nsew signal input
rlabel metal3 s 31600 230160 32000 230216 6 itasel[748]
port 1655 nsew signal input
rlabel metal3 s 31600 230440 32000 230496 6 itasel[749]
port 1656 nsew signal input
rlabel metal3 s 31600 25760 32000 25816 6 itasel[74]
port 1657 nsew signal input
rlabel metal3 s 31600 230720 32000 230776 6 itasel[750]
port 1658 nsew signal input
rlabel metal3 s 31600 231000 32000 231056 6 itasel[751]
port 1659 nsew signal input
rlabel metal3 s 31600 231280 32000 231336 6 itasel[752]
port 1660 nsew signal input
rlabel metal3 s 31600 231560 32000 231616 6 itasel[753]
port 1661 nsew signal input
rlabel metal3 s 31600 231840 32000 231896 6 itasel[754]
port 1662 nsew signal input
rlabel metal3 s 31600 232120 32000 232176 6 itasel[755]
port 1663 nsew signal input
rlabel metal3 s 31600 232400 32000 232456 6 itasel[756]
port 1664 nsew signal input
rlabel metal3 s 31600 232680 32000 232736 6 itasel[757]
port 1665 nsew signal input
rlabel metal3 s 31600 232960 32000 233016 6 itasel[758]
port 1666 nsew signal input
rlabel metal3 s 31600 233240 32000 233296 6 itasel[759]
port 1667 nsew signal input
rlabel metal3 s 31600 26040 32000 26096 6 itasel[75]
port 1668 nsew signal input
rlabel metal3 s 31600 233520 32000 233576 6 itasel[760]
port 1669 nsew signal input
rlabel metal3 s 31600 233800 32000 233856 6 itasel[761]
port 1670 nsew signal input
rlabel metal3 s 31600 234080 32000 234136 6 itasel[762]
port 1671 nsew signal input
rlabel metal3 s 31600 234360 32000 234416 6 itasel[763]
port 1672 nsew signal input
rlabel metal3 s 31600 234640 32000 234696 6 itasel[764]
port 1673 nsew signal input
rlabel metal3 s 31600 234920 32000 234976 6 itasel[765]
port 1674 nsew signal input
rlabel metal3 s 31600 235200 32000 235256 6 itasel[766]
port 1675 nsew signal input
rlabel metal3 s 31600 235480 32000 235536 6 itasel[767]
port 1676 nsew signal input
rlabel metal3 s 31600 26320 32000 26376 6 itasel[76]
port 1677 nsew signal input
rlabel metal3 s 31600 26600 32000 26656 6 itasel[77]
port 1678 nsew signal input
rlabel metal3 s 31600 26880 32000 26936 6 itasel[78]
port 1679 nsew signal input
rlabel metal3 s 31600 27160 32000 27216 6 itasel[79]
port 1680 nsew signal input
rlabel metal3 s 0 20440 400 20496 6 itasel[7]
port 1681 nsew signal input
rlabel metal3 s 31600 27440 32000 27496 6 itasel[80]
port 1682 nsew signal input
rlabel metal3 s 31600 27720 32000 27776 6 itasel[81]
port 1683 nsew signal input
rlabel metal3 s 31600 28000 32000 28056 6 itasel[82]
port 1684 nsew signal input
rlabel metal3 s 31600 28280 32000 28336 6 itasel[83]
port 1685 nsew signal input
rlabel metal3 s 31600 28560 32000 28616 6 itasel[84]
port 1686 nsew signal input
rlabel metal3 s 31600 28840 32000 28896 6 itasel[85]
port 1687 nsew signal input
rlabel metal3 s 31600 29120 32000 29176 6 itasel[86]
port 1688 nsew signal input
rlabel metal3 s 31600 29400 32000 29456 6 itasel[87]
port 1689 nsew signal input
rlabel metal3 s 31600 29680 32000 29736 6 itasel[88]
port 1690 nsew signal input
rlabel metal3 s 31600 29960 32000 30016 6 itasel[89]
port 1691 nsew signal input
rlabel metal3 s 0 20720 400 20776 6 itasel[8]
port 1692 nsew signal input
rlabel metal3 s 31600 30240 32000 30296 6 itasel[90]
port 1693 nsew signal input
rlabel metal3 s 31600 30520 32000 30576 6 itasel[91]
port 1694 nsew signal input
rlabel metal3 s 31600 30800 32000 30856 6 itasel[92]
port 1695 nsew signal input
rlabel metal3 s 31600 31080 32000 31136 6 itasel[93]
port 1696 nsew signal input
rlabel metal3 s 31600 31360 32000 31416 6 itasel[94]
port 1697 nsew signal input
rlabel metal3 s 31600 31640 32000 31696 6 itasel[95]
port 1698 nsew signal input
rlabel metal3 s 0 47600 400 47656 6 itasel[96]
port 1699 nsew signal input
rlabel metal3 s 0 47880 400 47936 6 itasel[97]
port 1700 nsew signal input
rlabel metal3 s 0 48160 400 48216 6 itasel[98]
port 1701 nsew signal input
rlabel metal3 s 0 48440 400 48496 6 itasel[99]
port 1702 nsew signal input
rlabel metal3 s 0 21000 400 21056 6 itasel[9]
port 1703 nsew signal input
rlabel metal2 s 560 269800 616 270200 6 nsel[0]
port 1704 nsew signal input
rlabel metal2 s 1120 269800 1176 270200 6 nsel[1]
port 1705 nsew signal input
rlabel metal2 s 1680 269800 1736 270200 6 nsel[2]
port 1706 nsew signal input
rlabel metal2 s 2240 269800 2296 270200 6 nsel[3]
port 1707 nsew signal input
rlabel metal2 s 2800 269800 2856 270200 6 nsel[4]
port 1708 nsew signal input
rlabel metal2 s 3360 269800 3416 270200 6 nsel[5]
port 1709 nsew signal input
rlabel metal2 s 3136 0 3192 400 6 segm[0]
port 1710 nsew signal output
rlabel metal2 s 24416 0 24472 400 6 segm[10]
port 1711 nsew signal output
rlabel metal2 s 26544 0 26600 400 6 segm[11]
port 1712 nsew signal output
rlabel metal2 s 28672 0 28728 400 6 segm[12]
port 1713 nsew signal output
rlabel metal2 s 30800 0 30856 400 6 segm[13]
port 1714 nsew signal output
rlabel metal2 s 5264 0 5320 400 6 segm[1]
port 1715 nsew signal output
rlabel metal2 s 7392 0 7448 400 6 segm[2]
port 1716 nsew signal output
rlabel metal2 s 9520 0 9576 400 6 segm[3]
port 1717 nsew signal output
rlabel metal2 s 11648 0 11704 400 6 segm[4]
port 1718 nsew signal output
rlabel metal2 s 13776 0 13832 400 6 segm[5]
port 1719 nsew signal output
rlabel metal2 s 15904 0 15960 400 6 segm[6]
port 1720 nsew signal output
rlabel metal2 s 18032 0 18088 400 6 segm[7]
port 1721 nsew signal output
rlabel metal2 s 20160 0 20216 400 6 segm[8]
port 1722 nsew signal output
rlabel metal2 s 22288 0 22344 400 6 segm[9]
port 1723 nsew signal output
rlabel metal2 s 3920 269800 3976 270200 6 sel[0]
port 1724 nsew signal output
rlabel metal2 s 9520 269800 9576 270200 6 sel[10]
port 1725 nsew signal output
rlabel metal2 s 10080 269800 10136 270200 6 sel[11]
port 1726 nsew signal output
rlabel metal2 s 4480 269800 4536 270200 6 sel[1]
port 1727 nsew signal output
rlabel metal2 s 5040 269800 5096 270200 6 sel[2]
port 1728 nsew signal output
rlabel metal2 s 5600 269800 5656 270200 6 sel[3]
port 1729 nsew signal output
rlabel metal2 s 6160 269800 6216 270200 6 sel[4]
port 1730 nsew signal output
rlabel metal2 s 6720 269800 6776 270200 6 sel[5]
port 1731 nsew signal output
rlabel metal2 s 7280 269800 7336 270200 6 sel[6]
port 1732 nsew signal output
rlabel metal2 s 7840 269800 7896 270200 6 sel[7]
port 1733 nsew signal output
rlabel metal2 s 8400 269800 8456 270200 6 sel[8]
port 1734 nsew signal output
rlabel metal2 s 8960 269800 9016 270200 6 sel[9]
port 1735 nsew signal output
rlabel metal4 s 2224 1538 2384 268550 6 vdd
port 1736 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 268550 6 vdd
port 1736 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 268550 6 vss
port 1737 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 268550 6 vss
port 1737 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32000 270200
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11760226
string GDS_FILE /home/urielcho/Proyectos_caravel/ITA23_GFMPW1b/openlane/ita/runs/23_11_11_07_55/results/signoff/ita.magic.gds
string GDS_START 312436
<< end >>

