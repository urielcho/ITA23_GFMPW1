VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ita53
  CLASS BLOCK ;
  FOREIGN ita53 ;
  ORIGIN 0.000 0.000 ;
  SIZE 210.000 BY 210.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.400 4.000 134.960 ;
    END
  END clk
  PIN segm[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END segm[0]
  PIN segm[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 206.000 121.520 210.000 ;
    END
  END segm[10]
  PIN segm[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 206.000 111.440 210.000 ;
    END
  END segm[11]
  PIN segm[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 77.280 210.000 77.840 ;
    END
  END segm[12]
  PIN segm[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.240 4.000 114.800 ;
    END
  END segm[13]
  PIN segm[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 114.240 210.000 114.800 ;
    END
  END segm[1]
  PIN segm[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 206.000 87.920 210.000 ;
    END
  END segm[2]
  PIN segm[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.880 4.000 111.440 ;
    END
  END segm[3]
  PIN segm[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 110.880 210.000 111.440 ;
    END
  END segm[4]
  PIN segm[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 206.000 81.200 210.000 ;
    END
  END segm[5]
  PIN segm[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END segm[6]
  PIN segm[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 206.000 84.560 210.000 ;
    END
  END segm[7]
  PIN segm[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 134.400 210.000 134.960 ;
    END
  END segm[8]
  PIN segm[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 131.040 210.000 131.600 ;
    END
  END segm[9]
  PIN sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 0.000 87.920 4.000 ;
    END
  END sel[0]
  PIN sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.360 4.000 87.920 ;
    END
  END sel[10]
  PIN sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 0.000 128.240 4.000 ;
    END
  END sel[11]
  PIN sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 100.800 210.000 101.360 ;
    END
  END sel[1]
  PIN sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 206.000 91.280 210.000 ;
    END
  END sel[2]
  PIN sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 4.000 ;
    END
  END sel[3]
  PIN sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 0.000 108.080 4.000 ;
    END
  END sel[4]
  PIN sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 206.000 104.720 210.000 ;
    END
  END sel[5]
  PIN sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 117.600 210.000 118.160 ;
    END
  END sel[6]
  PIN sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 84.000 210.000 84.560 ;
    END
  END sel[7]
  PIN sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.800 4.000 101.360 ;
    END
  END sel[8]
  PIN sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 97.440 210.000 98.000 ;
    END
  END sel[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 192.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 192.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 192.380 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 203.280 192.380 ;
      LAYER Metal2 ;
        RECT 9.660 205.700 80.340 206.000 ;
        RECT 81.500 205.700 83.700 206.000 ;
        RECT 84.860 205.700 87.060 206.000 ;
        RECT 88.220 205.700 90.420 206.000 ;
        RECT 91.580 205.700 103.860 206.000 ;
        RECT 105.020 205.700 110.580 206.000 ;
        RECT 111.740 205.700 120.660 206.000 ;
        RECT 121.820 205.700 200.340 206.000 ;
        RECT 9.660 4.300 200.340 205.700 ;
        RECT 9.660 4.000 87.060 4.300 ;
        RECT 88.220 4.000 90.420 4.300 ;
        RECT 91.580 4.000 107.220 4.300 ;
        RECT 108.380 4.000 110.580 4.300 ;
        RECT 111.740 4.000 127.380 4.300 ;
        RECT 128.540 4.000 200.340 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 135.260 206.000 192.220 ;
        RECT 4.300 134.100 205.700 135.260 ;
        RECT 4.000 131.900 206.000 134.100 ;
        RECT 4.000 130.740 205.700 131.900 ;
        RECT 4.000 118.460 206.000 130.740 ;
        RECT 4.300 117.300 205.700 118.460 ;
        RECT 4.000 115.100 206.000 117.300 ;
        RECT 4.300 113.940 205.700 115.100 ;
        RECT 4.000 111.740 206.000 113.940 ;
        RECT 4.300 110.580 205.700 111.740 ;
        RECT 4.000 101.660 206.000 110.580 ;
        RECT 4.300 100.500 205.700 101.660 ;
        RECT 4.000 98.300 206.000 100.500 ;
        RECT 4.000 97.140 205.700 98.300 ;
        RECT 4.000 88.220 206.000 97.140 ;
        RECT 4.300 87.060 206.000 88.220 ;
        RECT 4.000 84.860 206.000 87.060 ;
        RECT 4.000 83.700 205.700 84.860 ;
        RECT 4.000 78.140 206.000 83.700 ;
        RECT 4.000 76.980 205.700 78.140 ;
        RECT 4.000 15.540 206.000 76.980 ;
      LAYER Metal4 ;
        RECT 92.540 106.490 92.820 118.070 ;
  END
END ita53
END LIBRARY

