// This is the unpowered netlist.
module user_project_wrapper (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire \itasegm1[0] ;
 wire \itasegm1[100] ;
 wire \itasegm1[101] ;
 wire \itasegm1[102] ;
 wire \itasegm1[103] ;
 wire \itasegm1[104] ;
 wire \itasegm1[105] ;
 wire \itasegm1[106] ;
 wire \itasegm1[107] ;
 wire \itasegm1[108] ;
 wire \itasegm1[109] ;
 wire \itasegm1[10] ;
 wire \itasegm1[110] ;
 wire \itasegm1[111] ;
 wire \itasegm1[112] ;
 wire \itasegm1[113] ;
 wire \itasegm1[114] ;
 wire \itasegm1[115] ;
 wire \itasegm1[116] ;
 wire \itasegm1[117] ;
 wire \itasegm1[118] ;
 wire \itasegm1[119] ;
 wire \itasegm1[11] ;
 wire \itasegm1[120] ;
 wire \itasegm1[121] ;
 wire \itasegm1[122] ;
 wire \itasegm1[123] ;
 wire \itasegm1[124] ;
 wire \itasegm1[125] ;
 wire \itasegm1[126] ;
 wire \itasegm1[127] ;
 wire \itasegm1[128] ;
 wire \itasegm1[129] ;
 wire \itasegm1[12] ;
 wire \itasegm1[130] ;
 wire \itasegm1[131] ;
 wire \itasegm1[132] ;
 wire \itasegm1[133] ;
 wire \itasegm1[134] ;
 wire \itasegm1[135] ;
 wire \itasegm1[136] ;
 wire \itasegm1[137] ;
 wire \itasegm1[138] ;
 wire \itasegm1[139] ;
 wire \itasegm1[13] ;
 wire \itasegm1[140] ;
 wire \itasegm1[141] ;
 wire \itasegm1[142] ;
 wire \itasegm1[143] ;
 wire \itasegm1[144] ;
 wire \itasegm1[145] ;
 wire \itasegm1[146] ;
 wire \itasegm1[147] ;
 wire \itasegm1[148] ;
 wire \itasegm1[149] ;
 wire \itasegm1[14] ;
 wire \itasegm1[150] ;
 wire \itasegm1[151] ;
 wire \itasegm1[152] ;
 wire \itasegm1[153] ;
 wire \itasegm1[154] ;
 wire \itasegm1[155] ;
 wire \itasegm1[156] ;
 wire \itasegm1[157] ;
 wire \itasegm1[158] ;
 wire \itasegm1[159] ;
 wire \itasegm1[15] ;
 wire \itasegm1[160] ;
 wire \itasegm1[161] ;
 wire \itasegm1[162] ;
 wire \itasegm1[163] ;
 wire \itasegm1[164] ;
 wire \itasegm1[165] ;
 wire \itasegm1[166] ;
 wire \itasegm1[167] ;
 wire \itasegm1[168] ;
 wire \itasegm1[169] ;
 wire \itasegm1[16] ;
 wire \itasegm1[170] ;
 wire \itasegm1[171] ;
 wire \itasegm1[172] ;
 wire \itasegm1[173] ;
 wire \itasegm1[174] ;
 wire \itasegm1[175] ;
 wire \itasegm1[176] ;
 wire \itasegm1[177] ;
 wire \itasegm1[178] ;
 wire \itasegm1[179] ;
 wire \itasegm1[17] ;
 wire \itasegm1[180] ;
 wire \itasegm1[181] ;
 wire \itasegm1[182] ;
 wire \itasegm1[183] ;
 wire \itasegm1[184] ;
 wire \itasegm1[185] ;
 wire \itasegm1[186] ;
 wire \itasegm1[187] ;
 wire \itasegm1[188] ;
 wire \itasegm1[189] ;
 wire \itasegm1[18] ;
 wire \itasegm1[190] ;
 wire \itasegm1[191] ;
 wire \itasegm1[192] ;
 wire \itasegm1[193] ;
 wire \itasegm1[194] ;
 wire \itasegm1[195] ;
 wire \itasegm1[196] ;
 wire \itasegm1[197] ;
 wire \itasegm1[198] ;
 wire \itasegm1[199] ;
 wire \itasegm1[19] ;
 wire \itasegm1[1] ;
 wire \itasegm1[200] ;
 wire \itasegm1[201] ;
 wire \itasegm1[202] ;
 wire \itasegm1[203] ;
 wire \itasegm1[204] ;
 wire \itasegm1[205] ;
 wire \itasegm1[206] ;
 wire \itasegm1[207] ;
 wire \itasegm1[208] ;
 wire \itasegm1[209] ;
 wire \itasegm1[20] ;
 wire \itasegm1[210] ;
 wire \itasegm1[211] ;
 wire \itasegm1[212] ;
 wire \itasegm1[213] ;
 wire \itasegm1[214] ;
 wire \itasegm1[215] ;
 wire \itasegm1[216] ;
 wire \itasegm1[217] ;
 wire \itasegm1[218] ;
 wire \itasegm1[219] ;
 wire \itasegm1[21] ;
 wire \itasegm1[220] ;
 wire \itasegm1[221] ;
 wire \itasegm1[222] ;
 wire \itasegm1[223] ;
 wire \itasegm1[224] ;
 wire \itasegm1[225] ;
 wire \itasegm1[226] ;
 wire \itasegm1[227] ;
 wire \itasegm1[228] ;
 wire \itasegm1[229] ;
 wire \itasegm1[22] ;
 wire \itasegm1[230] ;
 wire \itasegm1[231] ;
 wire \itasegm1[232] ;
 wire \itasegm1[233] ;
 wire \itasegm1[234] ;
 wire \itasegm1[235] ;
 wire \itasegm1[236] ;
 wire \itasegm1[237] ;
 wire \itasegm1[238] ;
 wire \itasegm1[239] ;
 wire \itasegm1[23] ;
 wire \itasegm1[240] ;
 wire \itasegm1[241] ;
 wire \itasegm1[242] ;
 wire \itasegm1[243] ;
 wire \itasegm1[244] ;
 wire \itasegm1[245] ;
 wire \itasegm1[246] ;
 wire \itasegm1[247] ;
 wire \itasegm1[248] ;
 wire \itasegm1[249] ;
 wire \itasegm1[24] ;
 wire \itasegm1[250] ;
 wire \itasegm1[251] ;
 wire \itasegm1[252] ;
 wire \itasegm1[253] ;
 wire \itasegm1[254] ;
 wire \itasegm1[255] ;
 wire \itasegm1[256] ;
 wire \itasegm1[257] ;
 wire \itasegm1[258] ;
 wire \itasegm1[259] ;
 wire \itasegm1[25] ;
 wire \itasegm1[260] ;
 wire \itasegm1[261] ;
 wire \itasegm1[262] ;
 wire \itasegm1[263] ;
 wire \itasegm1[264] ;
 wire \itasegm1[265] ;
 wire \itasegm1[266] ;
 wire \itasegm1[267] ;
 wire \itasegm1[268] ;
 wire \itasegm1[269] ;
 wire \itasegm1[26] ;
 wire \itasegm1[270] ;
 wire \itasegm1[271] ;
 wire \itasegm1[272] ;
 wire \itasegm1[273] ;
 wire \itasegm1[274] ;
 wire \itasegm1[275] ;
 wire \itasegm1[276] ;
 wire \itasegm1[277] ;
 wire \itasegm1[278] ;
 wire \itasegm1[279] ;
 wire \itasegm1[27] ;
 wire \itasegm1[280] ;
 wire \itasegm1[281] ;
 wire \itasegm1[282] ;
 wire \itasegm1[283] ;
 wire \itasegm1[284] ;
 wire \itasegm1[285] ;
 wire \itasegm1[286] ;
 wire \itasegm1[287] ;
 wire \itasegm1[288] ;
 wire \itasegm1[289] ;
 wire \itasegm1[28] ;
 wire \itasegm1[290] ;
 wire \itasegm1[291] ;
 wire \itasegm1[292] ;
 wire \itasegm1[293] ;
 wire \itasegm1[294] ;
 wire \itasegm1[295] ;
 wire \itasegm1[296] ;
 wire \itasegm1[297] ;
 wire \itasegm1[298] ;
 wire \itasegm1[299] ;
 wire \itasegm1[29] ;
 wire \itasegm1[2] ;
 wire \itasegm1[300] ;
 wire \itasegm1[301] ;
 wire \itasegm1[302] ;
 wire \itasegm1[303] ;
 wire \itasegm1[304] ;
 wire \itasegm1[305] ;
 wire \itasegm1[306] ;
 wire \itasegm1[307] ;
 wire \itasegm1[308] ;
 wire \itasegm1[309] ;
 wire \itasegm1[30] ;
 wire \itasegm1[310] ;
 wire \itasegm1[311] ;
 wire \itasegm1[312] ;
 wire \itasegm1[313] ;
 wire \itasegm1[314] ;
 wire \itasegm1[315] ;
 wire \itasegm1[316] ;
 wire \itasegm1[317] ;
 wire \itasegm1[318] ;
 wire \itasegm1[319] ;
 wire \itasegm1[31] ;
 wire \itasegm1[320] ;
 wire \itasegm1[321] ;
 wire \itasegm1[322] ;
 wire \itasegm1[323] ;
 wire \itasegm1[324] ;
 wire \itasegm1[325] ;
 wire \itasegm1[326] ;
 wire \itasegm1[327] ;
 wire \itasegm1[328] ;
 wire \itasegm1[329] ;
 wire \itasegm1[32] ;
 wire \itasegm1[330] ;
 wire \itasegm1[331] ;
 wire \itasegm1[332] ;
 wire \itasegm1[333] ;
 wire \itasegm1[334] ;
 wire \itasegm1[335] ;
 wire \itasegm1[336] ;
 wire \itasegm1[337] ;
 wire \itasegm1[338] ;
 wire \itasegm1[339] ;
 wire \itasegm1[33] ;
 wire \itasegm1[340] ;
 wire \itasegm1[341] ;
 wire \itasegm1[342] ;
 wire \itasegm1[343] ;
 wire \itasegm1[344] ;
 wire \itasegm1[345] ;
 wire \itasegm1[346] ;
 wire \itasegm1[347] ;
 wire \itasegm1[348] ;
 wire \itasegm1[349] ;
 wire \itasegm1[34] ;
 wire \itasegm1[350] ;
 wire \itasegm1[351] ;
 wire \itasegm1[352] ;
 wire \itasegm1[353] ;
 wire \itasegm1[354] ;
 wire \itasegm1[355] ;
 wire \itasegm1[356] ;
 wire \itasegm1[357] ;
 wire \itasegm1[358] ;
 wire \itasegm1[359] ;
 wire \itasegm1[35] ;
 wire \itasegm1[360] ;
 wire \itasegm1[361] ;
 wire \itasegm1[362] ;
 wire \itasegm1[363] ;
 wire \itasegm1[364] ;
 wire \itasegm1[365] ;
 wire \itasegm1[366] ;
 wire \itasegm1[367] ;
 wire \itasegm1[368] ;
 wire \itasegm1[369] ;
 wire \itasegm1[36] ;
 wire \itasegm1[370] ;
 wire \itasegm1[371] ;
 wire \itasegm1[372] ;
 wire \itasegm1[373] ;
 wire \itasegm1[374] ;
 wire \itasegm1[375] ;
 wire \itasegm1[376] ;
 wire \itasegm1[377] ;
 wire \itasegm1[378] ;
 wire \itasegm1[379] ;
 wire \itasegm1[37] ;
 wire \itasegm1[380] ;
 wire \itasegm1[381] ;
 wire \itasegm1[382] ;
 wire \itasegm1[383] ;
 wire \itasegm1[384] ;
 wire \itasegm1[385] ;
 wire \itasegm1[386] ;
 wire \itasegm1[387] ;
 wire \itasegm1[388] ;
 wire \itasegm1[389] ;
 wire \itasegm1[38] ;
 wire \itasegm1[390] ;
 wire \itasegm1[391] ;
 wire \itasegm1[392] ;
 wire \itasegm1[393] ;
 wire \itasegm1[394] ;
 wire \itasegm1[395] ;
 wire \itasegm1[396] ;
 wire \itasegm1[397] ;
 wire \itasegm1[398] ;
 wire \itasegm1[399] ;
 wire \itasegm1[39] ;
 wire \itasegm1[3] ;
 wire \itasegm1[400] ;
 wire \itasegm1[401] ;
 wire \itasegm1[402] ;
 wire \itasegm1[403] ;
 wire \itasegm1[404] ;
 wire \itasegm1[405] ;
 wire \itasegm1[406] ;
 wire \itasegm1[407] ;
 wire \itasegm1[408] ;
 wire \itasegm1[409] ;
 wire \itasegm1[40] ;
 wire \itasegm1[410] ;
 wire \itasegm1[411] ;
 wire \itasegm1[412] ;
 wire \itasegm1[413] ;
 wire \itasegm1[414] ;
 wire \itasegm1[415] ;
 wire \itasegm1[416] ;
 wire \itasegm1[417] ;
 wire \itasegm1[418] ;
 wire \itasegm1[419] ;
 wire \itasegm1[41] ;
 wire \itasegm1[420] ;
 wire \itasegm1[421] ;
 wire \itasegm1[422] ;
 wire \itasegm1[423] ;
 wire \itasegm1[424] ;
 wire \itasegm1[425] ;
 wire \itasegm1[426] ;
 wire \itasegm1[427] ;
 wire \itasegm1[428] ;
 wire \itasegm1[429] ;
 wire \itasegm1[42] ;
 wire \itasegm1[430] ;
 wire \itasegm1[431] ;
 wire \itasegm1[432] ;
 wire \itasegm1[433] ;
 wire \itasegm1[434] ;
 wire \itasegm1[435] ;
 wire \itasegm1[436] ;
 wire \itasegm1[437] ;
 wire \itasegm1[438] ;
 wire \itasegm1[439] ;
 wire \itasegm1[43] ;
 wire \itasegm1[440] ;
 wire \itasegm1[441] ;
 wire \itasegm1[442] ;
 wire \itasegm1[443] ;
 wire \itasegm1[444] ;
 wire \itasegm1[445] ;
 wire \itasegm1[446] ;
 wire \itasegm1[447] ;
 wire \itasegm1[448] ;
 wire \itasegm1[449] ;
 wire \itasegm1[44] ;
 wire \itasegm1[450] ;
 wire \itasegm1[451] ;
 wire \itasegm1[452] ;
 wire \itasegm1[453] ;
 wire \itasegm1[454] ;
 wire \itasegm1[455] ;
 wire \itasegm1[456] ;
 wire \itasegm1[457] ;
 wire \itasegm1[458] ;
 wire \itasegm1[459] ;
 wire \itasegm1[45] ;
 wire \itasegm1[460] ;
 wire \itasegm1[461] ;
 wire \itasegm1[462] ;
 wire \itasegm1[463] ;
 wire \itasegm1[464] ;
 wire \itasegm1[465] ;
 wire \itasegm1[466] ;
 wire \itasegm1[467] ;
 wire \itasegm1[468] ;
 wire \itasegm1[469] ;
 wire \itasegm1[46] ;
 wire \itasegm1[470] ;
 wire \itasegm1[471] ;
 wire \itasegm1[472] ;
 wire \itasegm1[473] ;
 wire \itasegm1[474] ;
 wire \itasegm1[475] ;
 wire \itasegm1[476] ;
 wire \itasegm1[477] ;
 wire \itasegm1[478] ;
 wire \itasegm1[479] ;
 wire \itasegm1[47] ;
 wire \itasegm1[480] ;
 wire \itasegm1[481] ;
 wire \itasegm1[482] ;
 wire \itasegm1[483] ;
 wire \itasegm1[484] ;
 wire \itasegm1[485] ;
 wire \itasegm1[486] ;
 wire \itasegm1[487] ;
 wire \itasegm1[488] ;
 wire \itasegm1[489] ;
 wire \itasegm1[48] ;
 wire \itasegm1[490] ;
 wire \itasegm1[491] ;
 wire \itasegm1[492] ;
 wire \itasegm1[493] ;
 wire \itasegm1[494] ;
 wire \itasegm1[495] ;
 wire \itasegm1[496] ;
 wire \itasegm1[497] ;
 wire \itasegm1[498] ;
 wire \itasegm1[499] ;
 wire \itasegm1[49] ;
 wire \itasegm1[4] ;
 wire \itasegm1[500] ;
 wire \itasegm1[501] ;
 wire \itasegm1[502] ;
 wire \itasegm1[503] ;
 wire \itasegm1[504] ;
 wire \itasegm1[505] ;
 wire \itasegm1[506] ;
 wire \itasegm1[507] ;
 wire \itasegm1[508] ;
 wire \itasegm1[509] ;
 wire \itasegm1[50] ;
 wire \itasegm1[510] ;
 wire \itasegm1[511] ;
 wire \itasegm1[512] ;
 wire \itasegm1[513] ;
 wire \itasegm1[514] ;
 wire \itasegm1[515] ;
 wire \itasegm1[516] ;
 wire \itasegm1[517] ;
 wire \itasegm1[518] ;
 wire \itasegm1[519] ;
 wire \itasegm1[51] ;
 wire \itasegm1[520] ;
 wire \itasegm1[521] ;
 wire \itasegm1[522] ;
 wire \itasegm1[523] ;
 wire \itasegm1[524] ;
 wire \itasegm1[525] ;
 wire \itasegm1[526] ;
 wire \itasegm1[527] ;
 wire \itasegm1[528] ;
 wire \itasegm1[529] ;
 wire \itasegm1[52] ;
 wire \itasegm1[530] ;
 wire \itasegm1[531] ;
 wire \itasegm1[532] ;
 wire \itasegm1[533] ;
 wire \itasegm1[534] ;
 wire \itasegm1[535] ;
 wire \itasegm1[536] ;
 wire \itasegm1[537] ;
 wire \itasegm1[538] ;
 wire \itasegm1[539] ;
 wire \itasegm1[53] ;
 wire \itasegm1[540] ;
 wire \itasegm1[541] ;
 wire \itasegm1[542] ;
 wire \itasegm1[543] ;
 wire \itasegm1[544] ;
 wire \itasegm1[545] ;
 wire \itasegm1[546] ;
 wire \itasegm1[547] ;
 wire \itasegm1[548] ;
 wire \itasegm1[549] ;
 wire \itasegm1[54] ;
 wire \itasegm1[550] ;
 wire \itasegm1[551] ;
 wire \itasegm1[552] ;
 wire \itasegm1[553] ;
 wire \itasegm1[554] ;
 wire \itasegm1[555] ;
 wire \itasegm1[556] ;
 wire \itasegm1[557] ;
 wire \itasegm1[558] ;
 wire \itasegm1[559] ;
 wire \itasegm1[55] ;
 wire \itasegm1[560] ;
 wire \itasegm1[561] ;
 wire \itasegm1[562] ;
 wire \itasegm1[563] ;
 wire \itasegm1[564] ;
 wire \itasegm1[565] ;
 wire \itasegm1[566] ;
 wire \itasegm1[567] ;
 wire \itasegm1[568] ;
 wire \itasegm1[569] ;
 wire \itasegm1[56] ;
 wire \itasegm1[570] ;
 wire \itasegm1[571] ;
 wire \itasegm1[572] ;
 wire \itasegm1[573] ;
 wire \itasegm1[574] ;
 wire \itasegm1[575] ;
 wire \itasegm1[576] ;
 wire \itasegm1[577] ;
 wire \itasegm1[578] ;
 wire \itasegm1[579] ;
 wire \itasegm1[57] ;
 wire \itasegm1[580] ;
 wire \itasegm1[581] ;
 wire \itasegm1[582] ;
 wire \itasegm1[583] ;
 wire \itasegm1[584] ;
 wire \itasegm1[585] ;
 wire \itasegm1[586] ;
 wire \itasegm1[587] ;
 wire \itasegm1[588] ;
 wire \itasegm1[589] ;
 wire \itasegm1[58] ;
 wire \itasegm1[590] ;
 wire \itasegm1[591] ;
 wire \itasegm1[592] ;
 wire \itasegm1[593] ;
 wire \itasegm1[594] ;
 wire \itasegm1[595] ;
 wire \itasegm1[596] ;
 wire \itasegm1[597] ;
 wire \itasegm1[598] ;
 wire \itasegm1[599] ;
 wire \itasegm1[59] ;
 wire \itasegm1[5] ;
 wire \itasegm1[600] ;
 wire \itasegm1[601] ;
 wire \itasegm1[602] ;
 wire \itasegm1[603] ;
 wire \itasegm1[604] ;
 wire \itasegm1[605] ;
 wire \itasegm1[606] ;
 wire \itasegm1[607] ;
 wire \itasegm1[608] ;
 wire \itasegm1[609] ;
 wire \itasegm1[60] ;
 wire \itasegm1[610] ;
 wire \itasegm1[611] ;
 wire \itasegm1[612] ;
 wire \itasegm1[613] ;
 wire \itasegm1[614] ;
 wire \itasegm1[615] ;
 wire \itasegm1[616] ;
 wire \itasegm1[617] ;
 wire \itasegm1[618] ;
 wire \itasegm1[619] ;
 wire \itasegm1[61] ;
 wire \itasegm1[620] ;
 wire \itasegm1[621] ;
 wire \itasegm1[622] ;
 wire \itasegm1[623] ;
 wire \itasegm1[624] ;
 wire \itasegm1[625] ;
 wire \itasegm1[626] ;
 wire \itasegm1[627] ;
 wire \itasegm1[628] ;
 wire \itasegm1[629] ;
 wire \itasegm1[62] ;
 wire \itasegm1[630] ;
 wire \itasegm1[631] ;
 wire \itasegm1[632] ;
 wire \itasegm1[633] ;
 wire \itasegm1[634] ;
 wire \itasegm1[635] ;
 wire \itasegm1[636] ;
 wire \itasegm1[637] ;
 wire \itasegm1[638] ;
 wire \itasegm1[639] ;
 wire \itasegm1[63] ;
 wire \itasegm1[640] ;
 wire \itasegm1[641] ;
 wire \itasegm1[642] ;
 wire \itasegm1[643] ;
 wire \itasegm1[644] ;
 wire \itasegm1[645] ;
 wire \itasegm1[646] ;
 wire \itasegm1[647] ;
 wire \itasegm1[648] ;
 wire \itasegm1[649] ;
 wire \itasegm1[64] ;
 wire \itasegm1[650] ;
 wire \itasegm1[651] ;
 wire \itasegm1[652] ;
 wire \itasegm1[653] ;
 wire \itasegm1[654] ;
 wire \itasegm1[655] ;
 wire \itasegm1[656] ;
 wire \itasegm1[657] ;
 wire \itasegm1[658] ;
 wire \itasegm1[659] ;
 wire \itasegm1[65] ;
 wire \itasegm1[660] ;
 wire \itasegm1[661] ;
 wire \itasegm1[662] ;
 wire \itasegm1[663] ;
 wire \itasegm1[664] ;
 wire \itasegm1[665] ;
 wire \itasegm1[666] ;
 wire \itasegm1[667] ;
 wire \itasegm1[668] ;
 wire \itasegm1[669] ;
 wire \itasegm1[66] ;
 wire \itasegm1[670] ;
 wire \itasegm1[671] ;
 wire \itasegm1[672] ;
 wire \itasegm1[673] ;
 wire \itasegm1[674] ;
 wire \itasegm1[675] ;
 wire \itasegm1[676] ;
 wire \itasegm1[677] ;
 wire \itasegm1[678] ;
 wire \itasegm1[679] ;
 wire \itasegm1[67] ;
 wire \itasegm1[680] ;
 wire \itasegm1[681] ;
 wire \itasegm1[682] ;
 wire \itasegm1[683] ;
 wire \itasegm1[684] ;
 wire \itasegm1[685] ;
 wire \itasegm1[686] ;
 wire \itasegm1[687] ;
 wire \itasegm1[688] ;
 wire \itasegm1[689] ;
 wire \itasegm1[68] ;
 wire \itasegm1[690] ;
 wire \itasegm1[691] ;
 wire \itasegm1[692] ;
 wire \itasegm1[693] ;
 wire \itasegm1[694] ;
 wire \itasegm1[695] ;
 wire \itasegm1[696] ;
 wire \itasegm1[697] ;
 wire \itasegm1[698] ;
 wire \itasegm1[699] ;
 wire \itasegm1[69] ;
 wire \itasegm1[6] ;
 wire \itasegm1[700] ;
 wire \itasegm1[701] ;
 wire \itasegm1[702] ;
 wire \itasegm1[703] ;
 wire \itasegm1[704] ;
 wire \itasegm1[705] ;
 wire \itasegm1[706] ;
 wire \itasegm1[707] ;
 wire \itasegm1[708] ;
 wire \itasegm1[709] ;
 wire \itasegm1[70] ;
 wire \itasegm1[710] ;
 wire \itasegm1[711] ;
 wire \itasegm1[712] ;
 wire \itasegm1[713] ;
 wire \itasegm1[714] ;
 wire \itasegm1[715] ;
 wire \itasegm1[716] ;
 wire \itasegm1[717] ;
 wire \itasegm1[718] ;
 wire \itasegm1[719] ;
 wire \itasegm1[71] ;
 wire \itasegm1[720] ;
 wire \itasegm1[721] ;
 wire \itasegm1[722] ;
 wire \itasegm1[723] ;
 wire \itasegm1[724] ;
 wire \itasegm1[725] ;
 wire \itasegm1[726] ;
 wire \itasegm1[727] ;
 wire \itasegm1[728] ;
 wire \itasegm1[729] ;
 wire \itasegm1[72] ;
 wire \itasegm1[730] ;
 wire \itasegm1[731] ;
 wire \itasegm1[732] ;
 wire \itasegm1[733] ;
 wire \itasegm1[734] ;
 wire \itasegm1[735] ;
 wire \itasegm1[736] ;
 wire \itasegm1[737] ;
 wire \itasegm1[738] ;
 wire \itasegm1[739] ;
 wire \itasegm1[73] ;
 wire \itasegm1[740] ;
 wire \itasegm1[741] ;
 wire \itasegm1[742] ;
 wire \itasegm1[743] ;
 wire \itasegm1[744] ;
 wire \itasegm1[745] ;
 wire \itasegm1[746] ;
 wire \itasegm1[747] ;
 wire \itasegm1[748] ;
 wire \itasegm1[749] ;
 wire \itasegm1[74] ;
 wire \itasegm1[750] ;
 wire \itasegm1[751] ;
 wire \itasegm1[752] ;
 wire \itasegm1[753] ;
 wire \itasegm1[754] ;
 wire \itasegm1[755] ;
 wire \itasegm1[756] ;
 wire \itasegm1[757] ;
 wire \itasegm1[758] ;
 wire \itasegm1[759] ;
 wire \itasegm1[75] ;
 wire \itasegm1[760] ;
 wire \itasegm1[761] ;
 wire \itasegm1[762] ;
 wire \itasegm1[763] ;
 wire \itasegm1[764] ;
 wire \itasegm1[765] ;
 wire \itasegm1[766] ;
 wire \itasegm1[767] ;
 wire \itasegm1[768] ;
 wire \itasegm1[769] ;
 wire \itasegm1[76] ;
 wire \itasegm1[770] ;
 wire \itasegm1[771] ;
 wire \itasegm1[772] ;
 wire \itasegm1[773] ;
 wire \itasegm1[774] ;
 wire \itasegm1[775] ;
 wire \itasegm1[776] ;
 wire \itasegm1[777] ;
 wire \itasegm1[778] ;
 wire \itasegm1[779] ;
 wire \itasegm1[77] ;
 wire \itasegm1[780] ;
 wire \itasegm1[781] ;
 wire \itasegm1[782] ;
 wire \itasegm1[783] ;
 wire \itasegm1[784] ;
 wire \itasegm1[785] ;
 wire \itasegm1[786] ;
 wire \itasegm1[787] ;
 wire \itasegm1[788] ;
 wire \itasegm1[789] ;
 wire \itasegm1[78] ;
 wire \itasegm1[790] ;
 wire \itasegm1[791] ;
 wire \itasegm1[792] ;
 wire \itasegm1[793] ;
 wire \itasegm1[794] ;
 wire \itasegm1[795] ;
 wire \itasegm1[796] ;
 wire \itasegm1[797] ;
 wire \itasegm1[798] ;
 wire \itasegm1[799] ;
 wire \itasegm1[79] ;
 wire \itasegm1[7] ;
 wire \itasegm1[800] ;
 wire \itasegm1[801] ;
 wire \itasegm1[802] ;
 wire \itasegm1[803] ;
 wire \itasegm1[804] ;
 wire \itasegm1[805] ;
 wire \itasegm1[806] ;
 wire \itasegm1[807] ;
 wire \itasegm1[808] ;
 wire \itasegm1[809] ;
 wire \itasegm1[80] ;
 wire \itasegm1[810] ;
 wire \itasegm1[811] ;
 wire \itasegm1[812] ;
 wire \itasegm1[813] ;
 wire \itasegm1[814] ;
 wire \itasegm1[815] ;
 wire \itasegm1[816] ;
 wire \itasegm1[817] ;
 wire \itasegm1[818] ;
 wire \itasegm1[819] ;
 wire \itasegm1[81] ;
 wire \itasegm1[820] ;
 wire \itasegm1[821] ;
 wire \itasegm1[822] ;
 wire \itasegm1[823] ;
 wire \itasegm1[824] ;
 wire \itasegm1[825] ;
 wire \itasegm1[826] ;
 wire \itasegm1[827] ;
 wire \itasegm1[828] ;
 wire \itasegm1[829] ;
 wire \itasegm1[82] ;
 wire \itasegm1[830] ;
 wire \itasegm1[831] ;
 wire \itasegm1[832] ;
 wire \itasegm1[833] ;
 wire \itasegm1[834] ;
 wire \itasegm1[835] ;
 wire \itasegm1[836] ;
 wire \itasegm1[837] ;
 wire \itasegm1[838] ;
 wire \itasegm1[839] ;
 wire \itasegm1[83] ;
 wire \itasegm1[840] ;
 wire \itasegm1[841] ;
 wire \itasegm1[842] ;
 wire \itasegm1[843] ;
 wire \itasegm1[844] ;
 wire \itasegm1[845] ;
 wire \itasegm1[846] ;
 wire \itasegm1[847] ;
 wire \itasegm1[848] ;
 wire \itasegm1[849] ;
 wire \itasegm1[84] ;
 wire \itasegm1[850] ;
 wire \itasegm1[851] ;
 wire \itasegm1[852] ;
 wire \itasegm1[853] ;
 wire \itasegm1[854] ;
 wire \itasegm1[855] ;
 wire \itasegm1[856] ;
 wire \itasegm1[857] ;
 wire \itasegm1[858] ;
 wire \itasegm1[859] ;
 wire \itasegm1[85] ;
 wire \itasegm1[860] ;
 wire \itasegm1[861] ;
 wire \itasegm1[862] ;
 wire \itasegm1[863] ;
 wire \itasegm1[864] ;
 wire \itasegm1[865] ;
 wire \itasegm1[866] ;
 wire \itasegm1[867] ;
 wire \itasegm1[868] ;
 wire \itasegm1[869] ;
 wire \itasegm1[86] ;
 wire \itasegm1[870] ;
 wire \itasegm1[871] ;
 wire \itasegm1[872] ;
 wire \itasegm1[873] ;
 wire \itasegm1[874] ;
 wire \itasegm1[875] ;
 wire \itasegm1[876] ;
 wire \itasegm1[877] ;
 wire \itasegm1[878] ;
 wire \itasegm1[879] ;
 wire \itasegm1[87] ;
 wire \itasegm1[880] ;
 wire \itasegm1[881] ;
 wire \itasegm1[882] ;
 wire \itasegm1[883] ;
 wire \itasegm1[884] ;
 wire \itasegm1[885] ;
 wire \itasegm1[886] ;
 wire \itasegm1[887] ;
 wire \itasegm1[888] ;
 wire \itasegm1[889] ;
 wire \itasegm1[88] ;
 wire \itasegm1[890] ;
 wire \itasegm1[891] ;
 wire \itasegm1[892] ;
 wire \itasegm1[893] ;
 wire \itasegm1[894] ;
 wire \itasegm1[895] ;
 wire \itasegm1[89] ;
 wire \itasegm1[8] ;
 wire \itasegm1[90] ;
 wire \itasegm1[91] ;
 wire \itasegm1[92] ;
 wire \itasegm1[93] ;
 wire \itasegm1[94] ;
 wire \itasegm1[95] ;
 wire \itasegm1[96] ;
 wire \itasegm1[97] ;
 wire \itasegm1[98] ;
 wire \itasegm1[99] ;
 wire \itasegm1[9] ;
 wire \itasel1[0] ;
 wire \itasel1[100] ;
 wire \itasel1[101] ;
 wire \itasel1[102] ;
 wire \itasel1[103] ;
 wire \itasel1[104] ;
 wire \itasel1[105] ;
 wire \itasel1[106] ;
 wire \itasel1[107] ;
 wire \itasel1[108] ;
 wire \itasel1[109] ;
 wire \itasel1[10] ;
 wire \itasel1[110] ;
 wire \itasel1[111] ;
 wire \itasel1[112] ;
 wire \itasel1[113] ;
 wire \itasel1[114] ;
 wire \itasel1[115] ;
 wire \itasel1[116] ;
 wire \itasel1[117] ;
 wire \itasel1[118] ;
 wire \itasel1[119] ;
 wire \itasel1[11] ;
 wire \itasel1[120] ;
 wire \itasel1[121] ;
 wire \itasel1[122] ;
 wire \itasel1[123] ;
 wire \itasel1[124] ;
 wire \itasel1[125] ;
 wire \itasel1[126] ;
 wire \itasel1[127] ;
 wire \itasel1[128] ;
 wire \itasel1[129] ;
 wire \itasel1[12] ;
 wire \itasel1[130] ;
 wire \itasel1[131] ;
 wire \itasel1[132] ;
 wire \itasel1[133] ;
 wire \itasel1[134] ;
 wire \itasel1[135] ;
 wire \itasel1[136] ;
 wire \itasel1[137] ;
 wire \itasel1[138] ;
 wire \itasel1[139] ;
 wire \itasel1[13] ;
 wire \itasel1[140] ;
 wire \itasel1[141] ;
 wire \itasel1[142] ;
 wire \itasel1[143] ;
 wire \itasel1[144] ;
 wire \itasel1[145] ;
 wire \itasel1[146] ;
 wire \itasel1[147] ;
 wire \itasel1[148] ;
 wire \itasel1[149] ;
 wire \itasel1[14] ;
 wire \itasel1[150] ;
 wire \itasel1[151] ;
 wire \itasel1[152] ;
 wire \itasel1[153] ;
 wire \itasel1[154] ;
 wire \itasel1[155] ;
 wire \itasel1[156] ;
 wire \itasel1[157] ;
 wire \itasel1[158] ;
 wire \itasel1[159] ;
 wire \itasel1[15] ;
 wire \itasel1[160] ;
 wire \itasel1[161] ;
 wire \itasel1[162] ;
 wire \itasel1[163] ;
 wire \itasel1[164] ;
 wire \itasel1[165] ;
 wire \itasel1[166] ;
 wire \itasel1[167] ;
 wire \itasel1[168] ;
 wire \itasel1[169] ;
 wire \itasel1[16] ;
 wire \itasel1[170] ;
 wire \itasel1[171] ;
 wire \itasel1[172] ;
 wire \itasel1[173] ;
 wire \itasel1[174] ;
 wire \itasel1[175] ;
 wire \itasel1[176] ;
 wire \itasel1[177] ;
 wire \itasel1[178] ;
 wire \itasel1[179] ;
 wire \itasel1[17] ;
 wire \itasel1[180] ;
 wire \itasel1[181] ;
 wire \itasel1[182] ;
 wire \itasel1[183] ;
 wire \itasel1[184] ;
 wire \itasel1[185] ;
 wire \itasel1[186] ;
 wire \itasel1[187] ;
 wire \itasel1[188] ;
 wire \itasel1[189] ;
 wire \itasel1[18] ;
 wire \itasel1[190] ;
 wire \itasel1[191] ;
 wire \itasel1[192] ;
 wire \itasel1[193] ;
 wire \itasel1[194] ;
 wire \itasel1[195] ;
 wire \itasel1[196] ;
 wire \itasel1[197] ;
 wire \itasel1[198] ;
 wire \itasel1[199] ;
 wire \itasel1[19] ;
 wire \itasel1[1] ;
 wire \itasel1[200] ;
 wire \itasel1[201] ;
 wire \itasel1[202] ;
 wire \itasel1[203] ;
 wire \itasel1[204] ;
 wire \itasel1[205] ;
 wire \itasel1[206] ;
 wire \itasel1[207] ;
 wire \itasel1[208] ;
 wire \itasel1[209] ;
 wire \itasel1[20] ;
 wire \itasel1[210] ;
 wire \itasel1[211] ;
 wire \itasel1[212] ;
 wire \itasel1[213] ;
 wire \itasel1[214] ;
 wire \itasel1[215] ;
 wire \itasel1[216] ;
 wire \itasel1[217] ;
 wire \itasel1[218] ;
 wire \itasel1[219] ;
 wire \itasel1[21] ;
 wire \itasel1[220] ;
 wire \itasel1[221] ;
 wire \itasel1[222] ;
 wire \itasel1[223] ;
 wire \itasel1[224] ;
 wire \itasel1[225] ;
 wire \itasel1[226] ;
 wire \itasel1[227] ;
 wire \itasel1[228] ;
 wire \itasel1[229] ;
 wire \itasel1[22] ;
 wire \itasel1[230] ;
 wire \itasel1[231] ;
 wire \itasel1[232] ;
 wire \itasel1[233] ;
 wire \itasel1[234] ;
 wire \itasel1[235] ;
 wire \itasel1[236] ;
 wire \itasel1[237] ;
 wire \itasel1[238] ;
 wire \itasel1[239] ;
 wire \itasel1[23] ;
 wire \itasel1[240] ;
 wire \itasel1[241] ;
 wire \itasel1[242] ;
 wire \itasel1[243] ;
 wire \itasel1[244] ;
 wire \itasel1[245] ;
 wire \itasel1[246] ;
 wire \itasel1[247] ;
 wire \itasel1[248] ;
 wire \itasel1[249] ;
 wire \itasel1[24] ;
 wire \itasel1[250] ;
 wire \itasel1[251] ;
 wire \itasel1[252] ;
 wire \itasel1[253] ;
 wire \itasel1[254] ;
 wire \itasel1[255] ;
 wire \itasel1[256] ;
 wire \itasel1[257] ;
 wire \itasel1[258] ;
 wire \itasel1[259] ;
 wire \itasel1[25] ;
 wire \itasel1[260] ;
 wire \itasel1[261] ;
 wire \itasel1[262] ;
 wire \itasel1[263] ;
 wire \itasel1[264] ;
 wire \itasel1[265] ;
 wire \itasel1[266] ;
 wire \itasel1[267] ;
 wire \itasel1[268] ;
 wire \itasel1[269] ;
 wire \itasel1[26] ;
 wire \itasel1[270] ;
 wire \itasel1[271] ;
 wire \itasel1[272] ;
 wire \itasel1[273] ;
 wire \itasel1[274] ;
 wire \itasel1[275] ;
 wire \itasel1[276] ;
 wire \itasel1[277] ;
 wire \itasel1[278] ;
 wire \itasel1[279] ;
 wire \itasel1[27] ;
 wire \itasel1[280] ;
 wire \itasel1[281] ;
 wire \itasel1[282] ;
 wire \itasel1[283] ;
 wire \itasel1[284] ;
 wire \itasel1[285] ;
 wire \itasel1[286] ;
 wire \itasel1[287] ;
 wire \itasel1[288] ;
 wire \itasel1[289] ;
 wire \itasel1[28] ;
 wire \itasel1[290] ;
 wire \itasel1[291] ;
 wire \itasel1[292] ;
 wire \itasel1[293] ;
 wire \itasel1[294] ;
 wire \itasel1[295] ;
 wire \itasel1[296] ;
 wire \itasel1[297] ;
 wire \itasel1[298] ;
 wire \itasel1[299] ;
 wire \itasel1[29] ;
 wire \itasel1[2] ;
 wire \itasel1[300] ;
 wire \itasel1[301] ;
 wire \itasel1[302] ;
 wire \itasel1[303] ;
 wire \itasel1[304] ;
 wire \itasel1[305] ;
 wire \itasel1[306] ;
 wire \itasel1[307] ;
 wire \itasel1[308] ;
 wire \itasel1[309] ;
 wire \itasel1[30] ;
 wire \itasel1[310] ;
 wire \itasel1[311] ;
 wire \itasel1[312] ;
 wire \itasel1[313] ;
 wire \itasel1[314] ;
 wire \itasel1[315] ;
 wire \itasel1[316] ;
 wire \itasel1[317] ;
 wire \itasel1[318] ;
 wire \itasel1[319] ;
 wire \itasel1[31] ;
 wire \itasel1[320] ;
 wire \itasel1[321] ;
 wire \itasel1[322] ;
 wire \itasel1[323] ;
 wire \itasel1[324] ;
 wire \itasel1[325] ;
 wire \itasel1[326] ;
 wire \itasel1[327] ;
 wire \itasel1[328] ;
 wire \itasel1[329] ;
 wire \itasel1[32] ;
 wire \itasel1[330] ;
 wire \itasel1[331] ;
 wire \itasel1[332] ;
 wire \itasel1[333] ;
 wire \itasel1[334] ;
 wire \itasel1[335] ;
 wire \itasel1[336] ;
 wire \itasel1[337] ;
 wire \itasel1[338] ;
 wire \itasel1[339] ;
 wire \itasel1[33] ;
 wire \itasel1[340] ;
 wire \itasel1[341] ;
 wire \itasel1[342] ;
 wire \itasel1[343] ;
 wire \itasel1[344] ;
 wire \itasel1[345] ;
 wire \itasel1[346] ;
 wire \itasel1[347] ;
 wire \itasel1[348] ;
 wire \itasel1[349] ;
 wire \itasel1[34] ;
 wire \itasel1[350] ;
 wire \itasel1[351] ;
 wire \itasel1[352] ;
 wire \itasel1[353] ;
 wire \itasel1[354] ;
 wire \itasel1[355] ;
 wire \itasel1[356] ;
 wire \itasel1[357] ;
 wire \itasel1[358] ;
 wire \itasel1[359] ;
 wire \itasel1[35] ;
 wire \itasel1[360] ;
 wire \itasel1[361] ;
 wire \itasel1[362] ;
 wire \itasel1[363] ;
 wire \itasel1[364] ;
 wire \itasel1[365] ;
 wire \itasel1[366] ;
 wire \itasel1[367] ;
 wire \itasel1[368] ;
 wire \itasel1[369] ;
 wire \itasel1[36] ;
 wire \itasel1[370] ;
 wire \itasel1[371] ;
 wire \itasel1[372] ;
 wire \itasel1[373] ;
 wire \itasel1[374] ;
 wire \itasel1[375] ;
 wire \itasel1[376] ;
 wire \itasel1[377] ;
 wire \itasel1[378] ;
 wire \itasel1[379] ;
 wire \itasel1[37] ;
 wire \itasel1[380] ;
 wire \itasel1[381] ;
 wire \itasel1[382] ;
 wire \itasel1[383] ;
 wire \itasel1[384] ;
 wire \itasel1[385] ;
 wire \itasel1[386] ;
 wire \itasel1[387] ;
 wire \itasel1[388] ;
 wire \itasel1[389] ;
 wire \itasel1[38] ;
 wire \itasel1[390] ;
 wire \itasel1[391] ;
 wire \itasel1[392] ;
 wire \itasel1[393] ;
 wire \itasel1[394] ;
 wire \itasel1[395] ;
 wire \itasel1[396] ;
 wire \itasel1[397] ;
 wire \itasel1[398] ;
 wire \itasel1[399] ;
 wire \itasel1[39] ;
 wire \itasel1[3] ;
 wire \itasel1[400] ;
 wire \itasel1[401] ;
 wire \itasel1[402] ;
 wire \itasel1[403] ;
 wire \itasel1[404] ;
 wire \itasel1[405] ;
 wire \itasel1[406] ;
 wire \itasel1[407] ;
 wire \itasel1[408] ;
 wire \itasel1[409] ;
 wire \itasel1[40] ;
 wire \itasel1[410] ;
 wire \itasel1[411] ;
 wire \itasel1[412] ;
 wire \itasel1[413] ;
 wire \itasel1[414] ;
 wire \itasel1[415] ;
 wire \itasel1[416] ;
 wire \itasel1[417] ;
 wire \itasel1[418] ;
 wire \itasel1[419] ;
 wire \itasel1[41] ;
 wire \itasel1[420] ;
 wire \itasel1[421] ;
 wire \itasel1[422] ;
 wire \itasel1[423] ;
 wire \itasel1[424] ;
 wire \itasel1[425] ;
 wire \itasel1[426] ;
 wire \itasel1[427] ;
 wire \itasel1[428] ;
 wire \itasel1[429] ;
 wire \itasel1[42] ;
 wire \itasel1[430] ;
 wire \itasel1[431] ;
 wire \itasel1[432] ;
 wire \itasel1[433] ;
 wire \itasel1[434] ;
 wire \itasel1[435] ;
 wire \itasel1[436] ;
 wire \itasel1[437] ;
 wire \itasel1[438] ;
 wire \itasel1[439] ;
 wire \itasel1[43] ;
 wire \itasel1[440] ;
 wire \itasel1[441] ;
 wire \itasel1[442] ;
 wire \itasel1[443] ;
 wire \itasel1[444] ;
 wire \itasel1[445] ;
 wire \itasel1[446] ;
 wire \itasel1[447] ;
 wire \itasel1[448] ;
 wire \itasel1[449] ;
 wire \itasel1[44] ;
 wire \itasel1[450] ;
 wire \itasel1[451] ;
 wire \itasel1[452] ;
 wire \itasel1[453] ;
 wire \itasel1[454] ;
 wire \itasel1[455] ;
 wire \itasel1[456] ;
 wire \itasel1[457] ;
 wire \itasel1[458] ;
 wire \itasel1[459] ;
 wire \itasel1[45] ;
 wire \itasel1[460] ;
 wire \itasel1[461] ;
 wire \itasel1[462] ;
 wire \itasel1[463] ;
 wire \itasel1[464] ;
 wire \itasel1[465] ;
 wire \itasel1[466] ;
 wire \itasel1[467] ;
 wire \itasel1[468] ;
 wire \itasel1[469] ;
 wire \itasel1[46] ;
 wire \itasel1[470] ;
 wire \itasel1[471] ;
 wire \itasel1[472] ;
 wire \itasel1[473] ;
 wire \itasel1[474] ;
 wire \itasel1[475] ;
 wire \itasel1[476] ;
 wire \itasel1[477] ;
 wire \itasel1[478] ;
 wire \itasel1[479] ;
 wire \itasel1[47] ;
 wire \itasel1[480] ;
 wire \itasel1[481] ;
 wire \itasel1[482] ;
 wire \itasel1[483] ;
 wire \itasel1[484] ;
 wire \itasel1[485] ;
 wire \itasel1[486] ;
 wire \itasel1[487] ;
 wire \itasel1[488] ;
 wire \itasel1[489] ;
 wire \itasel1[48] ;
 wire \itasel1[490] ;
 wire \itasel1[491] ;
 wire \itasel1[492] ;
 wire \itasel1[493] ;
 wire \itasel1[494] ;
 wire \itasel1[495] ;
 wire \itasel1[496] ;
 wire \itasel1[497] ;
 wire \itasel1[498] ;
 wire \itasel1[499] ;
 wire \itasel1[49] ;
 wire \itasel1[4] ;
 wire \itasel1[500] ;
 wire \itasel1[501] ;
 wire \itasel1[502] ;
 wire \itasel1[503] ;
 wire \itasel1[504] ;
 wire \itasel1[505] ;
 wire \itasel1[506] ;
 wire \itasel1[507] ;
 wire \itasel1[508] ;
 wire \itasel1[509] ;
 wire \itasel1[50] ;
 wire \itasel1[510] ;
 wire \itasel1[511] ;
 wire \itasel1[512] ;
 wire \itasel1[513] ;
 wire \itasel1[514] ;
 wire \itasel1[515] ;
 wire \itasel1[516] ;
 wire \itasel1[517] ;
 wire \itasel1[518] ;
 wire \itasel1[519] ;
 wire \itasel1[51] ;
 wire \itasel1[520] ;
 wire \itasel1[521] ;
 wire \itasel1[522] ;
 wire \itasel1[523] ;
 wire \itasel1[524] ;
 wire \itasel1[525] ;
 wire \itasel1[526] ;
 wire \itasel1[527] ;
 wire \itasel1[528] ;
 wire \itasel1[529] ;
 wire \itasel1[52] ;
 wire \itasel1[530] ;
 wire \itasel1[531] ;
 wire \itasel1[532] ;
 wire \itasel1[533] ;
 wire \itasel1[534] ;
 wire \itasel1[535] ;
 wire \itasel1[536] ;
 wire \itasel1[537] ;
 wire \itasel1[538] ;
 wire \itasel1[539] ;
 wire \itasel1[53] ;
 wire \itasel1[540] ;
 wire \itasel1[541] ;
 wire \itasel1[542] ;
 wire \itasel1[543] ;
 wire \itasel1[544] ;
 wire \itasel1[545] ;
 wire \itasel1[546] ;
 wire \itasel1[547] ;
 wire \itasel1[548] ;
 wire \itasel1[549] ;
 wire \itasel1[54] ;
 wire \itasel1[550] ;
 wire \itasel1[551] ;
 wire \itasel1[552] ;
 wire \itasel1[553] ;
 wire \itasel1[554] ;
 wire \itasel1[555] ;
 wire \itasel1[556] ;
 wire \itasel1[557] ;
 wire \itasel1[558] ;
 wire \itasel1[559] ;
 wire \itasel1[55] ;
 wire \itasel1[560] ;
 wire \itasel1[561] ;
 wire \itasel1[562] ;
 wire \itasel1[563] ;
 wire \itasel1[564] ;
 wire \itasel1[565] ;
 wire \itasel1[566] ;
 wire \itasel1[567] ;
 wire \itasel1[568] ;
 wire \itasel1[569] ;
 wire \itasel1[56] ;
 wire \itasel1[570] ;
 wire \itasel1[571] ;
 wire \itasel1[572] ;
 wire \itasel1[573] ;
 wire \itasel1[574] ;
 wire \itasel1[575] ;
 wire \itasel1[576] ;
 wire \itasel1[577] ;
 wire \itasel1[578] ;
 wire \itasel1[579] ;
 wire \itasel1[57] ;
 wire \itasel1[580] ;
 wire \itasel1[581] ;
 wire \itasel1[582] ;
 wire \itasel1[583] ;
 wire \itasel1[584] ;
 wire \itasel1[585] ;
 wire \itasel1[586] ;
 wire \itasel1[587] ;
 wire \itasel1[588] ;
 wire \itasel1[589] ;
 wire \itasel1[58] ;
 wire \itasel1[590] ;
 wire \itasel1[591] ;
 wire \itasel1[592] ;
 wire \itasel1[593] ;
 wire \itasel1[594] ;
 wire \itasel1[595] ;
 wire \itasel1[596] ;
 wire \itasel1[597] ;
 wire \itasel1[598] ;
 wire \itasel1[599] ;
 wire \itasel1[59] ;
 wire \itasel1[5] ;
 wire \itasel1[600] ;
 wire \itasel1[601] ;
 wire \itasel1[602] ;
 wire \itasel1[603] ;
 wire \itasel1[604] ;
 wire \itasel1[605] ;
 wire \itasel1[606] ;
 wire \itasel1[607] ;
 wire \itasel1[608] ;
 wire \itasel1[609] ;
 wire \itasel1[60] ;
 wire \itasel1[610] ;
 wire \itasel1[611] ;
 wire \itasel1[612] ;
 wire \itasel1[613] ;
 wire \itasel1[614] ;
 wire \itasel1[615] ;
 wire \itasel1[616] ;
 wire \itasel1[617] ;
 wire \itasel1[618] ;
 wire \itasel1[619] ;
 wire \itasel1[61] ;
 wire \itasel1[620] ;
 wire \itasel1[621] ;
 wire \itasel1[622] ;
 wire \itasel1[623] ;
 wire \itasel1[624] ;
 wire \itasel1[625] ;
 wire \itasel1[626] ;
 wire \itasel1[627] ;
 wire \itasel1[628] ;
 wire \itasel1[629] ;
 wire \itasel1[62] ;
 wire \itasel1[630] ;
 wire \itasel1[631] ;
 wire \itasel1[632] ;
 wire \itasel1[633] ;
 wire \itasel1[634] ;
 wire \itasel1[635] ;
 wire \itasel1[636] ;
 wire \itasel1[637] ;
 wire \itasel1[638] ;
 wire \itasel1[639] ;
 wire \itasel1[63] ;
 wire \itasel1[640] ;
 wire \itasel1[641] ;
 wire \itasel1[642] ;
 wire \itasel1[643] ;
 wire \itasel1[644] ;
 wire \itasel1[645] ;
 wire \itasel1[646] ;
 wire \itasel1[647] ;
 wire \itasel1[648] ;
 wire \itasel1[649] ;
 wire \itasel1[64] ;
 wire \itasel1[650] ;
 wire \itasel1[651] ;
 wire \itasel1[652] ;
 wire \itasel1[653] ;
 wire \itasel1[654] ;
 wire \itasel1[655] ;
 wire \itasel1[656] ;
 wire \itasel1[657] ;
 wire \itasel1[658] ;
 wire \itasel1[659] ;
 wire \itasel1[65] ;
 wire \itasel1[660] ;
 wire \itasel1[661] ;
 wire \itasel1[662] ;
 wire \itasel1[663] ;
 wire \itasel1[664] ;
 wire \itasel1[665] ;
 wire \itasel1[666] ;
 wire \itasel1[667] ;
 wire \itasel1[668] ;
 wire \itasel1[669] ;
 wire \itasel1[66] ;
 wire \itasel1[670] ;
 wire \itasel1[671] ;
 wire \itasel1[672] ;
 wire \itasel1[673] ;
 wire \itasel1[674] ;
 wire \itasel1[675] ;
 wire \itasel1[676] ;
 wire \itasel1[677] ;
 wire \itasel1[678] ;
 wire \itasel1[679] ;
 wire \itasel1[67] ;
 wire \itasel1[680] ;
 wire \itasel1[681] ;
 wire \itasel1[682] ;
 wire \itasel1[683] ;
 wire \itasel1[684] ;
 wire \itasel1[685] ;
 wire \itasel1[686] ;
 wire \itasel1[687] ;
 wire \itasel1[688] ;
 wire \itasel1[689] ;
 wire \itasel1[68] ;
 wire \itasel1[690] ;
 wire \itasel1[691] ;
 wire \itasel1[692] ;
 wire \itasel1[693] ;
 wire \itasel1[694] ;
 wire \itasel1[695] ;
 wire \itasel1[696] ;
 wire \itasel1[697] ;
 wire \itasel1[698] ;
 wire \itasel1[699] ;
 wire \itasel1[69] ;
 wire \itasel1[6] ;
 wire \itasel1[700] ;
 wire \itasel1[701] ;
 wire \itasel1[702] ;
 wire \itasel1[703] ;
 wire \itasel1[704] ;
 wire \itasel1[705] ;
 wire \itasel1[706] ;
 wire \itasel1[707] ;
 wire \itasel1[708] ;
 wire \itasel1[709] ;
 wire \itasel1[70] ;
 wire \itasel1[710] ;
 wire \itasel1[711] ;
 wire \itasel1[712] ;
 wire \itasel1[713] ;
 wire \itasel1[714] ;
 wire \itasel1[715] ;
 wire \itasel1[716] ;
 wire \itasel1[717] ;
 wire \itasel1[718] ;
 wire \itasel1[719] ;
 wire \itasel1[71] ;
 wire \itasel1[720] ;
 wire \itasel1[721] ;
 wire \itasel1[722] ;
 wire \itasel1[723] ;
 wire \itasel1[724] ;
 wire \itasel1[725] ;
 wire \itasel1[726] ;
 wire \itasel1[727] ;
 wire \itasel1[728] ;
 wire \itasel1[729] ;
 wire \itasel1[72] ;
 wire \itasel1[730] ;
 wire \itasel1[731] ;
 wire \itasel1[732] ;
 wire \itasel1[733] ;
 wire \itasel1[734] ;
 wire \itasel1[735] ;
 wire \itasel1[736] ;
 wire \itasel1[737] ;
 wire \itasel1[738] ;
 wire \itasel1[739] ;
 wire \itasel1[73] ;
 wire \itasel1[740] ;
 wire \itasel1[741] ;
 wire \itasel1[742] ;
 wire \itasel1[743] ;
 wire \itasel1[744] ;
 wire \itasel1[745] ;
 wire \itasel1[746] ;
 wire \itasel1[747] ;
 wire \itasel1[748] ;
 wire \itasel1[749] ;
 wire \itasel1[74] ;
 wire \itasel1[750] ;
 wire \itasel1[751] ;
 wire \itasel1[752] ;
 wire \itasel1[753] ;
 wire \itasel1[754] ;
 wire \itasel1[755] ;
 wire \itasel1[756] ;
 wire \itasel1[757] ;
 wire \itasel1[758] ;
 wire \itasel1[759] ;
 wire \itasel1[75] ;
 wire \itasel1[760] ;
 wire \itasel1[761] ;
 wire \itasel1[762] ;
 wire \itasel1[763] ;
 wire \itasel1[764] ;
 wire \itasel1[765] ;
 wire \itasel1[766] ;
 wire \itasel1[767] ;
 wire \itasel1[76] ;
 wire \itasel1[77] ;
 wire \itasel1[78] ;
 wire \itasel1[79] ;
 wire \itasel1[7] ;
 wire \itasel1[80] ;
 wire \itasel1[81] ;
 wire \itasel1[82] ;
 wire \itasel1[83] ;
 wire \itasel1[84] ;
 wire \itasel1[85] ;
 wire \itasel1[86] ;
 wire \itasel1[87] ;
 wire \itasel1[88] ;
 wire \itasel1[89] ;
 wire \itasel1[8] ;
 wire \itasel1[90] ;
 wire \itasel1[91] ;
 wire \itasel1[92] ;
 wire \itasel1[93] ;
 wire \itasel1[94] ;
 wire \itasel1[95] ;
 wire \itasel1[96] ;
 wire \itasel1[97] ;
 wire \itasel1[98] ;
 wire \itasel1[99] ;
 wire \itasel1[9] ;

 ita ita (.clk(wb_clk_i),
    .io_oeb({io_oeb[37],
    io_oeb[36],
    io_oeb[35],
    io_oeb[34],
    io_oeb[33],
    io_oeb[32],
    io_oeb[31],
    io_oeb[30],
    io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24],
    io_oeb[23],
    io_oeb[22],
    io_oeb[21],
    io_oeb[20],
    io_oeb[19],
    io_oeb[18],
    io_oeb[17],
    io_oeb[16],
    io_oeb[15],
    io_oeb[14],
    io_oeb[13],
    io_oeb[12],
    io_oeb[11],
    io_oeb[10],
    io_oeb[9],
    io_oeb[8],
    io_oeb[7],
    io_oeb[6],
    io_oeb[5],
    io_oeb[4],
    io_oeb[3],
    io_oeb[2],
    io_oeb[1],
    io_oeb[0]}),
    .itasegm({\itasegm1[895] ,
    \itasegm1[894] ,
    \itasegm1[893] ,
    \itasegm1[892] ,
    \itasegm1[891] ,
    \itasegm1[890] ,
    \itasegm1[889] ,
    \itasegm1[888] ,
    \itasegm1[887] ,
    \itasegm1[886] ,
    \itasegm1[885] ,
    \itasegm1[884] ,
    \itasegm1[883] ,
    \itasegm1[882] ,
    \itasegm1[881] ,
    \itasegm1[880] ,
    \itasegm1[879] ,
    \itasegm1[878] ,
    \itasegm1[877] ,
    \itasegm1[876] ,
    \itasegm1[875] ,
    \itasegm1[874] ,
    \itasegm1[873] ,
    \itasegm1[872] ,
    \itasegm1[871] ,
    \itasegm1[870] ,
    \itasegm1[869] ,
    \itasegm1[868] ,
    \itasegm1[867] ,
    \itasegm1[866] ,
    \itasegm1[865] ,
    \itasegm1[864] ,
    \itasegm1[863] ,
    \itasegm1[862] ,
    \itasegm1[861] ,
    \itasegm1[860] ,
    \itasegm1[859] ,
    \itasegm1[858] ,
    \itasegm1[857] ,
    \itasegm1[856] ,
    \itasegm1[855] ,
    \itasegm1[854] ,
    \itasegm1[853] ,
    \itasegm1[852] ,
    \itasegm1[851] ,
    \itasegm1[850] ,
    \itasegm1[849] ,
    \itasegm1[848] ,
    \itasegm1[847] ,
    \itasegm1[846] ,
    \itasegm1[845] ,
    \itasegm1[844] ,
    \itasegm1[843] ,
    \itasegm1[842] ,
    \itasegm1[841] ,
    \itasegm1[840] ,
    \itasegm1[839] ,
    \itasegm1[838] ,
    \itasegm1[837] ,
    \itasegm1[836] ,
    \itasegm1[835] ,
    \itasegm1[834] ,
    \itasegm1[833] ,
    \itasegm1[832] ,
    \itasegm1[831] ,
    \itasegm1[830] ,
    \itasegm1[829] ,
    \itasegm1[828] ,
    \itasegm1[827] ,
    \itasegm1[826] ,
    \itasegm1[825] ,
    \itasegm1[824] ,
    \itasegm1[823] ,
    \itasegm1[822] ,
    \itasegm1[821] ,
    \itasegm1[820] ,
    \itasegm1[819] ,
    \itasegm1[818] ,
    \itasegm1[817] ,
    \itasegm1[816] ,
    \itasegm1[815] ,
    \itasegm1[814] ,
    \itasegm1[813] ,
    \itasegm1[812] ,
    \itasegm1[811] ,
    \itasegm1[810] ,
    \itasegm1[809] ,
    \itasegm1[808] ,
    \itasegm1[807] ,
    \itasegm1[806] ,
    \itasegm1[805] ,
    \itasegm1[804] ,
    \itasegm1[803] ,
    \itasegm1[802] ,
    \itasegm1[801] ,
    \itasegm1[800] ,
    \itasegm1[799] ,
    \itasegm1[798] ,
    \itasegm1[797] ,
    \itasegm1[796] ,
    \itasegm1[795] ,
    \itasegm1[794] ,
    \itasegm1[793] ,
    \itasegm1[792] ,
    \itasegm1[791] ,
    \itasegm1[790] ,
    \itasegm1[789] ,
    \itasegm1[788] ,
    \itasegm1[787] ,
    \itasegm1[786] ,
    \itasegm1[785] ,
    \itasegm1[784] ,
    \itasegm1[783] ,
    \itasegm1[782] ,
    \itasegm1[781] ,
    \itasegm1[780] ,
    \itasegm1[779] ,
    \itasegm1[778] ,
    \itasegm1[777] ,
    \itasegm1[776] ,
    \itasegm1[775] ,
    \itasegm1[774] ,
    \itasegm1[773] ,
    \itasegm1[772] ,
    \itasegm1[771] ,
    \itasegm1[770] ,
    \itasegm1[769] ,
    \itasegm1[768] ,
    \itasegm1[767] ,
    \itasegm1[766] ,
    \itasegm1[765] ,
    \itasegm1[764] ,
    \itasegm1[763] ,
    \itasegm1[762] ,
    \itasegm1[761] ,
    \itasegm1[760] ,
    \itasegm1[759] ,
    \itasegm1[758] ,
    \itasegm1[757] ,
    \itasegm1[756] ,
    \itasegm1[755] ,
    \itasegm1[754] ,
    \itasegm1[753] ,
    \itasegm1[752] ,
    \itasegm1[751] ,
    \itasegm1[750] ,
    \itasegm1[749] ,
    \itasegm1[748] ,
    \itasegm1[747] ,
    \itasegm1[746] ,
    \itasegm1[745] ,
    \itasegm1[744] ,
    \itasegm1[743] ,
    \itasegm1[742] ,
    \itasegm1[741] ,
    \itasegm1[740] ,
    \itasegm1[739] ,
    \itasegm1[738] ,
    \itasegm1[737] ,
    \itasegm1[736] ,
    \itasegm1[735] ,
    \itasegm1[734] ,
    \itasegm1[733] ,
    \itasegm1[732] ,
    \itasegm1[731] ,
    \itasegm1[730] ,
    \itasegm1[729] ,
    \itasegm1[728] ,
    \itasegm1[727] ,
    \itasegm1[726] ,
    \itasegm1[725] ,
    \itasegm1[724] ,
    \itasegm1[723] ,
    \itasegm1[722] ,
    \itasegm1[721] ,
    \itasegm1[720] ,
    \itasegm1[719] ,
    \itasegm1[718] ,
    \itasegm1[717] ,
    \itasegm1[716] ,
    \itasegm1[715] ,
    \itasegm1[714] ,
    \itasegm1[713] ,
    \itasegm1[712] ,
    \itasegm1[711] ,
    \itasegm1[710] ,
    \itasegm1[709] ,
    \itasegm1[708] ,
    \itasegm1[707] ,
    \itasegm1[706] ,
    \itasegm1[705] ,
    \itasegm1[704] ,
    \itasegm1[703] ,
    \itasegm1[702] ,
    \itasegm1[701] ,
    \itasegm1[700] ,
    \itasegm1[699] ,
    \itasegm1[698] ,
    \itasegm1[697] ,
    \itasegm1[696] ,
    \itasegm1[695] ,
    \itasegm1[694] ,
    \itasegm1[693] ,
    \itasegm1[692] ,
    \itasegm1[691] ,
    \itasegm1[690] ,
    \itasegm1[689] ,
    \itasegm1[688] ,
    \itasegm1[687] ,
    \itasegm1[686] ,
    \itasegm1[685] ,
    \itasegm1[684] ,
    \itasegm1[683] ,
    \itasegm1[682] ,
    \itasegm1[681] ,
    \itasegm1[680] ,
    \itasegm1[679] ,
    \itasegm1[678] ,
    \itasegm1[677] ,
    \itasegm1[676] ,
    \itasegm1[675] ,
    \itasegm1[674] ,
    \itasegm1[673] ,
    \itasegm1[672] ,
    \itasegm1[671] ,
    \itasegm1[670] ,
    \itasegm1[669] ,
    \itasegm1[668] ,
    \itasegm1[667] ,
    \itasegm1[666] ,
    \itasegm1[665] ,
    \itasegm1[664] ,
    \itasegm1[663] ,
    \itasegm1[662] ,
    \itasegm1[661] ,
    \itasegm1[660] ,
    \itasegm1[659] ,
    \itasegm1[658] ,
    \itasegm1[657] ,
    \itasegm1[656] ,
    \itasegm1[655] ,
    \itasegm1[654] ,
    \itasegm1[653] ,
    \itasegm1[652] ,
    \itasegm1[651] ,
    \itasegm1[650] ,
    \itasegm1[649] ,
    \itasegm1[648] ,
    \itasegm1[647] ,
    \itasegm1[646] ,
    \itasegm1[645] ,
    \itasegm1[644] ,
    \itasegm1[643] ,
    \itasegm1[642] ,
    \itasegm1[641] ,
    \itasegm1[640] ,
    \itasegm1[639] ,
    \itasegm1[638] ,
    \itasegm1[637] ,
    \itasegm1[636] ,
    \itasegm1[635] ,
    \itasegm1[634] ,
    \itasegm1[633] ,
    \itasegm1[632] ,
    \itasegm1[631] ,
    \itasegm1[630] ,
    \itasegm1[629] ,
    \itasegm1[628] ,
    \itasegm1[627] ,
    \itasegm1[626] ,
    \itasegm1[625] ,
    \itasegm1[624] ,
    \itasegm1[623] ,
    \itasegm1[622] ,
    \itasegm1[621] ,
    \itasegm1[620] ,
    \itasegm1[619] ,
    \itasegm1[618] ,
    \itasegm1[617] ,
    \itasegm1[616] ,
    \itasegm1[615] ,
    \itasegm1[614] ,
    \itasegm1[613] ,
    \itasegm1[612] ,
    \itasegm1[611] ,
    \itasegm1[610] ,
    \itasegm1[609] ,
    \itasegm1[608] ,
    \itasegm1[607] ,
    \itasegm1[606] ,
    \itasegm1[605] ,
    \itasegm1[604] ,
    \itasegm1[603] ,
    \itasegm1[602] ,
    \itasegm1[601] ,
    \itasegm1[600] ,
    \itasegm1[599] ,
    \itasegm1[598] ,
    \itasegm1[597] ,
    \itasegm1[596] ,
    \itasegm1[595] ,
    \itasegm1[594] ,
    \itasegm1[593] ,
    \itasegm1[592] ,
    \itasegm1[591] ,
    \itasegm1[590] ,
    \itasegm1[589] ,
    \itasegm1[588] ,
    \itasegm1[587] ,
    \itasegm1[586] ,
    \itasegm1[585] ,
    \itasegm1[584] ,
    \itasegm1[583] ,
    \itasegm1[582] ,
    \itasegm1[581] ,
    \itasegm1[580] ,
    \itasegm1[579] ,
    \itasegm1[578] ,
    \itasegm1[577] ,
    \itasegm1[576] ,
    \itasegm1[575] ,
    \itasegm1[574] ,
    \itasegm1[573] ,
    \itasegm1[572] ,
    \itasegm1[571] ,
    \itasegm1[570] ,
    \itasegm1[569] ,
    \itasegm1[568] ,
    \itasegm1[567] ,
    \itasegm1[566] ,
    \itasegm1[565] ,
    \itasegm1[564] ,
    \itasegm1[563] ,
    \itasegm1[562] ,
    \itasegm1[561] ,
    \itasegm1[560] ,
    \itasegm1[559] ,
    \itasegm1[558] ,
    \itasegm1[557] ,
    \itasegm1[556] ,
    \itasegm1[555] ,
    \itasegm1[554] ,
    \itasegm1[553] ,
    \itasegm1[552] ,
    \itasegm1[551] ,
    \itasegm1[550] ,
    \itasegm1[549] ,
    \itasegm1[548] ,
    \itasegm1[547] ,
    \itasegm1[546] ,
    \itasegm1[545] ,
    \itasegm1[544] ,
    \itasegm1[543] ,
    \itasegm1[542] ,
    \itasegm1[541] ,
    \itasegm1[540] ,
    \itasegm1[539] ,
    \itasegm1[538] ,
    \itasegm1[537] ,
    \itasegm1[536] ,
    \itasegm1[535] ,
    \itasegm1[534] ,
    \itasegm1[533] ,
    \itasegm1[532] ,
    \itasegm1[531] ,
    \itasegm1[530] ,
    \itasegm1[529] ,
    \itasegm1[528] ,
    \itasegm1[527] ,
    \itasegm1[526] ,
    \itasegm1[525] ,
    \itasegm1[524] ,
    \itasegm1[523] ,
    \itasegm1[522] ,
    \itasegm1[521] ,
    \itasegm1[520] ,
    \itasegm1[519] ,
    \itasegm1[518] ,
    \itasegm1[517] ,
    \itasegm1[516] ,
    \itasegm1[515] ,
    \itasegm1[514] ,
    \itasegm1[513] ,
    \itasegm1[512] ,
    \itasegm1[511] ,
    \itasegm1[510] ,
    \itasegm1[509] ,
    \itasegm1[508] ,
    \itasegm1[507] ,
    \itasegm1[506] ,
    \itasegm1[505] ,
    \itasegm1[504] ,
    \itasegm1[503] ,
    \itasegm1[502] ,
    \itasegm1[501] ,
    \itasegm1[500] ,
    \itasegm1[499] ,
    \itasegm1[498] ,
    \itasegm1[497] ,
    \itasegm1[496] ,
    \itasegm1[495] ,
    \itasegm1[494] ,
    \itasegm1[493] ,
    \itasegm1[492] ,
    \itasegm1[491] ,
    \itasegm1[490] ,
    \itasegm1[489] ,
    \itasegm1[488] ,
    \itasegm1[487] ,
    \itasegm1[486] ,
    \itasegm1[485] ,
    \itasegm1[484] ,
    \itasegm1[483] ,
    \itasegm1[482] ,
    \itasegm1[481] ,
    \itasegm1[480] ,
    \itasegm1[479] ,
    \itasegm1[478] ,
    \itasegm1[477] ,
    \itasegm1[476] ,
    \itasegm1[475] ,
    \itasegm1[474] ,
    \itasegm1[473] ,
    \itasegm1[472] ,
    \itasegm1[471] ,
    \itasegm1[470] ,
    \itasegm1[469] ,
    \itasegm1[468] ,
    \itasegm1[467] ,
    \itasegm1[466] ,
    \itasegm1[465] ,
    \itasegm1[464] ,
    \itasegm1[463] ,
    \itasegm1[462] ,
    \itasegm1[461] ,
    \itasegm1[460] ,
    \itasegm1[459] ,
    \itasegm1[458] ,
    \itasegm1[457] ,
    \itasegm1[456] ,
    \itasegm1[455] ,
    \itasegm1[454] ,
    \itasegm1[453] ,
    \itasegm1[452] ,
    \itasegm1[451] ,
    \itasegm1[450] ,
    \itasegm1[449] ,
    \itasegm1[448] ,
    \itasegm1[447] ,
    \itasegm1[446] ,
    \itasegm1[445] ,
    \itasegm1[444] ,
    \itasegm1[443] ,
    \itasegm1[442] ,
    \itasegm1[441] ,
    \itasegm1[440] ,
    \itasegm1[439] ,
    \itasegm1[438] ,
    \itasegm1[437] ,
    \itasegm1[436] ,
    \itasegm1[435] ,
    \itasegm1[434] ,
    \itasegm1[433] ,
    \itasegm1[432] ,
    \itasegm1[431] ,
    \itasegm1[430] ,
    \itasegm1[429] ,
    \itasegm1[428] ,
    \itasegm1[427] ,
    \itasegm1[426] ,
    \itasegm1[425] ,
    \itasegm1[424] ,
    \itasegm1[423] ,
    \itasegm1[422] ,
    \itasegm1[421] ,
    \itasegm1[420] ,
    \itasegm1[419] ,
    \itasegm1[418] ,
    \itasegm1[417] ,
    \itasegm1[416] ,
    \itasegm1[415] ,
    \itasegm1[414] ,
    \itasegm1[413] ,
    \itasegm1[412] ,
    \itasegm1[411] ,
    \itasegm1[410] ,
    \itasegm1[409] ,
    \itasegm1[408] ,
    \itasegm1[407] ,
    \itasegm1[406] ,
    \itasegm1[405] ,
    \itasegm1[404] ,
    \itasegm1[403] ,
    \itasegm1[402] ,
    \itasegm1[401] ,
    \itasegm1[400] ,
    \itasegm1[399] ,
    \itasegm1[398] ,
    \itasegm1[397] ,
    \itasegm1[396] ,
    \itasegm1[395] ,
    \itasegm1[394] ,
    \itasegm1[393] ,
    \itasegm1[392] ,
    \itasegm1[391] ,
    \itasegm1[390] ,
    \itasegm1[389] ,
    \itasegm1[388] ,
    \itasegm1[387] ,
    \itasegm1[386] ,
    \itasegm1[385] ,
    \itasegm1[384] ,
    \itasegm1[383] ,
    \itasegm1[382] ,
    \itasegm1[381] ,
    \itasegm1[380] ,
    \itasegm1[379] ,
    \itasegm1[378] ,
    \itasegm1[377] ,
    \itasegm1[376] ,
    \itasegm1[375] ,
    \itasegm1[374] ,
    \itasegm1[373] ,
    \itasegm1[372] ,
    \itasegm1[371] ,
    \itasegm1[370] ,
    \itasegm1[369] ,
    \itasegm1[368] ,
    \itasegm1[367] ,
    \itasegm1[366] ,
    \itasegm1[365] ,
    \itasegm1[364] ,
    \itasegm1[363] ,
    \itasegm1[362] ,
    \itasegm1[361] ,
    \itasegm1[360] ,
    \itasegm1[359] ,
    \itasegm1[358] ,
    \itasegm1[357] ,
    \itasegm1[356] ,
    \itasegm1[355] ,
    \itasegm1[354] ,
    \itasegm1[353] ,
    \itasegm1[352] ,
    \itasegm1[351] ,
    \itasegm1[350] ,
    \itasegm1[349] ,
    \itasegm1[348] ,
    \itasegm1[347] ,
    \itasegm1[346] ,
    \itasegm1[345] ,
    \itasegm1[344] ,
    \itasegm1[343] ,
    \itasegm1[342] ,
    \itasegm1[341] ,
    \itasegm1[340] ,
    \itasegm1[339] ,
    \itasegm1[338] ,
    \itasegm1[337] ,
    \itasegm1[336] ,
    \itasegm1[335] ,
    \itasegm1[334] ,
    \itasegm1[333] ,
    \itasegm1[332] ,
    \itasegm1[331] ,
    \itasegm1[330] ,
    \itasegm1[329] ,
    \itasegm1[328] ,
    \itasegm1[327] ,
    \itasegm1[326] ,
    \itasegm1[325] ,
    \itasegm1[324] ,
    \itasegm1[323] ,
    \itasegm1[322] ,
    \itasegm1[321] ,
    \itasegm1[320] ,
    \itasegm1[319] ,
    \itasegm1[318] ,
    \itasegm1[317] ,
    \itasegm1[316] ,
    \itasegm1[315] ,
    \itasegm1[314] ,
    \itasegm1[313] ,
    \itasegm1[312] ,
    \itasegm1[311] ,
    \itasegm1[310] ,
    \itasegm1[309] ,
    \itasegm1[308] ,
    \itasegm1[307] ,
    \itasegm1[306] ,
    \itasegm1[305] ,
    \itasegm1[304] ,
    \itasegm1[303] ,
    \itasegm1[302] ,
    \itasegm1[301] ,
    \itasegm1[300] ,
    \itasegm1[299] ,
    \itasegm1[298] ,
    \itasegm1[297] ,
    \itasegm1[296] ,
    \itasegm1[295] ,
    \itasegm1[294] ,
    \itasegm1[293] ,
    \itasegm1[292] ,
    \itasegm1[291] ,
    \itasegm1[290] ,
    \itasegm1[289] ,
    \itasegm1[288] ,
    \itasegm1[287] ,
    \itasegm1[286] ,
    \itasegm1[285] ,
    \itasegm1[284] ,
    \itasegm1[283] ,
    \itasegm1[282] ,
    \itasegm1[281] ,
    \itasegm1[280] ,
    \itasegm1[279] ,
    \itasegm1[278] ,
    \itasegm1[277] ,
    \itasegm1[276] ,
    \itasegm1[275] ,
    \itasegm1[274] ,
    \itasegm1[273] ,
    \itasegm1[272] ,
    \itasegm1[271] ,
    \itasegm1[270] ,
    \itasegm1[269] ,
    \itasegm1[268] ,
    \itasegm1[267] ,
    \itasegm1[266] ,
    \itasegm1[265] ,
    \itasegm1[264] ,
    \itasegm1[263] ,
    \itasegm1[262] ,
    \itasegm1[261] ,
    \itasegm1[260] ,
    \itasegm1[259] ,
    \itasegm1[258] ,
    \itasegm1[257] ,
    \itasegm1[256] ,
    \itasegm1[255] ,
    \itasegm1[254] ,
    \itasegm1[253] ,
    \itasegm1[252] ,
    \itasegm1[251] ,
    \itasegm1[250] ,
    \itasegm1[249] ,
    \itasegm1[248] ,
    \itasegm1[247] ,
    \itasegm1[246] ,
    \itasegm1[245] ,
    \itasegm1[244] ,
    \itasegm1[243] ,
    \itasegm1[242] ,
    \itasegm1[241] ,
    \itasegm1[240] ,
    \itasegm1[239] ,
    \itasegm1[238] ,
    \itasegm1[237] ,
    \itasegm1[236] ,
    \itasegm1[235] ,
    \itasegm1[234] ,
    \itasegm1[233] ,
    \itasegm1[232] ,
    \itasegm1[231] ,
    \itasegm1[230] ,
    \itasegm1[229] ,
    \itasegm1[228] ,
    \itasegm1[227] ,
    \itasegm1[226] ,
    \itasegm1[225] ,
    \itasegm1[224] ,
    \itasegm1[223] ,
    \itasegm1[222] ,
    \itasegm1[221] ,
    \itasegm1[220] ,
    \itasegm1[219] ,
    \itasegm1[218] ,
    \itasegm1[217] ,
    \itasegm1[216] ,
    \itasegm1[215] ,
    \itasegm1[214] ,
    \itasegm1[213] ,
    \itasegm1[212] ,
    \itasegm1[211] ,
    \itasegm1[210] ,
    \itasegm1[209] ,
    \itasegm1[208] ,
    \itasegm1[207] ,
    \itasegm1[206] ,
    \itasegm1[205] ,
    \itasegm1[204] ,
    \itasegm1[203] ,
    \itasegm1[202] ,
    \itasegm1[201] ,
    \itasegm1[200] ,
    \itasegm1[199] ,
    \itasegm1[198] ,
    \itasegm1[197] ,
    \itasegm1[196] ,
    \itasegm1[195] ,
    \itasegm1[194] ,
    \itasegm1[193] ,
    \itasegm1[192] ,
    \itasegm1[191] ,
    \itasegm1[190] ,
    \itasegm1[189] ,
    \itasegm1[188] ,
    \itasegm1[187] ,
    \itasegm1[186] ,
    \itasegm1[185] ,
    \itasegm1[184] ,
    \itasegm1[183] ,
    \itasegm1[182] ,
    \itasegm1[181] ,
    \itasegm1[180] ,
    \itasegm1[179] ,
    \itasegm1[178] ,
    \itasegm1[177] ,
    \itasegm1[176] ,
    \itasegm1[175] ,
    \itasegm1[174] ,
    \itasegm1[173] ,
    \itasegm1[172] ,
    \itasegm1[171] ,
    \itasegm1[170] ,
    \itasegm1[169] ,
    \itasegm1[168] ,
    \itasegm1[167] ,
    \itasegm1[166] ,
    \itasegm1[165] ,
    \itasegm1[164] ,
    \itasegm1[163] ,
    \itasegm1[162] ,
    \itasegm1[161] ,
    \itasegm1[160] ,
    \itasegm1[159] ,
    \itasegm1[158] ,
    \itasegm1[157] ,
    \itasegm1[156] ,
    \itasegm1[155] ,
    \itasegm1[154] ,
    \itasegm1[153] ,
    \itasegm1[152] ,
    \itasegm1[151] ,
    \itasegm1[150] ,
    \itasegm1[149] ,
    \itasegm1[148] ,
    \itasegm1[147] ,
    \itasegm1[146] ,
    \itasegm1[145] ,
    \itasegm1[144] ,
    \itasegm1[143] ,
    \itasegm1[142] ,
    \itasegm1[141] ,
    \itasegm1[140] ,
    \itasegm1[139] ,
    \itasegm1[138] ,
    \itasegm1[137] ,
    \itasegm1[136] ,
    \itasegm1[135] ,
    \itasegm1[134] ,
    \itasegm1[133] ,
    \itasegm1[132] ,
    \itasegm1[131] ,
    \itasegm1[130] ,
    \itasegm1[129] ,
    \itasegm1[128] ,
    \itasegm1[127] ,
    \itasegm1[126] ,
    \itasegm1[125] ,
    \itasegm1[124] ,
    \itasegm1[123] ,
    \itasegm1[122] ,
    \itasegm1[121] ,
    \itasegm1[120] ,
    \itasegm1[119] ,
    \itasegm1[118] ,
    \itasegm1[117] ,
    \itasegm1[116] ,
    \itasegm1[115] ,
    \itasegm1[114] ,
    \itasegm1[113] ,
    \itasegm1[112] ,
    \itasegm1[111] ,
    \itasegm1[110] ,
    \itasegm1[109] ,
    \itasegm1[108] ,
    \itasegm1[107] ,
    \itasegm1[106] ,
    \itasegm1[105] ,
    \itasegm1[104] ,
    \itasegm1[103] ,
    \itasegm1[102] ,
    \itasegm1[101] ,
    \itasegm1[100] ,
    \itasegm1[99] ,
    \itasegm1[98] ,
    \itasegm1[97] ,
    \itasegm1[96] ,
    \itasegm1[95] ,
    \itasegm1[94] ,
    \itasegm1[93] ,
    \itasegm1[92] ,
    \itasegm1[91] ,
    \itasegm1[90] ,
    \itasegm1[89] ,
    \itasegm1[88] ,
    \itasegm1[87] ,
    \itasegm1[86] ,
    \itasegm1[85] ,
    \itasegm1[84] ,
    \itasegm1[83] ,
    \itasegm1[82] ,
    \itasegm1[81] ,
    \itasegm1[80] ,
    \itasegm1[79] ,
    \itasegm1[78] ,
    \itasegm1[77] ,
    \itasegm1[76] ,
    \itasegm1[75] ,
    \itasegm1[74] ,
    \itasegm1[73] ,
    \itasegm1[72] ,
    \itasegm1[71] ,
    \itasegm1[70] ,
    \itasegm1[69] ,
    \itasegm1[68] ,
    \itasegm1[67] ,
    \itasegm1[66] ,
    \itasegm1[65] ,
    \itasegm1[64] ,
    \itasegm1[63] ,
    \itasegm1[62] ,
    \itasegm1[61] ,
    \itasegm1[60] ,
    \itasegm1[59] ,
    \itasegm1[58] ,
    \itasegm1[57] ,
    \itasegm1[56] ,
    \itasegm1[55] ,
    \itasegm1[54] ,
    \itasegm1[53] ,
    \itasegm1[52] ,
    \itasegm1[51] ,
    \itasegm1[50] ,
    \itasegm1[49] ,
    \itasegm1[48] ,
    \itasegm1[47] ,
    \itasegm1[46] ,
    \itasegm1[45] ,
    \itasegm1[44] ,
    \itasegm1[43] ,
    \itasegm1[42] ,
    \itasegm1[41] ,
    \itasegm1[40] ,
    \itasegm1[39] ,
    \itasegm1[38] ,
    \itasegm1[37] ,
    \itasegm1[36] ,
    \itasegm1[35] ,
    \itasegm1[34] ,
    \itasegm1[33] ,
    \itasegm1[32] ,
    \itasegm1[31] ,
    \itasegm1[30] ,
    \itasegm1[29] ,
    \itasegm1[28] ,
    \itasegm1[27] ,
    \itasegm1[26] ,
    \itasegm1[25] ,
    \itasegm1[24] ,
    \itasegm1[23] ,
    \itasegm1[22] ,
    \itasegm1[21] ,
    \itasegm1[20] ,
    \itasegm1[19] ,
    \itasegm1[18] ,
    \itasegm1[17] ,
    \itasegm1[16] ,
    \itasegm1[15] ,
    \itasegm1[14] ,
    \itasegm1[13] ,
    \itasegm1[12] ,
    \itasegm1[11] ,
    \itasegm1[10] ,
    \itasegm1[9] ,
    \itasegm1[8] ,
    \itasegm1[7] ,
    \itasegm1[6] ,
    \itasegm1[5] ,
    \itasegm1[4] ,
    \itasegm1[3] ,
    \itasegm1[2] ,
    \itasegm1[1] ,
    \itasegm1[0] }),
    .itasel({\itasel1[767] ,
    \itasel1[766] ,
    \itasel1[765] ,
    \itasel1[764] ,
    \itasel1[763] ,
    \itasel1[762] ,
    \itasel1[761] ,
    \itasel1[760] ,
    \itasel1[759] ,
    \itasel1[758] ,
    \itasel1[757] ,
    \itasel1[756] ,
    \itasel1[755] ,
    \itasel1[754] ,
    \itasel1[753] ,
    \itasel1[752] ,
    \itasel1[751] ,
    \itasel1[750] ,
    \itasel1[749] ,
    \itasel1[748] ,
    \itasel1[747] ,
    \itasel1[746] ,
    \itasel1[745] ,
    \itasel1[744] ,
    \itasel1[743] ,
    \itasel1[742] ,
    \itasel1[741] ,
    \itasel1[740] ,
    \itasel1[739] ,
    \itasel1[738] ,
    \itasel1[737] ,
    \itasel1[736] ,
    \itasel1[735] ,
    \itasel1[734] ,
    \itasel1[733] ,
    \itasel1[732] ,
    \itasel1[731] ,
    \itasel1[730] ,
    \itasel1[729] ,
    \itasel1[728] ,
    \itasel1[727] ,
    \itasel1[726] ,
    \itasel1[725] ,
    \itasel1[724] ,
    \itasel1[723] ,
    \itasel1[722] ,
    \itasel1[721] ,
    \itasel1[720] ,
    \itasel1[719] ,
    \itasel1[718] ,
    \itasel1[717] ,
    \itasel1[716] ,
    \itasel1[715] ,
    \itasel1[714] ,
    \itasel1[713] ,
    \itasel1[712] ,
    \itasel1[711] ,
    \itasel1[710] ,
    \itasel1[709] ,
    \itasel1[708] ,
    \itasel1[707] ,
    \itasel1[706] ,
    \itasel1[705] ,
    \itasel1[704] ,
    \itasel1[703] ,
    \itasel1[702] ,
    \itasel1[701] ,
    \itasel1[700] ,
    \itasel1[699] ,
    \itasel1[698] ,
    \itasel1[697] ,
    \itasel1[696] ,
    \itasel1[695] ,
    \itasel1[694] ,
    \itasel1[693] ,
    \itasel1[692] ,
    \itasel1[691] ,
    \itasel1[690] ,
    \itasel1[689] ,
    \itasel1[688] ,
    \itasel1[687] ,
    \itasel1[686] ,
    \itasel1[685] ,
    \itasel1[684] ,
    \itasel1[683] ,
    \itasel1[682] ,
    \itasel1[681] ,
    \itasel1[680] ,
    \itasel1[679] ,
    \itasel1[678] ,
    \itasel1[677] ,
    \itasel1[676] ,
    \itasel1[675] ,
    \itasel1[674] ,
    \itasel1[673] ,
    \itasel1[672] ,
    \itasel1[671] ,
    \itasel1[670] ,
    \itasel1[669] ,
    \itasel1[668] ,
    \itasel1[667] ,
    \itasel1[666] ,
    \itasel1[665] ,
    \itasel1[664] ,
    \itasel1[663] ,
    \itasel1[662] ,
    \itasel1[661] ,
    \itasel1[660] ,
    \itasel1[659] ,
    \itasel1[658] ,
    \itasel1[657] ,
    \itasel1[656] ,
    \itasel1[655] ,
    \itasel1[654] ,
    \itasel1[653] ,
    \itasel1[652] ,
    \itasel1[651] ,
    \itasel1[650] ,
    \itasel1[649] ,
    \itasel1[648] ,
    \itasel1[647] ,
    \itasel1[646] ,
    \itasel1[645] ,
    \itasel1[644] ,
    \itasel1[643] ,
    \itasel1[642] ,
    \itasel1[641] ,
    \itasel1[640] ,
    \itasel1[639] ,
    \itasel1[638] ,
    \itasel1[637] ,
    \itasel1[636] ,
    \itasel1[635] ,
    \itasel1[634] ,
    \itasel1[633] ,
    \itasel1[632] ,
    \itasel1[631] ,
    \itasel1[630] ,
    \itasel1[629] ,
    \itasel1[628] ,
    \itasel1[627] ,
    \itasel1[626] ,
    \itasel1[625] ,
    \itasel1[624] ,
    \itasel1[623] ,
    \itasel1[622] ,
    \itasel1[621] ,
    \itasel1[620] ,
    \itasel1[619] ,
    \itasel1[618] ,
    \itasel1[617] ,
    \itasel1[616] ,
    \itasel1[615] ,
    \itasel1[614] ,
    \itasel1[613] ,
    \itasel1[612] ,
    \itasel1[611] ,
    \itasel1[610] ,
    \itasel1[609] ,
    \itasel1[608] ,
    \itasel1[607] ,
    \itasel1[606] ,
    \itasel1[605] ,
    \itasel1[604] ,
    \itasel1[603] ,
    \itasel1[602] ,
    \itasel1[601] ,
    \itasel1[600] ,
    \itasel1[599] ,
    \itasel1[598] ,
    \itasel1[597] ,
    \itasel1[596] ,
    \itasel1[595] ,
    \itasel1[594] ,
    \itasel1[593] ,
    \itasel1[592] ,
    \itasel1[591] ,
    \itasel1[590] ,
    \itasel1[589] ,
    \itasel1[588] ,
    \itasel1[587] ,
    \itasel1[586] ,
    \itasel1[585] ,
    \itasel1[584] ,
    \itasel1[583] ,
    \itasel1[582] ,
    \itasel1[581] ,
    \itasel1[580] ,
    \itasel1[579] ,
    \itasel1[578] ,
    \itasel1[577] ,
    \itasel1[576] ,
    \itasel1[575] ,
    \itasel1[574] ,
    \itasel1[573] ,
    \itasel1[572] ,
    \itasel1[571] ,
    \itasel1[570] ,
    \itasel1[569] ,
    \itasel1[568] ,
    \itasel1[567] ,
    \itasel1[566] ,
    \itasel1[565] ,
    \itasel1[564] ,
    \itasel1[563] ,
    \itasel1[562] ,
    \itasel1[561] ,
    \itasel1[560] ,
    \itasel1[559] ,
    \itasel1[558] ,
    \itasel1[557] ,
    \itasel1[556] ,
    \itasel1[555] ,
    \itasel1[554] ,
    \itasel1[553] ,
    \itasel1[552] ,
    \itasel1[551] ,
    \itasel1[550] ,
    \itasel1[549] ,
    \itasel1[548] ,
    \itasel1[547] ,
    \itasel1[546] ,
    \itasel1[545] ,
    \itasel1[544] ,
    \itasel1[543] ,
    \itasel1[542] ,
    \itasel1[541] ,
    \itasel1[540] ,
    \itasel1[539] ,
    \itasel1[538] ,
    \itasel1[537] ,
    \itasel1[536] ,
    \itasel1[535] ,
    \itasel1[534] ,
    \itasel1[533] ,
    \itasel1[532] ,
    \itasel1[531] ,
    \itasel1[530] ,
    \itasel1[529] ,
    \itasel1[528] ,
    \itasel1[527] ,
    \itasel1[526] ,
    \itasel1[525] ,
    \itasel1[524] ,
    \itasel1[523] ,
    \itasel1[522] ,
    \itasel1[521] ,
    \itasel1[520] ,
    \itasel1[519] ,
    \itasel1[518] ,
    \itasel1[517] ,
    \itasel1[516] ,
    \itasel1[515] ,
    \itasel1[514] ,
    \itasel1[513] ,
    \itasel1[512] ,
    \itasel1[511] ,
    \itasel1[510] ,
    \itasel1[509] ,
    \itasel1[508] ,
    \itasel1[507] ,
    \itasel1[506] ,
    \itasel1[505] ,
    \itasel1[504] ,
    \itasel1[503] ,
    \itasel1[502] ,
    \itasel1[501] ,
    \itasel1[500] ,
    \itasel1[499] ,
    \itasel1[498] ,
    \itasel1[497] ,
    \itasel1[496] ,
    \itasel1[495] ,
    \itasel1[494] ,
    \itasel1[493] ,
    \itasel1[492] ,
    \itasel1[491] ,
    \itasel1[490] ,
    \itasel1[489] ,
    \itasel1[488] ,
    \itasel1[487] ,
    \itasel1[486] ,
    \itasel1[485] ,
    \itasel1[484] ,
    \itasel1[483] ,
    \itasel1[482] ,
    \itasel1[481] ,
    \itasel1[480] ,
    \itasel1[479] ,
    \itasel1[478] ,
    \itasel1[477] ,
    \itasel1[476] ,
    \itasel1[475] ,
    \itasel1[474] ,
    \itasel1[473] ,
    \itasel1[472] ,
    \itasel1[471] ,
    \itasel1[470] ,
    \itasel1[469] ,
    \itasel1[468] ,
    \itasel1[467] ,
    \itasel1[466] ,
    \itasel1[465] ,
    \itasel1[464] ,
    \itasel1[463] ,
    \itasel1[462] ,
    \itasel1[461] ,
    \itasel1[460] ,
    \itasel1[459] ,
    \itasel1[458] ,
    \itasel1[457] ,
    \itasel1[456] ,
    \itasel1[455] ,
    \itasel1[454] ,
    \itasel1[453] ,
    \itasel1[452] ,
    \itasel1[451] ,
    \itasel1[450] ,
    \itasel1[449] ,
    \itasel1[448] ,
    \itasel1[447] ,
    \itasel1[446] ,
    \itasel1[445] ,
    \itasel1[444] ,
    \itasel1[443] ,
    \itasel1[442] ,
    \itasel1[441] ,
    \itasel1[440] ,
    \itasel1[439] ,
    \itasel1[438] ,
    \itasel1[437] ,
    \itasel1[436] ,
    \itasel1[435] ,
    \itasel1[434] ,
    \itasel1[433] ,
    \itasel1[432] ,
    \itasel1[431] ,
    \itasel1[430] ,
    \itasel1[429] ,
    \itasel1[428] ,
    \itasel1[427] ,
    \itasel1[426] ,
    \itasel1[425] ,
    \itasel1[424] ,
    \itasel1[423] ,
    \itasel1[422] ,
    \itasel1[421] ,
    \itasel1[420] ,
    \itasel1[419] ,
    \itasel1[418] ,
    \itasel1[417] ,
    \itasel1[416] ,
    \itasel1[415] ,
    \itasel1[414] ,
    \itasel1[413] ,
    \itasel1[412] ,
    \itasel1[411] ,
    \itasel1[410] ,
    \itasel1[409] ,
    \itasel1[408] ,
    \itasel1[407] ,
    \itasel1[406] ,
    \itasel1[405] ,
    \itasel1[404] ,
    \itasel1[403] ,
    \itasel1[402] ,
    \itasel1[401] ,
    \itasel1[400] ,
    \itasel1[399] ,
    \itasel1[398] ,
    \itasel1[397] ,
    \itasel1[396] ,
    \itasel1[395] ,
    \itasel1[394] ,
    \itasel1[393] ,
    \itasel1[392] ,
    \itasel1[391] ,
    \itasel1[390] ,
    \itasel1[389] ,
    \itasel1[388] ,
    \itasel1[387] ,
    \itasel1[386] ,
    \itasel1[385] ,
    \itasel1[384] ,
    \itasel1[383] ,
    \itasel1[382] ,
    \itasel1[381] ,
    \itasel1[380] ,
    \itasel1[379] ,
    \itasel1[378] ,
    \itasel1[377] ,
    \itasel1[376] ,
    \itasel1[375] ,
    \itasel1[374] ,
    \itasel1[373] ,
    \itasel1[372] ,
    \itasel1[371] ,
    \itasel1[370] ,
    \itasel1[369] ,
    \itasel1[368] ,
    \itasel1[367] ,
    \itasel1[366] ,
    \itasel1[365] ,
    \itasel1[364] ,
    \itasel1[363] ,
    \itasel1[362] ,
    \itasel1[361] ,
    \itasel1[360] ,
    \itasel1[359] ,
    \itasel1[358] ,
    \itasel1[357] ,
    \itasel1[356] ,
    \itasel1[355] ,
    \itasel1[354] ,
    \itasel1[353] ,
    \itasel1[352] ,
    \itasel1[351] ,
    \itasel1[350] ,
    \itasel1[349] ,
    \itasel1[348] ,
    \itasel1[347] ,
    \itasel1[346] ,
    \itasel1[345] ,
    \itasel1[344] ,
    \itasel1[343] ,
    \itasel1[342] ,
    \itasel1[341] ,
    \itasel1[340] ,
    \itasel1[339] ,
    \itasel1[338] ,
    \itasel1[337] ,
    \itasel1[336] ,
    \itasel1[335] ,
    \itasel1[334] ,
    \itasel1[333] ,
    \itasel1[332] ,
    \itasel1[331] ,
    \itasel1[330] ,
    \itasel1[329] ,
    \itasel1[328] ,
    \itasel1[327] ,
    \itasel1[326] ,
    \itasel1[325] ,
    \itasel1[324] ,
    \itasel1[323] ,
    \itasel1[322] ,
    \itasel1[321] ,
    \itasel1[320] ,
    \itasel1[319] ,
    \itasel1[318] ,
    \itasel1[317] ,
    \itasel1[316] ,
    \itasel1[315] ,
    \itasel1[314] ,
    \itasel1[313] ,
    \itasel1[312] ,
    \itasel1[311] ,
    \itasel1[310] ,
    \itasel1[309] ,
    \itasel1[308] ,
    \itasel1[307] ,
    \itasel1[306] ,
    \itasel1[305] ,
    \itasel1[304] ,
    \itasel1[303] ,
    \itasel1[302] ,
    \itasel1[301] ,
    \itasel1[300] ,
    \itasel1[299] ,
    \itasel1[298] ,
    \itasel1[297] ,
    \itasel1[296] ,
    \itasel1[295] ,
    \itasel1[294] ,
    \itasel1[293] ,
    \itasel1[292] ,
    \itasel1[291] ,
    \itasel1[290] ,
    \itasel1[289] ,
    \itasel1[288] ,
    \itasel1[287] ,
    \itasel1[286] ,
    \itasel1[285] ,
    \itasel1[284] ,
    \itasel1[283] ,
    \itasel1[282] ,
    \itasel1[281] ,
    \itasel1[280] ,
    \itasel1[279] ,
    \itasel1[278] ,
    \itasel1[277] ,
    \itasel1[276] ,
    \itasel1[275] ,
    \itasel1[274] ,
    \itasel1[273] ,
    \itasel1[272] ,
    \itasel1[271] ,
    \itasel1[270] ,
    \itasel1[269] ,
    \itasel1[268] ,
    \itasel1[267] ,
    \itasel1[266] ,
    \itasel1[265] ,
    \itasel1[264] ,
    \itasel1[263] ,
    \itasel1[262] ,
    \itasel1[261] ,
    \itasel1[260] ,
    \itasel1[259] ,
    \itasel1[258] ,
    \itasel1[257] ,
    \itasel1[256] ,
    \itasel1[255] ,
    \itasel1[254] ,
    \itasel1[253] ,
    \itasel1[252] ,
    \itasel1[251] ,
    \itasel1[250] ,
    \itasel1[249] ,
    \itasel1[248] ,
    \itasel1[247] ,
    \itasel1[246] ,
    \itasel1[245] ,
    \itasel1[244] ,
    \itasel1[243] ,
    \itasel1[242] ,
    \itasel1[241] ,
    \itasel1[240] ,
    \itasel1[239] ,
    \itasel1[238] ,
    \itasel1[237] ,
    \itasel1[236] ,
    \itasel1[235] ,
    \itasel1[234] ,
    \itasel1[233] ,
    \itasel1[232] ,
    \itasel1[231] ,
    \itasel1[230] ,
    \itasel1[229] ,
    \itasel1[228] ,
    \itasel1[227] ,
    \itasel1[226] ,
    \itasel1[225] ,
    \itasel1[224] ,
    \itasel1[223] ,
    \itasel1[222] ,
    \itasel1[221] ,
    \itasel1[220] ,
    \itasel1[219] ,
    \itasel1[218] ,
    \itasel1[217] ,
    \itasel1[216] ,
    \itasel1[215] ,
    \itasel1[214] ,
    \itasel1[213] ,
    \itasel1[212] ,
    \itasel1[211] ,
    \itasel1[210] ,
    \itasel1[209] ,
    \itasel1[208] ,
    \itasel1[207] ,
    \itasel1[206] ,
    \itasel1[205] ,
    \itasel1[204] ,
    \itasel1[203] ,
    \itasel1[202] ,
    \itasel1[201] ,
    \itasel1[200] ,
    \itasel1[199] ,
    \itasel1[198] ,
    \itasel1[197] ,
    \itasel1[196] ,
    \itasel1[195] ,
    \itasel1[194] ,
    \itasel1[193] ,
    \itasel1[192] ,
    \itasel1[191] ,
    \itasel1[190] ,
    \itasel1[189] ,
    \itasel1[188] ,
    \itasel1[187] ,
    \itasel1[186] ,
    \itasel1[185] ,
    \itasel1[184] ,
    \itasel1[183] ,
    \itasel1[182] ,
    \itasel1[181] ,
    \itasel1[180] ,
    \itasel1[179] ,
    \itasel1[178] ,
    \itasel1[177] ,
    \itasel1[176] ,
    \itasel1[175] ,
    \itasel1[174] ,
    \itasel1[173] ,
    \itasel1[172] ,
    \itasel1[171] ,
    \itasel1[170] ,
    \itasel1[169] ,
    \itasel1[168] ,
    \itasel1[167] ,
    \itasel1[166] ,
    \itasel1[165] ,
    \itasel1[164] ,
    \itasel1[163] ,
    \itasel1[162] ,
    \itasel1[161] ,
    \itasel1[160] ,
    \itasel1[159] ,
    \itasel1[158] ,
    \itasel1[157] ,
    \itasel1[156] ,
    \itasel1[155] ,
    \itasel1[154] ,
    \itasel1[153] ,
    \itasel1[152] ,
    \itasel1[151] ,
    \itasel1[150] ,
    \itasel1[149] ,
    \itasel1[148] ,
    \itasel1[147] ,
    \itasel1[146] ,
    \itasel1[145] ,
    \itasel1[144] ,
    \itasel1[143] ,
    \itasel1[142] ,
    \itasel1[141] ,
    \itasel1[140] ,
    \itasel1[139] ,
    \itasel1[138] ,
    \itasel1[137] ,
    \itasel1[136] ,
    \itasel1[135] ,
    \itasel1[134] ,
    \itasel1[133] ,
    \itasel1[132] ,
    \itasel1[131] ,
    \itasel1[130] ,
    \itasel1[129] ,
    \itasel1[128] ,
    \itasel1[127] ,
    \itasel1[126] ,
    \itasel1[125] ,
    \itasel1[124] ,
    \itasel1[123] ,
    \itasel1[122] ,
    \itasel1[121] ,
    \itasel1[120] ,
    \itasel1[119] ,
    \itasel1[118] ,
    \itasel1[117] ,
    \itasel1[116] ,
    \itasel1[115] ,
    \itasel1[114] ,
    \itasel1[113] ,
    \itasel1[112] ,
    \itasel1[111] ,
    \itasel1[110] ,
    \itasel1[109] ,
    \itasel1[108] ,
    \itasel1[107] ,
    \itasel1[106] ,
    \itasel1[105] ,
    \itasel1[104] ,
    \itasel1[103] ,
    \itasel1[102] ,
    \itasel1[101] ,
    \itasel1[100] ,
    \itasel1[99] ,
    \itasel1[98] ,
    \itasel1[97] ,
    \itasel1[96] ,
    \itasel1[95] ,
    \itasel1[94] ,
    \itasel1[93] ,
    \itasel1[92] ,
    \itasel1[91] ,
    \itasel1[90] ,
    \itasel1[89] ,
    \itasel1[88] ,
    \itasel1[87] ,
    \itasel1[86] ,
    \itasel1[85] ,
    \itasel1[84] ,
    \itasel1[83] ,
    \itasel1[82] ,
    \itasel1[81] ,
    \itasel1[80] ,
    \itasel1[79] ,
    \itasel1[78] ,
    \itasel1[77] ,
    \itasel1[76] ,
    \itasel1[75] ,
    \itasel1[74] ,
    \itasel1[73] ,
    \itasel1[72] ,
    \itasel1[71] ,
    \itasel1[70] ,
    \itasel1[69] ,
    \itasel1[68] ,
    \itasel1[67] ,
    \itasel1[66] ,
    \itasel1[65] ,
    \itasel1[64] ,
    \itasel1[63] ,
    \itasel1[62] ,
    \itasel1[61] ,
    \itasel1[60] ,
    \itasel1[59] ,
    \itasel1[58] ,
    \itasel1[57] ,
    \itasel1[56] ,
    \itasel1[55] ,
    \itasel1[54] ,
    \itasel1[53] ,
    \itasel1[52] ,
    \itasel1[51] ,
    \itasel1[50] ,
    \itasel1[49] ,
    \itasel1[48] ,
    \itasel1[47] ,
    \itasel1[46] ,
    \itasel1[45] ,
    \itasel1[44] ,
    \itasel1[43] ,
    \itasel1[42] ,
    \itasel1[41] ,
    \itasel1[40] ,
    \itasel1[39] ,
    \itasel1[38] ,
    \itasel1[37] ,
    \itasel1[36] ,
    \itasel1[35] ,
    \itasel1[34] ,
    \itasel1[33] ,
    \itasel1[32] ,
    \itasel1[31] ,
    \itasel1[30] ,
    \itasel1[29] ,
    \itasel1[28] ,
    \itasel1[27] ,
    \itasel1[26] ,
    \itasel1[25] ,
    \itasel1[24] ,
    \itasel1[23] ,
    \itasel1[22] ,
    \itasel1[21] ,
    \itasel1[20] ,
    \itasel1[19] ,
    \itasel1[18] ,
    \itasel1[17] ,
    \itasel1[16] ,
    \itasel1[15] ,
    \itasel1[14] ,
    \itasel1[13] ,
    \itasel1[12] ,
    \itasel1[11] ,
    \itasel1[10] ,
    \itasel1[9] ,
    \itasel1[8] ,
    \itasel1[7] ,
    \itasel1[6] ,
    \itasel1[5] ,
    \itasel1[4] ,
    \itasel1[3] ,
    \itasel1[2] ,
    \itasel1[1] ,
    \itasel1[0] }),
    .nsel({io_in[11],
    io_in[10],
    io_in[9],
    io_in[8],
    io_in[7],
    io_in[6]}),
    .segm({io_out[37],
    io_out[36],
    io_out[35],
    io_out[34],
    io_out[33],
    io_out[32],
    io_out[31],
    io_out[30],
    io_out[29],
    io_out[28],
    io_out[27],
    io_out[26],
    io_out[25],
    io_out[24]}),
    .sel({io_out[23],
    io_out[22],
    io_out[21],
    io_out[20],
    io_out[19],
    io_out[18],
    io_out[17],
    io_out[16],
    io_out[15],
    io_out[14],
    io_out[13],
    io_out[12]}));
 ita1 ita1 (.clk(wb_clk_i),
    .segm({\itasegm1[13] ,
    \itasegm1[12] ,
    \itasegm1[11] ,
    \itasegm1[10] ,
    \itasegm1[9] ,
    \itasegm1[8] ,
    \itasegm1[7] ,
    \itasegm1[6] ,
    \itasegm1[5] ,
    \itasegm1[4] ,
    \itasegm1[3] ,
    \itasegm1[2] ,
    \itasegm1[1] ,
    \itasegm1[0] }),
    .sel({\itasel1[11] ,
    \itasel1[10] ,
    \itasel1[9] ,
    \itasel1[8] ,
    \itasel1[7] ,
    \itasel1[6] ,
    \itasel1[5] ,
    \itasel1[4] ,
    \itasel1[3] ,
    \itasel1[2] ,
    \itasel1[1] ,
    \itasel1[0] }));
 ita10 ita10 (.clk(wb_clk_i),
    .segm({\itasegm1[139] ,
    \itasegm1[138] ,
    \itasegm1[137] ,
    \itasegm1[136] ,
    \itasegm1[135] ,
    \itasegm1[134] ,
    \itasegm1[133] ,
    \itasegm1[132] ,
    \itasegm1[131] ,
    \itasegm1[130] ,
    \itasegm1[129] ,
    \itasegm1[128] ,
    \itasegm1[127] ,
    \itasegm1[126] }),
    .sel({\itasel1[119] ,
    \itasel1[118] ,
    \itasel1[117] ,
    \itasel1[116] ,
    \itasel1[115] ,
    \itasel1[114] ,
    \itasel1[113] ,
    \itasel1[112] ,
    \itasel1[111] ,
    \itasel1[110] ,
    \itasel1[109] ,
    \itasel1[108] }));
 ita11 ita11 (.clk(wb_clk_i),
    .segm({\itasegm1[153] ,
    \itasegm1[152] ,
    \itasegm1[151] ,
    \itasegm1[150] ,
    \itasegm1[149] ,
    \itasegm1[148] ,
    \itasegm1[147] ,
    \itasegm1[146] ,
    \itasegm1[145] ,
    \itasegm1[144] ,
    \itasegm1[143] ,
    \itasegm1[142] ,
    \itasegm1[141] ,
    \itasegm1[140] }),
    .sel({\itasel1[131] ,
    \itasel1[130] ,
    \itasel1[129] ,
    \itasel1[128] ,
    \itasel1[127] ,
    \itasel1[126] ,
    \itasel1[125] ,
    \itasel1[124] ,
    \itasel1[123] ,
    \itasel1[122] ,
    \itasel1[121] ,
    \itasel1[120] }));
 ita12 ita12 (.clk(wb_clk_i),
    .segm({\itasegm1[167] ,
    \itasegm1[166] ,
    \itasegm1[165] ,
    \itasegm1[164] ,
    \itasegm1[163] ,
    \itasegm1[162] ,
    \itasegm1[161] ,
    \itasegm1[160] ,
    \itasegm1[159] ,
    \itasegm1[158] ,
    \itasegm1[157] ,
    \itasegm1[156] ,
    \itasegm1[155] ,
    \itasegm1[154] }),
    .sel({\itasel1[143] ,
    \itasel1[142] ,
    \itasel1[141] ,
    \itasel1[140] ,
    \itasel1[139] ,
    \itasel1[138] ,
    \itasel1[137] ,
    \itasel1[136] ,
    \itasel1[135] ,
    \itasel1[134] ,
    \itasel1[133] ,
    \itasel1[132] }));
 ita13 ita13 (.clk(wb_clk_i),
    .segm({\itasegm1[181] ,
    \itasegm1[180] ,
    \itasegm1[179] ,
    \itasegm1[178] ,
    \itasegm1[177] ,
    \itasegm1[176] ,
    \itasegm1[175] ,
    \itasegm1[174] ,
    \itasegm1[173] ,
    \itasegm1[172] ,
    \itasegm1[171] ,
    \itasegm1[170] ,
    \itasegm1[169] ,
    \itasegm1[168] }),
    .sel({\itasel1[155] ,
    \itasel1[154] ,
    \itasel1[153] ,
    \itasel1[152] ,
    \itasel1[151] ,
    \itasel1[150] ,
    \itasel1[149] ,
    \itasel1[148] ,
    \itasel1[147] ,
    \itasel1[146] ,
    \itasel1[145] ,
    \itasel1[144] }));
 ita14 ita14 (.clk(wb_clk_i),
    .segm({\itasegm1[195] ,
    \itasegm1[194] ,
    \itasegm1[193] ,
    \itasegm1[192] ,
    \itasegm1[191] ,
    \itasegm1[190] ,
    \itasegm1[189] ,
    \itasegm1[188] ,
    \itasegm1[187] ,
    \itasegm1[186] ,
    \itasegm1[185] ,
    \itasegm1[184] ,
    \itasegm1[183] ,
    \itasegm1[182] }),
    .sel({\itasel1[167] ,
    \itasel1[166] ,
    \itasel1[165] ,
    \itasel1[164] ,
    \itasel1[163] ,
    \itasel1[162] ,
    \itasel1[161] ,
    \itasel1[160] ,
    \itasel1[159] ,
    \itasel1[158] ,
    \itasel1[157] ,
    \itasel1[156] }));
 ita15 ita15 (.clk(wb_clk_i),
    .segm({\itasegm1[209] ,
    \itasegm1[208] ,
    \itasegm1[207] ,
    \itasegm1[206] ,
    \itasegm1[205] ,
    \itasegm1[204] ,
    \itasegm1[203] ,
    \itasegm1[202] ,
    \itasegm1[201] ,
    \itasegm1[200] ,
    \itasegm1[199] ,
    \itasegm1[198] ,
    \itasegm1[197] ,
    \itasegm1[196] }),
    .sel({\itasel1[179] ,
    \itasel1[178] ,
    \itasel1[177] ,
    \itasel1[176] ,
    \itasel1[175] ,
    \itasel1[174] ,
    \itasel1[173] ,
    \itasel1[172] ,
    \itasel1[171] ,
    \itasel1[170] ,
    \itasel1[169] ,
    \itasel1[168] }));
 ita16 ita16 (.clk(wb_clk_i),
    .segm({\itasegm1[223] ,
    \itasegm1[222] ,
    \itasegm1[221] ,
    \itasegm1[220] ,
    \itasegm1[219] ,
    \itasegm1[218] ,
    \itasegm1[217] ,
    \itasegm1[216] ,
    \itasegm1[215] ,
    \itasegm1[214] ,
    \itasegm1[213] ,
    \itasegm1[212] ,
    \itasegm1[211] ,
    \itasegm1[210] }),
    .sel({\itasel1[191] ,
    \itasel1[190] ,
    \itasel1[189] ,
    \itasel1[188] ,
    \itasel1[187] ,
    \itasel1[186] ,
    \itasel1[185] ,
    \itasel1[184] ,
    \itasel1[183] ,
    \itasel1[182] ,
    \itasel1[181] ,
    \itasel1[180] }));
 ita17 ita17 (.clk(wb_clk_i),
    .segm({\itasegm1[237] ,
    \itasegm1[236] ,
    \itasegm1[235] ,
    \itasegm1[234] ,
    \itasegm1[233] ,
    \itasegm1[232] ,
    \itasegm1[231] ,
    \itasegm1[230] ,
    \itasegm1[229] ,
    \itasegm1[228] ,
    \itasegm1[227] ,
    \itasegm1[226] ,
    \itasegm1[225] ,
    \itasegm1[224] }),
    .sel({\itasel1[203] ,
    \itasel1[202] ,
    \itasel1[201] ,
    \itasel1[200] ,
    \itasel1[199] ,
    \itasel1[198] ,
    \itasel1[197] ,
    \itasel1[196] ,
    \itasel1[195] ,
    \itasel1[194] ,
    \itasel1[193] ,
    \itasel1[192] }));
 ita18 ita18 (.clk(wb_clk_i),
    .segm({\itasegm1[251] ,
    \itasegm1[250] ,
    \itasegm1[249] ,
    \itasegm1[248] ,
    \itasegm1[247] ,
    \itasegm1[246] ,
    \itasegm1[245] ,
    \itasegm1[244] ,
    \itasegm1[243] ,
    \itasegm1[242] ,
    \itasegm1[241] ,
    \itasegm1[240] ,
    \itasegm1[239] ,
    \itasegm1[238] }),
    .sel({\itasel1[215] ,
    \itasel1[214] ,
    \itasel1[213] ,
    \itasel1[212] ,
    \itasel1[211] ,
    \itasel1[210] ,
    \itasel1[209] ,
    \itasel1[208] ,
    \itasel1[207] ,
    \itasel1[206] ,
    \itasel1[205] ,
    \itasel1[204] }));
 ita19 ita19 (.clk(wb_clk_i),
    .segm({\itasegm1[265] ,
    \itasegm1[264] ,
    \itasegm1[263] ,
    \itasegm1[262] ,
    \itasegm1[261] ,
    \itasegm1[260] ,
    \itasegm1[259] ,
    \itasegm1[258] ,
    \itasegm1[257] ,
    \itasegm1[256] ,
    \itasegm1[255] ,
    \itasegm1[254] ,
    \itasegm1[253] ,
    \itasegm1[252] }),
    .sel({\itasel1[227] ,
    \itasel1[226] ,
    \itasel1[225] ,
    \itasel1[224] ,
    \itasel1[223] ,
    \itasel1[222] ,
    \itasel1[221] ,
    \itasel1[220] ,
    \itasel1[219] ,
    \itasel1[218] ,
    \itasel1[217] ,
    \itasel1[216] }));
 ita2 ita2 (.clk(wb_clk_i),
    .segm({\itasegm1[27] ,
    \itasegm1[26] ,
    \itasegm1[25] ,
    \itasegm1[24] ,
    \itasegm1[23] ,
    \itasegm1[22] ,
    \itasegm1[21] ,
    \itasegm1[20] ,
    \itasegm1[19] ,
    \itasegm1[18] ,
    \itasegm1[17] ,
    \itasegm1[16] ,
    \itasegm1[15] ,
    \itasegm1[14] }),
    .sel({\itasel1[23] ,
    \itasel1[22] ,
    \itasel1[21] ,
    \itasel1[20] ,
    \itasel1[19] ,
    \itasel1[18] ,
    \itasel1[17] ,
    \itasel1[16] ,
    \itasel1[15] ,
    \itasel1[14] ,
    \itasel1[13] ,
    \itasel1[12] }));
 ita20 ita20 (.clk(wb_clk_i),
    .segm({\itasegm1[279] ,
    \itasegm1[278] ,
    \itasegm1[277] ,
    \itasegm1[276] ,
    \itasegm1[275] ,
    \itasegm1[274] ,
    \itasegm1[273] ,
    \itasegm1[272] ,
    \itasegm1[271] ,
    \itasegm1[270] ,
    \itasegm1[269] ,
    \itasegm1[268] ,
    \itasegm1[267] ,
    \itasegm1[266] }),
    .sel({\itasel1[239] ,
    \itasel1[238] ,
    \itasel1[237] ,
    \itasel1[236] ,
    \itasel1[235] ,
    \itasel1[234] ,
    \itasel1[233] ,
    \itasel1[232] ,
    \itasel1[231] ,
    \itasel1[230] ,
    \itasel1[229] ,
    \itasel1[228] }));
 ita21 ita21 (.clk(wb_clk_i),
    .segm({\itasegm1[293] ,
    \itasegm1[292] ,
    \itasegm1[291] ,
    \itasegm1[290] ,
    \itasegm1[289] ,
    \itasegm1[288] ,
    \itasegm1[287] ,
    \itasegm1[286] ,
    \itasegm1[285] ,
    \itasegm1[284] ,
    \itasegm1[283] ,
    \itasegm1[282] ,
    \itasegm1[281] ,
    \itasegm1[280] }),
    .sel({\itasel1[251] ,
    \itasel1[250] ,
    \itasel1[249] ,
    \itasel1[248] ,
    \itasel1[247] ,
    \itasel1[246] ,
    \itasel1[245] ,
    \itasel1[244] ,
    \itasel1[243] ,
    \itasel1[242] ,
    \itasel1[241] ,
    \itasel1[240] }));
 ita22 ita22 (.clk(wb_clk_i),
    .segm({\itasegm1[307] ,
    \itasegm1[306] ,
    \itasegm1[305] ,
    \itasegm1[304] ,
    \itasegm1[303] ,
    \itasegm1[302] ,
    \itasegm1[301] ,
    \itasegm1[300] ,
    \itasegm1[299] ,
    \itasegm1[298] ,
    \itasegm1[297] ,
    \itasegm1[296] ,
    \itasegm1[295] ,
    \itasegm1[294] }),
    .sel({\itasel1[263] ,
    \itasel1[262] ,
    \itasel1[261] ,
    \itasel1[260] ,
    \itasel1[259] ,
    \itasel1[258] ,
    \itasel1[257] ,
    \itasel1[256] ,
    \itasel1[255] ,
    \itasel1[254] ,
    \itasel1[253] ,
    \itasel1[252] }));
 ita23 ita23 (.clk(wb_clk_i),
    .segm({\itasegm1[321] ,
    \itasegm1[320] ,
    \itasegm1[319] ,
    \itasegm1[318] ,
    \itasegm1[317] ,
    \itasegm1[316] ,
    \itasegm1[315] ,
    \itasegm1[314] ,
    \itasegm1[313] ,
    \itasegm1[312] ,
    \itasegm1[311] ,
    \itasegm1[310] ,
    \itasegm1[309] ,
    \itasegm1[308] }),
    .sel({\itasel1[275] ,
    \itasel1[274] ,
    \itasel1[273] ,
    \itasel1[272] ,
    \itasel1[271] ,
    \itasel1[270] ,
    \itasel1[269] ,
    \itasel1[268] ,
    \itasel1[267] ,
    \itasel1[266] ,
    \itasel1[265] ,
    \itasel1[264] }));
 ita24 ita24 (.clk(wb_clk_i),
    .segm({\itasegm1[335] ,
    \itasegm1[334] ,
    \itasegm1[333] ,
    \itasegm1[332] ,
    \itasegm1[331] ,
    \itasegm1[330] ,
    \itasegm1[329] ,
    \itasegm1[328] ,
    \itasegm1[327] ,
    \itasegm1[326] ,
    \itasegm1[325] ,
    \itasegm1[324] ,
    \itasegm1[323] ,
    \itasegm1[322] }),
    .sel({\itasel1[287] ,
    \itasel1[286] ,
    \itasel1[285] ,
    \itasel1[284] ,
    \itasel1[283] ,
    \itasel1[282] ,
    \itasel1[281] ,
    \itasel1[280] ,
    \itasel1[279] ,
    \itasel1[278] ,
    \itasel1[277] ,
    \itasel1[276] }));
 ita25 ita25 (.clk(wb_clk_i),
    .segm({\itasegm1[349] ,
    \itasegm1[348] ,
    \itasegm1[347] ,
    \itasegm1[346] ,
    \itasegm1[345] ,
    \itasegm1[344] ,
    \itasegm1[343] ,
    \itasegm1[342] ,
    \itasegm1[341] ,
    \itasegm1[340] ,
    \itasegm1[339] ,
    \itasegm1[338] ,
    \itasegm1[337] ,
    \itasegm1[336] }),
    .sel({\itasel1[299] ,
    \itasel1[298] ,
    \itasel1[297] ,
    \itasel1[296] ,
    \itasel1[295] ,
    \itasel1[294] ,
    \itasel1[293] ,
    \itasel1[292] ,
    \itasel1[291] ,
    \itasel1[290] ,
    \itasel1[289] ,
    \itasel1[288] }));
 ita26 ita26 (.clk(wb_clk_i),
    .segm({\itasegm1[363] ,
    \itasegm1[362] ,
    \itasegm1[361] ,
    \itasegm1[360] ,
    \itasegm1[359] ,
    \itasegm1[358] ,
    \itasegm1[357] ,
    \itasegm1[356] ,
    \itasegm1[355] ,
    \itasegm1[354] ,
    \itasegm1[353] ,
    \itasegm1[352] ,
    \itasegm1[351] ,
    \itasegm1[350] }),
    .sel({\itasel1[311] ,
    \itasel1[310] ,
    \itasel1[309] ,
    \itasel1[308] ,
    \itasel1[307] ,
    \itasel1[306] ,
    \itasel1[305] ,
    \itasel1[304] ,
    \itasel1[303] ,
    \itasel1[302] ,
    \itasel1[301] ,
    \itasel1[300] }));
 ita27 ita27 (.clk(wb_clk_i),
    .segm({\itasegm1[377] ,
    \itasegm1[376] ,
    \itasegm1[375] ,
    \itasegm1[374] ,
    \itasegm1[373] ,
    \itasegm1[372] ,
    \itasegm1[371] ,
    \itasegm1[370] ,
    \itasegm1[369] ,
    \itasegm1[368] ,
    \itasegm1[367] ,
    \itasegm1[366] ,
    \itasegm1[365] ,
    \itasegm1[364] }),
    .sel({\itasel1[323] ,
    \itasel1[322] ,
    \itasel1[321] ,
    \itasel1[320] ,
    \itasel1[319] ,
    \itasel1[318] ,
    \itasel1[317] ,
    \itasel1[316] ,
    \itasel1[315] ,
    \itasel1[314] ,
    \itasel1[313] ,
    \itasel1[312] }));
 ita28 ita28 (.clk(wb_clk_i),
    .segm({\itasegm1[391] ,
    \itasegm1[390] ,
    \itasegm1[389] ,
    \itasegm1[388] ,
    \itasegm1[387] ,
    \itasegm1[386] ,
    \itasegm1[385] ,
    \itasegm1[384] ,
    \itasegm1[383] ,
    \itasegm1[382] ,
    \itasegm1[381] ,
    \itasegm1[380] ,
    \itasegm1[379] ,
    \itasegm1[378] }),
    .sel({\itasel1[335] ,
    \itasel1[334] ,
    \itasel1[333] ,
    \itasel1[332] ,
    \itasel1[331] ,
    \itasel1[330] ,
    \itasel1[329] ,
    \itasel1[328] ,
    \itasel1[327] ,
    \itasel1[326] ,
    \itasel1[325] ,
    \itasel1[324] }));
 ita29 ita29 (.clk(wb_clk_i),
    .segm({\itasegm1[405] ,
    \itasegm1[404] ,
    \itasegm1[403] ,
    \itasegm1[402] ,
    \itasegm1[401] ,
    \itasegm1[400] ,
    \itasegm1[399] ,
    \itasegm1[398] ,
    \itasegm1[397] ,
    \itasegm1[396] ,
    \itasegm1[395] ,
    \itasegm1[394] ,
    \itasegm1[393] ,
    \itasegm1[392] }),
    .sel({\itasel1[347] ,
    \itasel1[346] ,
    \itasel1[345] ,
    \itasel1[344] ,
    \itasel1[343] ,
    \itasel1[342] ,
    \itasel1[341] ,
    \itasel1[340] ,
    \itasel1[339] ,
    \itasel1[338] ,
    \itasel1[337] ,
    \itasel1[336] }));
 ita3 ita3 (.clk(wb_clk_i),
    .segm({\itasegm1[41] ,
    \itasegm1[40] ,
    \itasegm1[39] ,
    \itasegm1[38] ,
    \itasegm1[37] ,
    \itasegm1[36] ,
    \itasegm1[35] ,
    \itasegm1[34] ,
    \itasegm1[33] ,
    \itasegm1[32] ,
    \itasegm1[31] ,
    \itasegm1[30] ,
    \itasegm1[29] ,
    \itasegm1[28] }),
    .sel({\itasel1[35] ,
    \itasel1[34] ,
    \itasel1[33] ,
    \itasel1[32] ,
    \itasel1[31] ,
    \itasel1[30] ,
    \itasel1[29] ,
    \itasel1[28] ,
    \itasel1[27] ,
    \itasel1[26] ,
    \itasel1[25] ,
    \itasel1[24] }));
 ita30 ita30 (.clk(wb_clk_i),
    .segm({\itasegm1[419] ,
    \itasegm1[418] ,
    \itasegm1[417] ,
    \itasegm1[416] ,
    \itasegm1[415] ,
    \itasegm1[414] ,
    \itasegm1[413] ,
    \itasegm1[412] ,
    \itasegm1[411] ,
    \itasegm1[410] ,
    \itasegm1[409] ,
    \itasegm1[408] ,
    \itasegm1[407] ,
    \itasegm1[406] }),
    .sel({\itasel1[359] ,
    \itasel1[358] ,
    \itasel1[357] ,
    \itasel1[356] ,
    \itasel1[355] ,
    \itasel1[354] ,
    \itasel1[353] ,
    \itasel1[352] ,
    \itasel1[351] ,
    \itasel1[350] ,
    \itasel1[349] ,
    \itasel1[348] }));
 ita31 ita31 (.clk(wb_clk_i),
    .segm({\itasegm1[433] ,
    \itasegm1[432] ,
    \itasegm1[431] ,
    \itasegm1[430] ,
    \itasegm1[429] ,
    \itasegm1[428] ,
    \itasegm1[427] ,
    \itasegm1[426] ,
    \itasegm1[425] ,
    \itasegm1[424] ,
    \itasegm1[423] ,
    \itasegm1[422] ,
    \itasegm1[421] ,
    \itasegm1[420] }),
    .sel({\itasel1[371] ,
    \itasel1[370] ,
    \itasel1[369] ,
    \itasel1[368] ,
    \itasel1[367] ,
    \itasel1[366] ,
    \itasel1[365] ,
    \itasel1[364] ,
    \itasel1[363] ,
    \itasel1[362] ,
    \itasel1[361] ,
    \itasel1[360] }));
 ita32 ita32 (.clk(wb_clk_i),
    .segm({\itasegm1[447] ,
    \itasegm1[446] ,
    \itasegm1[445] ,
    \itasegm1[444] ,
    \itasegm1[443] ,
    \itasegm1[442] ,
    \itasegm1[441] ,
    \itasegm1[440] ,
    \itasegm1[439] ,
    \itasegm1[438] ,
    \itasegm1[437] ,
    \itasegm1[436] ,
    \itasegm1[435] ,
    \itasegm1[434] }),
    .sel({\itasel1[383] ,
    \itasel1[382] ,
    \itasel1[381] ,
    \itasel1[380] ,
    \itasel1[379] ,
    \itasel1[378] ,
    \itasel1[377] ,
    \itasel1[376] ,
    \itasel1[375] ,
    \itasel1[374] ,
    \itasel1[373] ,
    \itasel1[372] }));
 ita33 ita33 (.clk(wb_clk_i),
    .segm({\itasegm1[461] ,
    \itasegm1[460] ,
    \itasegm1[459] ,
    \itasegm1[458] ,
    \itasegm1[457] ,
    \itasegm1[456] ,
    \itasegm1[455] ,
    \itasegm1[454] ,
    \itasegm1[453] ,
    \itasegm1[452] ,
    \itasegm1[451] ,
    \itasegm1[450] ,
    \itasegm1[449] ,
    \itasegm1[448] }),
    .sel({\itasel1[395] ,
    \itasel1[394] ,
    \itasel1[393] ,
    \itasel1[392] ,
    \itasel1[391] ,
    \itasel1[390] ,
    \itasel1[389] ,
    \itasel1[388] ,
    \itasel1[387] ,
    \itasel1[386] ,
    \itasel1[385] ,
    \itasel1[384] }));
 ita34 ita34 (.clk(wb_clk_i),
    .segm({\itasegm1[475] ,
    \itasegm1[474] ,
    \itasegm1[473] ,
    \itasegm1[472] ,
    \itasegm1[471] ,
    \itasegm1[470] ,
    \itasegm1[469] ,
    \itasegm1[468] ,
    \itasegm1[467] ,
    \itasegm1[466] ,
    \itasegm1[465] ,
    \itasegm1[464] ,
    \itasegm1[463] ,
    \itasegm1[462] }),
    .sel({\itasel1[407] ,
    \itasel1[406] ,
    \itasel1[405] ,
    \itasel1[404] ,
    \itasel1[403] ,
    \itasel1[402] ,
    \itasel1[401] ,
    \itasel1[400] ,
    \itasel1[399] ,
    \itasel1[398] ,
    \itasel1[397] ,
    \itasel1[396] }));
 ita35 ita35 (.clk(wb_clk_i),
    .segm({\itasegm1[489] ,
    \itasegm1[488] ,
    \itasegm1[487] ,
    \itasegm1[486] ,
    \itasegm1[485] ,
    \itasegm1[484] ,
    \itasegm1[483] ,
    \itasegm1[482] ,
    \itasegm1[481] ,
    \itasegm1[480] ,
    \itasegm1[479] ,
    \itasegm1[478] ,
    \itasegm1[477] ,
    \itasegm1[476] }),
    .sel({\itasel1[419] ,
    \itasel1[418] ,
    \itasel1[417] ,
    \itasel1[416] ,
    \itasel1[415] ,
    \itasel1[414] ,
    \itasel1[413] ,
    \itasel1[412] ,
    \itasel1[411] ,
    \itasel1[410] ,
    \itasel1[409] ,
    \itasel1[408] }));
 ita36 ita36 (.clk(wb_clk_i),
    .segm({\itasegm1[503] ,
    \itasegm1[502] ,
    \itasegm1[501] ,
    \itasegm1[500] ,
    \itasegm1[499] ,
    \itasegm1[498] ,
    \itasegm1[497] ,
    \itasegm1[496] ,
    \itasegm1[495] ,
    \itasegm1[494] ,
    \itasegm1[493] ,
    \itasegm1[492] ,
    \itasegm1[491] ,
    \itasegm1[490] }),
    .sel({\itasel1[431] ,
    \itasel1[430] ,
    \itasel1[429] ,
    \itasel1[428] ,
    \itasel1[427] ,
    \itasel1[426] ,
    \itasel1[425] ,
    \itasel1[424] ,
    \itasel1[423] ,
    \itasel1[422] ,
    \itasel1[421] ,
    \itasel1[420] }));
 ita37 ita37 (.clk(wb_clk_i),
    .segm({\itasegm1[517] ,
    \itasegm1[516] ,
    \itasegm1[515] ,
    \itasegm1[514] ,
    \itasegm1[513] ,
    \itasegm1[512] ,
    \itasegm1[511] ,
    \itasegm1[510] ,
    \itasegm1[509] ,
    \itasegm1[508] ,
    \itasegm1[507] ,
    \itasegm1[506] ,
    \itasegm1[505] ,
    \itasegm1[504] }),
    .sel({\itasel1[443] ,
    \itasel1[442] ,
    \itasel1[441] ,
    \itasel1[440] ,
    \itasel1[439] ,
    \itasel1[438] ,
    \itasel1[437] ,
    \itasel1[436] ,
    \itasel1[435] ,
    \itasel1[434] ,
    \itasel1[433] ,
    \itasel1[432] }));
 ita38 ita38 (.clk(wb_clk_i),
    .segm({\itasegm1[531] ,
    \itasegm1[530] ,
    \itasegm1[529] ,
    \itasegm1[528] ,
    \itasegm1[527] ,
    \itasegm1[526] ,
    \itasegm1[525] ,
    \itasegm1[524] ,
    \itasegm1[523] ,
    \itasegm1[522] ,
    \itasegm1[521] ,
    \itasegm1[520] ,
    \itasegm1[519] ,
    \itasegm1[518] }),
    .sel({\itasel1[455] ,
    \itasel1[454] ,
    \itasel1[453] ,
    \itasel1[452] ,
    \itasel1[451] ,
    \itasel1[450] ,
    \itasel1[449] ,
    \itasel1[448] ,
    \itasel1[447] ,
    \itasel1[446] ,
    \itasel1[445] ,
    \itasel1[444] }));
 ita39 ita39 (.clk(wb_clk_i),
    .segm({\itasegm1[545] ,
    \itasegm1[544] ,
    \itasegm1[543] ,
    \itasegm1[542] ,
    \itasegm1[541] ,
    \itasegm1[540] ,
    \itasegm1[539] ,
    \itasegm1[538] ,
    \itasegm1[537] ,
    \itasegm1[536] ,
    \itasegm1[535] ,
    \itasegm1[534] ,
    \itasegm1[533] ,
    \itasegm1[532] }),
    .sel({\itasel1[467] ,
    \itasel1[466] ,
    \itasel1[465] ,
    \itasel1[464] ,
    \itasel1[463] ,
    \itasel1[462] ,
    \itasel1[461] ,
    \itasel1[460] ,
    \itasel1[459] ,
    \itasel1[458] ,
    \itasel1[457] ,
    \itasel1[456] }));
 ita4 ita4 (.clk(wb_clk_i),
    .segm({\itasegm1[55] ,
    \itasegm1[54] ,
    \itasegm1[53] ,
    \itasegm1[52] ,
    \itasegm1[51] ,
    \itasegm1[50] ,
    \itasegm1[49] ,
    \itasegm1[48] ,
    \itasegm1[47] ,
    \itasegm1[46] ,
    \itasegm1[45] ,
    \itasegm1[44] ,
    \itasegm1[43] ,
    \itasegm1[42] }),
    .sel({\itasel1[47] ,
    \itasel1[46] ,
    \itasel1[45] ,
    \itasel1[44] ,
    \itasel1[43] ,
    \itasel1[42] ,
    \itasel1[41] ,
    \itasel1[40] ,
    \itasel1[39] ,
    \itasel1[38] ,
    \itasel1[37] ,
    \itasel1[36] }));
 ita40 ita40 (.clk(wb_clk_i),
    .segm({\itasegm1[559] ,
    \itasegm1[558] ,
    \itasegm1[557] ,
    \itasegm1[556] ,
    \itasegm1[555] ,
    \itasegm1[554] ,
    \itasegm1[553] ,
    \itasegm1[552] ,
    \itasegm1[551] ,
    \itasegm1[550] ,
    \itasegm1[549] ,
    \itasegm1[548] ,
    \itasegm1[547] ,
    \itasegm1[546] }),
    .sel({\itasel1[479] ,
    \itasel1[478] ,
    \itasel1[477] ,
    \itasel1[476] ,
    \itasel1[475] ,
    \itasel1[474] ,
    \itasel1[473] ,
    \itasel1[472] ,
    \itasel1[471] ,
    \itasel1[470] ,
    \itasel1[469] ,
    \itasel1[468] }));
 ita41 ita41 (.clk(wb_clk_i),
    .segm({\itasegm1[573] ,
    \itasegm1[572] ,
    \itasegm1[571] ,
    \itasegm1[570] ,
    \itasegm1[569] ,
    \itasegm1[568] ,
    \itasegm1[567] ,
    \itasegm1[566] ,
    \itasegm1[565] ,
    \itasegm1[564] ,
    \itasegm1[563] ,
    \itasegm1[562] ,
    \itasegm1[561] ,
    \itasegm1[560] }),
    .sel({\itasel1[491] ,
    \itasel1[490] ,
    \itasel1[489] ,
    \itasel1[488] ,
    \itasel1[487] ,
    \itasel1[486] ,
    \itasel1[485] ,
    \itasel1[484] ,
    \itasel1[483] ,
    \itasel1[482] ,
    \itasel1[481] ,
    \itasel1[480] }));
 ita42 ita42 (.clk(wb_clk_i),
    .segm({\itasegm1[587] ,
    \itasegm1[586] ,
    \itasegm1[585] ,
    \itasegm1[584] ,
    \itasegm1[583] ,
    \itasegm1[582] ,
    \itasegm1[581] ,
    \itasegm1[580] ,
    \itasegm1[579] ,
    \itasegm1[578] ,
    \itasegm1[577] ,
    \itasegm1[576] ,
    \itasegm1[575] ,
    \itasegm1[574] }),
    .sel({\itasel1[503] ,
    \itasel1[502] ,
    \itasel1[501] ,
    \itasel1[500] ,
    \itasel1[499] ,
    \itasel1[498] ,
    \itasel1[497] ,
    \itasel1[496] ,
    \itasel1[495] ,
    \itasel1[494] ,
    \itasel1[493] ,
    \itasel1[492] }));
 ita43 ita43 (.clk(wb_clk_i),
    .segm({\itasegm1[601] ,
    \itasegm1[600] ,
    \itasegm1[599] ,
    \itasegm1[598] ,
    \itasegm1[597] ,
    \itasegm1[596] ,
    \itasegm1[595] ,
    \itasegm1[594] ,
    \itasegm1[593] ,
    \itasegm1[592] ,
    \itasegm1[591] ,
    \itasegm1[590] ,
    \itasegm1[589] ,
    \itasegm1[588] }),
    .sel({\itasel1[515] ,
    \itasel1[514] ,
    \itasel1[513] ,
    \itasel1[512] ,
    \itasel1[511] ,
    \itasel1[510] ,
    \itasel1[509] ,
    \itasel1[508] ,
    \itasel1[507] ,
    \itasel1[506] ,
    \itasel1[505] ,
    \itasel1[504] }));
 ita44 ita44 (.clk(wb_clk_i),
    .segm({\itasegm1[615] ,
    \itasegm1[614] ,
    \itasegm1[613] ,
    \itasegm1[612] ,
    \itasegm1[611] ,
    \itasegm1[610] ,
    \itasegm1[609] ,
    \itasegm1[608] ,
    \itasegm1[607] ,
    \itasegm1[606] ,
    \itasegm1[605] ,
    \itasegm1[604] ,
    \itasegm1[603] ,
    \itasegm1[602] }),
    .sel({\itasel1[527] ,
    \itasel1[526] ,
    \itasel1[525] ,
    \itasel1[524] ,
    \itasel1[523] ,
    \itasel1[522] ,
    \itasel1[521] ,
    \itasel1[520] ,
    \itasel1[519] ,
    \itasel1[518] ,
    \itasel1[517] ,
    \itasel1[516] }));
 ita45 ita45 (.clk(wb_clk_i),
    .segm({\itasegm1[629] ,
    \itasegm1[628] ,
    \itasegm1[627] ,
    \itasegm1[626] ,
    \itasegm1[625] ,
    \itasegm1[624] ,
    \itasegm1[623] ,
    \itasegm1[622] ,
    \itasegm1[621] ,
    \itasegm1[620] ,
    \itasegm1[619] ,
    \itasegm1[618] ,
    \itasegm1[617] ,
    \itasegm1[616] }),
    .sel({\itasel1[539] ,
    \itasel1[538] ,
    \itasel1[537] ,
    \itasel1[536] ,
    \itasel1[535] ,
    \itasel1[534] ,
    \itasel1[533] ,
    \itasel1[532] ,
    \itasel1[531] ,
    \itasel1[530] ,
    \itasel1[529] ,
    \itasel1[528] }));
 ita46 ita46 (.clk(wb_clk_i),
    .segm({\itasegm1[643] ,
    \itasegm1[642] ,
    \itasegm1[641] ,
    \itasegm1[640] ,
    \itasegm1[639] ,
    \itasegm1[638] ,
    \itasegm1[637] ,
    \itasegm1[636] ,
    \itasegm1[635] ,
    \itasegm1[634] ,
    \itasegm1[633] ,
    \itasegm1[632] ,
    \itasegm1[631] ,
    \itasegm1[630] }),
    .sel({\itasel1[551] ,
    \itasel1[550] ,
    \itasel1[549] ,
    \itasel1[548] ,
    \itasel1[547] ,
    \itasel1[546] ,
    \itasel1[545] ,
    \itasel1[544] ,
    \itasel1[543] ,
    \itasel1[542] ,
    \itasel1[541] ,
    \itasel1[540] }));
 ita47 ita47 (.clk(wb_clk_i),
    .segm({\itasegm1[657] ,
    \itasegm1[656] ,
    \itasegm1[655] ,
    \itasegm1[654] ,
    \itasegm1[653] ,
    \itasegm1[652] ,
    \itasegm1[651] ,
    \itasegm1[650] ,
    \itasegm1[649] ,
    \itasegm1[648] ,
    \itasegm1[647] ,
    \itasegm1[646] ,
    \itasegm1[645] ,
    \itasegm1[644] }),
    .sel({\itasel1[563] ,
    \itasel1[562] ,
    \itasel1[561] ,
    \itasel1[560] ,
    \itasel1[559] ,
    \itasel1[558] ,
    \itasel1[557] ,
    \itasel1[556] ,
    \itasel1[555] ,
    \itasel1[554] ,
    \itasel1[553] ,
    \itasel1[552] }));
 ita48 ita48 (.clk(wb_clk_i),
    .segm({\itasegm1[671] ,
    \itasegm1[670] ,
    \itasegm1[669] ,
    \itasegm1[668] ,
    \itasegm1[667] ,
    \itasegm1[666] ,
    \itasegm1[665] ,
    \itasegm1[664] ,
    \itasegm1[663] ,
    \itasegm1[662] ,
    \itasegm1[661] ,
    \itasegm1[660] ,
    \itasegm1[659] ,
    \itasegm1[658] }),
    .sel({\itasel1[575] ,
    \itasel1[574] ,
    \itasel1[573] ,
    \itasel1[572] ,
    \itasel1[571] ,
    \itasel1[570] ,
    \itasel1[569] ,
    \itasel1[568] ,
    \itasel1[567] ,
    \itasel1[566] ,
    \itasel1[565] ,
    \itasel1[564] }));
 ita49 ita49 (.clk(wb_clk_i),
    .segm({\itasegm1[685] ,
    \itasegm1[684] ,
    \itasegm1[683] ,
    \itasegm1[682] ,
    \itasegm1[681] ,
    \itasegm1[680] ,
    \itasegm1[679] ,
    \itasegm1[678] ,
    \itasegm1[677] ,
    \itasegm1[676] ,
    \itasegm1[675] ,
    \itasegm1[674] ,
    \itasegm1[673] ,
    \itasegm1[672] }),
    .sel({\itasel1[587] ,
    \itasel1[586] ,
    \itasel1[585] ,
    \itasel1[584] ,
    \itasel1[583] ,
    \itasel1[582] ,
    \itasel1[581] ,
    \itasel1[580] ,
    \itasel1[579] ,
    \itasel1[578] ,
    \itasel1[577] ,
    \itasel1[576] }));
 ita5 ita5 (.clk(wb_clk_i),
    .segm({\itasegm1[69] ,
    \itasegm1[68] ,
    \itasegm1[67] ,
    \itasegm1[66] ,
    \itasegm1[65] ,
    \itasegm1[64] ,
    \itasegm1[63] ,
    \itasegm1[62] ,
    \itasegm1[61] ,
    \itasegm1[60] ,
    \itasegm1[59] ,
    \itasegm1[58] ,
    \itasegm1[57] ,
    \itasegm1[56] }),
    .sel({\itasel1[59] ,
    \itasel1[58] ,
    \itasel1[57] ,
    \itasel1[56] ,
    \itasel1[55] ,
    \itasel1[54] ,
    \itasel1[53] ,
    \itasel1[52] ,
    \itasel1[51] ,
    \itasel1[50] ,
    \itasel1[49] ,
    \itasel1[48] }));
 ita50 ita50 (.clk(wb_clk_i),
    .segm({\itasegm1[699] ,
    \itasegm1[698] ,
    \itasegm1[697] ,
    \itasegm1[696] ,
    \itasegm1[695] ,
    \itasegm1[694] ,
    \itasegm1[693] ,
    \itasegm1[692] ,
    \itasegm1[691] ,
    \itasegm1[690] ,
    \itasegm1[689] ,
    \itasegm1[688] ,
    \itasegm1[687] ,
    \itasegm1[686] }),
    .sel({\itasel1[599] ,
    \itasel1[598] ,
    \itasel1[597] ,
    \itasel1[596] ,
    \itasel1[595] ,
    \itasel1[594] ,
    \itasel1[593] ,
    \itasel1[592] ,
    \itasel1[591] ,
    \itasel1[590] ,
    \itasel1[589] ,
    \itasel1[588] }));
 ita51 ita51 (.clk(wb_clk_i),
    .segm({\itasegm1[713] ,
    \itasegm1[712] ,
    \itasegm1[711] ,
    \itasegm1[710] ,
    \itasegm1[709] ,
    \itasegm1[708] ,
    \itasegm1[707] ,
    \itasegm1[706] ,
    \itasegm1[705] ,
    \itasegm1[704] ,
    \itasegm1[703] ,
    \itasegm1[702] ,
    \itasegm1[701] ,
    \itasegm1[700] }),
    .sel({\itasel1[611] ,
    \itasel1[610] ,
    \itasel1[609] ,
    \itasel1[608] ,
    \itasel1[607] ,
    \itasel1[606] ,
    \itasel1[605] ,
    \itasel1[604] ,
    \itasel1[603] ,
    \itasel1[602] ,
    \itasel1[601] ,
    \itasel1[600] }));
 ita52 ita52 (.clk(wb_clk_i),
    .segm({\itasegm1[727] ,
    \itasegm1[726] ,
    \itasegm1[725] ,
    \itasegm1[724] ,
    \itasegm1[723] ,
    \itasegm1[722] ,
    \itasegm1[721] ,
    \itasegm1[720] ,
    \itasegm1[719] ,
    \itasegm1[718] ,
    \itasegm1[717] ,
    \itasegm1[716] ,
    \itasegm1[715] ,
    \itasegm1[714] }),
    .sel({\itasel1[623] ,
    \itasel1[622] ,
    \itasel1[621] ,
    \itasel1[620] ,
    \itasel1[619] ,
    \itasel1[618] ,
    \itasel1[617] ,
    \itasel1[616] ,
    \itasel1[615] ,
    \itasel1[614] ,
    \itasel1[613] ,
    \itasel1[612] }));
 ita53 ita53 (.clk(wb_clk_i),
    .segm({\itasegm1[741] ,
    \itasegm1[740] ,
    \itasegm1[739] ,
    \itasegm1[738] ,
    \itasegm1[737] ,
    \itasegm1[736] ,
    \itasegm1[735] ,
    \itasegm1[734] ,
    \itasegm1[733] ,
    \itasegm1[732] ,
    \itasegm1[731] ,
    \itasegm1[730] ,
    \itasegm1[729] ,
    \itasegm1[728] }),
    .sel({\itasel1[635] ,
    \itasel1[634] ,
    \itasel1[633] ,
    \itasel1[632] ,
    \itasel1[631] ,
    \itasel1[630] ,
    \itasel1[629] ,
    \itasel1[628] ,
    \itasel1[627] ,
    \itasel1[626] ,
    \itasel1[625] ,
    \itasel1[624] }));
 ita54 ita54 (.clk(wb_clk_i),
    .segm({\itasegm1[755] ,
    \itasegm1[754] ,
    \itasegm1[753] ,
    \itasegm1[752] ,
    \itasegm1[751] ,
    \itasegm1[750] ,
    \itasegm1[749] ,
    \itasegm1[748] ,
    \itasegm1[747] ,
    \itasegm1[746] ,
    \itasegm1[745] ,
    \itasegm1[744] ,
    \itasegm1[743] ,
    \itasegm1[742] }),
    .sel({\itasel1[647] ,
    \itasel1[646] ,
    \itasel1[645] ,
    \itasel1[644] ,
    \itasel1[643] ,
    \itasel1[642] ,
    \itasel1[641] ,
    \itasel1[640] ,
    \itasel1[639] ,
    \itasel1[638] ,
    \itasel1[637] ,
    \itasel1[636] }));
 ita55 ita55 (.clk(wb_clk_i),
    .segm({\itasegm1[769] ,
    \itasegm1[768] ,
    \itasegm1[767] ,
    \itasegm1[766] ,
    \itasegm1[765] ,
    \itasegm1[764] ,
    \itasegm1[763] ,
    \itasegm1[762] ,
    \itasegm1[761] ,
    \itasegm1[760] ,
    \itasegm1[759] ,
    \itasegm1[758] ,
    \itasegm1[757] ,
    \itasegm1[756] }),
    .sel({\itasel1[659] ,
    \itasel1[658] ,
    \itasel1[657] ,
    \itasel1[656] ,
    \itasel1[655] ,
    \itasel1[654] ,
    \itasel1[653] ,
    \itasel1[652] ,
    \itasel1[651] ,
    \itasel1[650] ,
    \itasel1[649] ,
    \itasel1[648] }));
 ita56 ita56 (.clk(wb_clk_i),
    .segm({\itasegm1[783] ,
    \itasegm1[782] ,
    \itasegm1[781] ,
    \itasegm1[780] ,
    \itasegm1[779] ,
    \itasegm1[778] ,
    \itasegm1[777] ,
    \itasegm1[776] ,
    \itasegm1[775] ,
    \itasegm1[774] ,
    \itasegm1[773] ,
    \itasegm1[772] ,
    \itasegm1[771] ,
    \itasegm1[770] }),
    .sel({\itasel1[671] ,
    \itasel1[670] ,
    \itasel1[669] ,
    \itasel1[668] ,
    \itasel1[667] ,
    \itasel1[666] ,
    \itasel1[665] ,
    \itasel1[664] ,
    \itasel1[663] ,
    \itasel1[662] ,
    \itasel1[661] ,
    \itasel1[660] }));
 ita57 ita57 (.clk(wb_clk_i),
    .segm({\itasegm1[797] ,
    \itasegm1[796] ,
    \itasegm1[795] ,
    \itasegm1[794] ,
    \itasegm1[793] ,
    \itasegm1[792] ,
    \itasegm1[791] ,
    \itasegm1[790] ,
    \itasegm1[789] ,
    \itasegm1[788] ,
    \itasegm1[787] ,
    \itasegm1[786] ,
    \itasegm1[785] ,
    \itasegm1[784] }),
    .sel({\itasel1[683] ,
    \itasel1[682] ,
    \itasel1[681] ,
    \itasel1[680] ,
    \itasel1[679] ,
    \itasel1[678] ,
    \itasel1[677] ,
    \itasel1[676] ,
    \itasel1[675] ,
    \itasel1[674] ,
    \itasel1[673] ,
    \itasel1[672] }));
 ita58 ita58 (.clk(wb_clk_i),
    .segm({\itasegm1[811] ,
    \itasegm1[810] ,
    \itasegm1[809] ,
    \itasegm1[808] ,
    \itasegm1[807] ,
    \itasegm1[806] ,
    \itasegm1[805] ,
    \itasegm1[804] ,
    \itasegm1[803] ,
    \itasegm1[802] ,
    \itasegm1[801] ,
    \itasegm1[800] ,
    \itasegm1[799] ,
    \itasegm1[798] }),
    .sel({\itasel1[695] ,
    \itasel1[694] ,
    \itasel1[693] ,
    \itasel1[692] ,
    \itasel1[691] ,
    \itasel1[690] ,
    \itasel1[689] ,
    \itasel1[688] ,
    \itasel1[687] ,
    \itasel1[686] ,
    \itasel1[685] ,
    \itasel1[684] }));
 ita59 ita59 (.clk(wb_clk_i),
    .segm({\itasegm1[825] ,
    \itasegm1[824] ,
    \itasegm1[823] ,
    \itasegm1[822] ,
    \itasegm1[821] ,
    \itasegm1[820] ,
    \itasegm1[819] ,
    \itasegm1[818] ,
    \itasegm1[817] ,
    \itasegm1[816] ,
    \itasegm1[815] ,
    \itasegm1[814] ,
    \itasegm1[813] ,
    \itasegm1[812] }),
    .sel({\itasel1[707] ,
    \itasel1[706] ,
    \itasel1[705] ,
    \itasel1[704] ,
    \itasel1[703] ,
    \itasel1[702] ,
    \itasel1[701] ,
    \itasel1[700] ,
    \itasel1[699] ,
    \itasel1[698] ,
    \itasel1[697] ,
    \itasel1[696] }));
 ita6 ita6 (.clk(wb_clk_i),
    .segm({\itasegm1[83] ,
    \itasegm1[82] ,
    \itasegm1[81] ,
    \itasegm1[80] ,
    \itasegm1[79] ,
    \itasegm1[78] ,
    \itasegm1[77] ,
    \itasegm1[76] ,
    \itasegm1[75] ,
    \itasegm1[74] ,
    \itasegm1[73] ,
    \itasegm1[72] ,
    \itasegm1[71] ,
    \itasegm1[70] }),
    .sel({\itasel1[71] ,
    \itasel1[70] ,
    \itasel1[69] ,
    \itasel1[68] ,
    \itasel1[67] ,
    \itasel1[66] ,
    \itasel1[65] ,
    \itasel1[64] ,
    \itasel1[63] ,
    \itasel1[62] ,
    \itasel1[61] ,
    \itasel1[60] }));
 ita60 ita60 (.clk(wb_clk_i),
    .segm({\itasegm1[839] ,
    \itasegm1[838] ,
    \itasegm1[837] ,
    \itasegm1[836] ,
    \itasegm1[835] ,
    \itasegm1[834] ,
    \itasegm1[833] ,
    \itasegm1[832] ,
    \itasegm1[831] ,
    \itasegm1[830] ,
    \itasegm1[829] ,
    \itasegm1[828] ,
    \itasegm1[827] ,
    \itasegm1[826] }),
    .sel({\itasel1[719] ,
    \itasel1[718] ,
    \itasel1[717] ,
    \itasel1[716] ,
    \itasel1[715] ,
    \itasel1[714] ,
    \itasel1[713] ,
    \itasel1[712] ,
    \itasel1[711] ,
    \itasel1[710] ,
    \itasel1[709] ,
    \itasel1[708] }));
 ita61 ita61 (.clk(wb_clk_i),
    .segm({\itasegm1[853] ,
    \itasegm1[852] ,
    \itasegm1[851] ,
    \itasegm1[850] ,
    \itasegm1[849] ,
    \itasegm1[848] ,
    \itasegm1[847] ,
    \itasegm1[846] ,
    \itasegm1[845] ,
    \itasegm1[844] ,
    \itasegm1[843] ,
    \itasegm1[842] ,
    \itasegm1[841] ,
    \itasegm1[840] }),
    .sel({\itasel1[731] ,
    \itasel1[730] ,
    \itasel1[729] ,
    \itasel1[728] ,
    \itasel1[727] ,
    \itasel1[726] ,
    \itasel1[725] ,
    \itasel1[724] ,
    \itasel1[723] ,
    \itasel1[722] ,
    \itasel1[721] ,
    \itasel1[720] }));
 ita62 ita62 (.clk(wb_clk_i),
    .segm({\itasegm1[867] ,
    \itasegm1[866] ,
    \itasegm1[865] ,
    \itasegm1[864] ,
    \itasegm1[863] ,
    \itasegm1[862] ,
    \itasegm1[861] ,
    \itasegm1[860] ,
    \itasegm1[859] ,
    \itasegm1[858] ,
    \itasegm1[857] ,
    \itasegm1[856] ,
    \itasegm1[855] ,
    \itasegm1[854] }),
    .sel({\itasel1[743] ,
    \itasel1[742] ,
    \itasel1[741] ,
    \itasel1[740] ,
    \itasel1[739] ,
    \itasel1[738] ,
    \itasel1[737] ,
    \itasel1[736] ,
    \itasel1[735] ,
    \itasel1[734] ,
    \itasel1[733] ,
    \itasel1[732] }));
 ita63 ita63 (.clk(wb_clk_i),
    .segm({\itasegm1[881] ,
    \itasegm1[880] ,
    \itasegm1[879] ,
    \itasegm1[878] ,
    \itasegm1[877] ,
    \itasegm1[876] ,
    \itasegm1[875] ,
    \itasegm1[874] ,
    \itasegm1[873] ,
    \itasegm1[872] ,
    \itasegm1[871] ,
    \itasegm1[870] ,
    \itasegm1[869] ,
    \itasegm1[868] }),
    .sel({\itasel1[755] ,
    \itasel1[754] ,
    \itasel1[753] ,
    \itasel1[752] ,
    \itasel1[751] ,
    \itasel1[750] ,
    \itasel1[749] ,
    \itasel1[748] ,
    \itasel1[747] ,
    \itasel1[746] ,
    \itasel1[745] ,
    \itasel1[744] }));
 ita64 ita64 (.clk(wb_clk_i),
    .segm({\itasegm1[895] ,
    \itasegm1[894] ,
    \itasegm1[893] ,
    \itasegm1[892] ,
    \itasegm1[891] ,
    \itasegm1[890] ,
    \itasegm1[889] ,
    \itasegm1[888] ,
    \itasegm1[887] ,
    \itasegm1[886] ,
    \itasegm1[885] ,
    \itasegm1[884] ,
    \itasegm1[883] ,
    \itasegm1[882] }),
    .sel({\itasel1[767] ,
    \itasel1[766] ,
    \itasel1[765] ,
    \itasel1[764] ,
    \itasel1[763] ,
    \itasel1[762] ,
    \itasel1[761] ,
    \itasel1[760] ,
    \itasel1[759] ,
    \itasel1[758] ,
    \itasel1[757] ,
    \itasel1[756] }));
 ita7 ita7 (.clk(wb_clk_i),
    .segm({\itasegm1[97] ,
    \itasegm1[96] ,
    \itasegm1[95] ,
    \itasegm1[94] ,
    \itasegm1[93] ,
    \itasegm1[92] ,
    \itasegm1[91] ,
    \itasegm1[90] ,
    \itasegm1[89] ,
    \itasegm1[88] ,
    \itasegm1[87] ,
    \itasegm1[86] ,
    \itasegm1[85] ,
    \itasegm1[84] }),
    .sel({\itasel1[83] ,
    \itasel1[82] ,
    \itasel1[81] ,
    \itasel1[80] ,
    \itasel1[79] ,
    \itasel1[78] ,
    \itasel1[77] ,
    \itasel1[76] ,
    \itasel1[75] ,
    \itasel1[74] ,
    \itasel1[73] ,
    \itasel1[72] }));
 ita8 ita8 (.clk(wb_clk_i),
    .segm({\itasegm1[111] ,
    \itasegm1[110] ,
    \itasegm1[109] ,
    \itasegm1[108] ,
    \itasegm1[107] ,
    \itasegm1[106] ,
    \itasegm1[105] ,
    \itasegm1[104] ,
    \itasegm1[103] ,
    \itasegm1[102] ,
    \itasegm1[101] ,
    \itasegm1[100] ,
    \itasegm1[99] ,
    \itasegm1[98] }),
    .sel({\itasel1[95] ,
    \itasel1[94] ,
    \itasel1[93] ,
    \itasel1[92] ,
    \itasel1[91] ,
    \itasel1[90] ,
    \itasel1[89] ,
    \itasel1[88] ,
    \itasel1[87] ,
    \itasel1[86] ,
    \itasel1[85] ,
    \itasel1[84] }));
 ita9 ita9 (.clk(wb_clk_i),
    .segm({\itasegm1[125] ,
    \itasegm1[124] ,
    \itasegm1[123] ,
    \itasegm1[122] ,
    \itasegm1[121] ,
    \itasegm1[120] ,
    \itasegm1[119] ,
    \itasegm1[118] ,
    \itasegm1[117] ,
    \itasegm1[116] ,
    \itasegm1[115] ,
    \itasegm1[114] ,
    \itasegm1[113] ,
    \itasegm1[112] }),
    .sel({\itasel1[107] ,
    \itasel1[106] ,
    \itasel1[105] ,
    \itasel1[104] ,
    \itasel1[103] ,
    \itasel1[102] ,
    \itasel1[101] ,
    \itasel1[100] ,
    \itasel1[99] ,
    \itasel1[98] ,
    \itasel1[97] ,
    \itasel1[96] }));
endmodule

