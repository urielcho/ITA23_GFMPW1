magic
tech gf180mcuD
magscale 1 10
timestamp 1699641626
<< metal1 >>
rect 27570 38558 27582 38610
rect 27634 38607 27646 38610
rect 28354 38607 28366 38610
rect 27634 38561 28366 38607
rect 27634 38558 27646 38561
rect 28354 38558 28366 38561
rect 28418 38558 28430 38610
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 18062 38274 18114 38286
rect 18062 38210 18114 38222
rect 22430 38274 22482 38286
rect 22430 38210 22482 38222
rect 26126 38274 26178 38286
rect 26126 38210 26178 38222
rect 17042 37998 17054 38050
rect 17106 37998 17118 38050
rect 21410 37998 21422 38050
rect 21474 37998 21486 38050
rect 25218 37998 25230 38050
rect 25282 37998 25294 38050
rect 28366 37938 28418 37950
rect 28366 37874 28418 37886
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 22094 37490 22146 37502
rect 22094 37426 22146 37438
rect 26798 37490 26850 37502
rect 26798 37426 26850 37438
rect 1710 37378 1762 37390
rect 1710 37314 1762 37326
rect 21074 37214 21086 37266
rect 21138 37214 21150 37266
rect 26002 37214 26014 37266
rect 26066 37214 26078 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 22318 36706 22370 36718
rect 22318 36642 22370 36654
rect 21298 36430 21310 36482
rect 21362 36430 21374 36482
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 21086 29314 21138 29326
rect 21086 29250 21138 29262
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 20738 28702 20750 28754
rect 20802 28702 20814 28754
rect 21646 28642 21698 28654
rect 17938 28590 17950 28642
rect 18002 28590 18014 28642
rect 21646 28578 21698 28590
rect 22094 28642 22146 28654
rect 22094 28578 22146 28590
rect 18610 28478 18622 28530
rect 18674 28478 18686 28530
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 18498 27806 18510 27858
rect 18562 27806 18574 27858
rect 21858 27806 21870 27858
rect 21922 27806 21934 27858
rect 19282 27694 19294 27746
rect 19346 27694 19358 27746
rect 21410 27694 21422 27746
rect 21474 27694 21486 27746
rect 22530 27694 22542 27746
rect 22594 27694 22606 27746
rect 24658 27694 24670 27746
rect 24722 27694 24734 27746
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 19630 27298 19682 27310
rect 19630 27234 19682 27246
rect 21310 27298 21362 27310
rect 21310 27234 21362 27246
rect 17390 27186 17442 27198
rect 16930 27134 16942 27186
rect 16994 27134 17006 27186
rect 26002 27134 26014 27186
rect 26066 27134 26078 27186
rect 17390 27122 17442 27134
rect 20526 27074 20578 27086
rect 22206 27074 22258 27086
rect 14130 27022 14142 27074
rect 14194 27022 14206 27074
rect 20738 27022 20750 27074
rect 20802 27022 20814 27074
rect 20526 27010 20578 27022
rect 22206 27010 22258 27022
rect 22542 27074 22594 27086
rect 23090 27022 23102 27074
rect 23154 27022 23166 27074
rect 22542 27010 22594 27022
rect 19742 26962 19794 26974
rect 14802 26910 14814 26962
rect 14866 26910 14878 26962
rect 19742 26898 19794 26910
rect 20078 26962 20130 26974
rect 20078 26898 20130 26910
rect 20414 26962 20466 26974
rect 20414 26898 20466 26910
rect 21422 26962 21474 26974
rect 21422 26898 21474 26910
rect 22654 26962 22706 26974
rect 23874 26910 23886 26962
rect 23938 26910 23950 26962
rect 22654 26898 22706 26910
rect 20302 26850 20354 26862
rect 20302 26786 20354 26798
rect 22318 26850 22370 26862
rect 22318 26786 22370 26798
rect 22430 26850 22482 26862
rect 22430 26786 22482 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 15710 26514 15762 26526
rect 15710 26450 15762 26462
rect 17838 26514 17890 26526
rect 17838 26450 17890 26462
rect 21646 26514 21698 26526
rect 21646 26450 21698 26462
rect 21870 26514 21922 26526
rect 21870 26450 21922 26462
rect 23662 26514 23714 26526
rect 23662 26450 23714 26462
rect 23886 26514 23938 26526
rect 23886 26450 23938 26462
rect 24446 26514 24498 26526
rect 24446 26450 24498 26462
rect 17390 26402 17442 26414
rect 17390 26338 17442 26350
rect 23102 26402 23154 26414
rect 23102 26338 23154 26350
rect 23438 26402 23490 26414
rect 23438 26338 23490 26350
rect 17614 26290 17666 26302
rect 17614 26226 17666 26238
rect 17950 26290 18002 26302
rect 21982 26290 22034 26302
rect 24558 26290 24610 26302
rect 21410 26238 21422 26290
rect 21474 26238 21486 26290
rect 24098 26238 24110 26290
rect 24162 26238 24174 26290
rect 17950 26226 18002 26238
rect 21982 26226 22034 26238
rect 24558 26226 24610 26238
rect 15822 26178 15874 26190
rect 15822 26114 15874 26126
rect 17726 26178 17778 26190
rect 22654 26178 22706 26190
rect 21522 26126 21534 26178
rect 21586 26126 21598 26178
rect 23986 26126 23998 26178
rect 24050 26126 24062 26178
rect 17726 26114 17778 26126
rect 22654 26114 22706 26126
rect 22990 26066 23042 26078
rect 22990 26002 23042 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 1934 25618 1986 25630
rect 40014 25618 40066 25630
rect 13906 25566 13918 25618
rect 13970 25566 13982 25618
rect 20402 25566 20414 25618
rect 20466 25566 20478 25618
rect 1934 25554 1986 25566
rect 40014 25554 40066 25566
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 16818 25454 16830 25506
rect 16882 25454 16894 25506
rect 17602 25454 17614 25506
rect 17666 25454 17678 25506
rect 37650 25454 37662 25506
rect 37714 25454 37726 25506
rect 26686 25394 26738 25406
rect 16034 25342 16046 25394
rect 16098 25342 16110 25394
rect 18274 25342 18286 25394
rect 18338 25342 18350 25394
rect 25554 25342 25566 25394
rect 25618 25342 25630 25394
rect 26686 25330 26738 25342
rect 26910 25394 26962 25406
rect 26910 25330 26962 25342
rect 27246 25394 27298 25406
rect 27246 25330 27298 25342
rect 27582 25394 27634 25406
rect 27582 25330 27634 25342
rect 21422 25282 21474 25294
rect 21422 25218 21474 25230
rect 25230 25282 25282 25294
rect 25230 25218 25282 25230
rect 27022 25282 27074 25294
rect 27022 25218 27074 25230
rect 27694 25282 27746 25294
rect 27694 25218 27746 25230
rect 27918 25282 27970 25294
rect 27918 25218 27970 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 16046 24946 16098 24958
rect 16046 24882 16098 24894
rect 17502 24946 17554 24958
rect 17502 24882 17554 24894
rect 18622 24946 18674 24958
rect 18622 24882 18674 24894
rect 28590 24946 28642 24958
rect 28590 24882 28642 24894
rect 15934 24834 15986 24846
rect 15934 24770 15986 24782
rect 28702 24834 28754 24846
rect 28702 24770 28754 24782
rect 18062 24722 18114 24734
rect 17826 24670 17838 24722
rect 17890 24670 17902 24722
rect 18062 24658 18114 24670
rect 18398 24722 18450 24734
rect 18610 24670 18622 24722
rect 18674 24670 18686 24722
rect 23874 24670 23886 24722
rect 23938 24670 23950 24722
rect 25330 24670 25342 24722
rect 25394 24670 25406 24722
rect 37650 24670 37662 24722
rect 37714 24670 37726 24722
rect 18398 24658 18450 24670
rect 18734 24610 18786 24622
rect 18734 24546 18786 24558
rect 19182 24610 19234 24622
rect 22642 24558 22654 24610
rect 22706 24558 22718 24610
rect 26114 24558 26126 24610
rect 26178 24558 26190 24610
rect 28242 24558 28254 24610
rect 28306 24558 28318 24610
rect 19182 24546 19234 24558
rect 16158 24498 16210 24510
rect 16158 24434 16210 24446
rect 40014 24498 40066 24510
rect 40014 24434 40066 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 19966 24162 20018 24174
rect 19966 24098 20018 24110
rect 1934 24050 1986 24062
rect 1934 23986 1986 23998
rect 15150 24050 15202 24062
rect 20078 24050 20130 24062
rect 16818 23998 16830 24050
rect 16882 23998 16894 24050
rect 15150 23986 15202 23998
rect 20078 23986 20130 23998
rect 21646 24050 21698 24062
rect 40014 24050 40066 24062
rect 24882 23998 24894 24050
rect 24946 23998 24958 24050
rect 26450 23998 26462 24050
rect 26514 23998 26526 24050
rect 28578 23998 28590 24050
rect 28642 23998 28654 24050
rect 21646 23986 21698 23998
rect 40014 23986 40066 23998
rect 17726 23938 17778 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 17726 23874 17778 23886
rect 18174 23938 18226 23950
rect 22082 23886 22094 23938
rect 22146 23886 22158 23938
rect 25666 23886 25678 23938
rect 25730 23886 25742 23938
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 18174 23874 18226 23886
rect 15822 23826 15874 23838
rect 15822 23762 15874 23774
rect 16830 23826 16882 23838
rect 16830 23762 16882 23774
rect 17278 23826 17330 23838
rect 22754 23774 22766 23826
rect 22818 23774 22830 23826
rect 17278 23762 17330 23774
rect 15598 23714 15650 23726
rect 15598 23650 15650 23662
rect 15710 23714 15762 23726
rect 15710 23650 15762 23662
rect 16718 23714 16770 23726
rect 16718 23650 16770 23662
rect 17054 23714 17106 23726
rect 17054 23650 17106 23662
rect 17838 23714 17890 23726
rect 17838 23650 17890 23662
rect 25342 23714 25394 23726
rect 25342 23650 25394 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 15486 23378 15538 23390
rect 15486 23314 15538 23326
rect 22318 23378 22370 23390
rect 22318 23314 22370 23326
rect 23102 23378 23154 23390
rect 23102 23314 23154 23326
rect 23662 23378 23714 23390
rect 23662 23314 23714 23326
rect 26126 23378 26178 23390
rect 26126 23314 26178 23326
rect 26350 23378 26402 23390
rect 26350 23314 26402 23326
rect 15598 23266 15650 23278
rect 14130 23214 14142 23266
rect 14194 23214 14206 23266
rect 15598 23202 15650 23214
rect 17838 23266 17890 23278
rect 17838 23202 17890 23214
rect 20750 23266 20802 23278
rect 20750 23202 20802 23214
rect 21198 23266 21250 23278
rect 21198 23202 21250 23214
rect 21534 23266 21586 23278
rect 21534 23202 21586 23214
rect 22654 23266 22706 23278
rect 22654 23202 22706 23214
rect 16046 23154 16098 23166
rect 4274 23102 4286 23154
rect 4338 23102 4350 23154
rect 14914 23102 14926 23154
rect 14978 23102 14990 23154
rect 16046 23090 16098 23102
rect 16158 23154 16210 23166
rect 16158 23090 16210 23102
rect 16606 23154 16658 23166
rect 16606 23090 16658 23102
rect 17950 23154 18002 23166
rect 21310 23154 21362 23166
rect 18162 23102 18174 23154
rect 18226 23102 18238 23154
rect 20962 23102 20974 23154
rect 21026 23102 21038 23154
rect 17950 23090 18002 23102
rect 21310 23090 21362 23102
rect 21870 23154 21922 23166
rect 21870 23090 21922 23102
rect 21982 23154 22034 23166
rect 22878 23154 22930 23166
rect 26014 23154 26066 23166
rect 22306 23102 22318 23154
rect 22370 23102 22382 23154
rect 23314 23102 23326 23154
rect 23378 23102 23390 23154
rect 21982 23090 22034 23102
rect 22878 23090 22930 23102
rect 26014 23090 26066 23102
rect 15822 23042 15874 23054
rect 12002 22990 12014 23042
rect 12066 22990 12078 23042
rect 15822 22978 15874 22990
rect 20526 23042 20578 23054
rect 20526 22978 20578 22990
rect 22990 23042 23042 23054
rect 22990 22978 23042 22990
rect 23774 23042 23826 23054
rect 23774 22978 23826 22990
rect 25342 23042 25394 23054
rect 25342 22978 25394 22990
rect 1934 22930 1986 22942
rect 17378 22878 17390 22930
rect 17442 22878 17454 22930
rect 1934 22866 1986 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 13806 22594 13858 22606
rect 21870 22594 21922 22606
rect 20066 22542 20078 22594
rect 20130 22542 20142 22594
rect 13806 22530 13858 22542
rect 21870 22530 21922 22542
rect 21982 22594 22034 22606
rect 21982 22530 22034 22542
rect 16158 22482 16210 22494
rect 16158 22418 16210 22430
rect 16830 22482 16882 22494
rect 16830 22418 16882 22430
rect 15262 22370 15314 22382
rect 15026 22318 15038 22370
rect 15090 22318 15102 22370
rect 15262 22306 15314 22318
rect 15486 22370 15538 22382
rect 16718 22370 16770 22382
rect 20302 22370 20354 22382
rect 21646 22370 21698 22382
rect 15698 22318 15710 22370
rect 15762 22318 15774 22370
rect 20066 22318 20078 22370
rect 20130 22318 20142 22370
rect 21410 22318 21422 22370
rect 21474 22318 21486 22370
rect 15486 22306 15538 22318
rect 16718 22306 16770 22318
rect 20302 22306 20354 22318
rect 21646 22306 21698 22318
rect 17602 22206 17614 22258
rect 17666 22206 17678 22258
rect 18610 22206 18622 22258
rect 18674 22206 18686 22258
rect 22978 22206 22990 22258
rect 23042 22206 23054 22258
rect 13582 22146 13634 22158
rect 13582 22082 13634 22094
rect 13694 22146 13746 22158
rect 13694 22082 13746 22094
rect 15374 22146 15426 22158
rect 15374 22082 15426 22094
rect 16942 22146 16994 22158
rect 16942 22082 16994 22094
rect 17166 22146 17218 22158
rect 17166 22082 17218 22094
rect 17950 22146 18002 22158
rect 17950 22082 18002 22094
rect 18958 22146 19010 22158
rect 18958 22082 19010 22094
rect 23326 22146 23378 22158
rect 23326 22082 23378 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 14814 21810 14866 21822
rect 25342 21810 25394 21822
rect 19170 21758 19182 21810
rect 19234 21758 19246 21810
rect 20514 21758 20526 21810
rect 20578 21758 20590 21810
rect 14814 21746 14866 21758
rect 25342 21746 25394 21758
rect 20190 21698 20242 21710
rect 25566 21698 25618 21710
rect 13570 21646 13582 21698
rect 13634 21646 13646 21698
rect 24098 21646 24110 21698
rect 24162 21646 24174 21698
rect 20190 21634 20242 21646
rect 25566 21634 25618 21646
rect 27022 21698 27074 21710
rect 27022 21634 27074 21646
rect 27470 21698 27522 21710
rect 27470 21634 27522 21646
rect 27582 21698 27634 21710
rect 27582 21634 27634 21646
rect 19518 21586 19570 21598
rect 20862 21586 20914 21598
rect 14354 21534 14366 21586
rect 14418 21534 14430 21586
rect 19842 21534 19854 21586
rect 19906 21534 19918 21586
rect 19518 21522 19570 21534
rect 20862 21522 20914 21534
rect 23774 21586 23826 21598
rect 23774 21522 23826 21534
rect 25230 21586 25282 21598
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 25230 21522 25282 21534
rect 25902 21474 25954 21486
rect 11442 21422 11454 21474
rect 11506 21422 11518 21474
rect 25902 21410 25954 21422
rect 19854 21362 19906 21374
rect 19854 21298 19906 21310
rect 27470 21362 27522 21374
rect 27470 21298 27522 21310
rect 40014 21362 40066 21374
rect 40014 21298 40066 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 17938 20974 17950 21026
rect 18002 20974 18014 21026
rect 1934 20914 1986 20926
rect 23874 20862 23886 20914
rect 23938 20862 23950 20914
rect 1934 20850 1986 20862
rect 18174 20802 18226 20814
rect 4274 20750 4286 20802
rect 4338 20750 4350 20802
rect 16706 20750 16718 20802
rect 16770 20750 16782 20802
rect 18174 20738 18226 20750
rect 18622 20802 18674 20814
rect 18622 20738 18674 20750
rect 19294 20802 19346 20814
rect 19294 20738 19346 20750
rect 20302 20802 20354 20814
rect 20302 20738 20354 20750
rect 20526 20802 20578 20814
rect 21298 20750 21310 20802
rect 21362 20750 21374 20802
rect 20526 20738 20578 20750
rect 14478 20690 14530 20702
rect 18958 20690 19010 20702
rect 16482 20638 16494 20690
rect 16546 20638 16558 20690
rect 14478 20626 14530 20638
rect 18958 20626 19010 20638
rect 14590 20578 14642 20590
rect 14590 20514 14642 20526
rect 19070 20578 19122 20590
rect 19070 20514 19122 20526
rect 20638 20578 20690 20590
rect 20638 20514 20690 20526
rect 20862 20578 20914 20590
rect 20862 20514 20914 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 15710 20242 15762 20254
rect 15710 20178 15762 20190
rect 22654 20242 22706 20254
rect 22654 20178 22706 20190
rect 15486 20130 15538 20142
rect 21534 20130 21586 20142
rect 22766 20130 22818 20142
rect 24334 20130 24386 20142
rect 19842 20078 19854 20130
rect 19906 20078 19918 20130
rect 20290 20078 20302 20130
rect 20354 20078 20366 20130
rect 21858 20078 21870 20130
rect 21922 20078 21934 20130
rect 23202 20078 23214 20130
rect 23266 20078 23278 20130
rect 26002 20078 26014 20130
rect 26066 20078 26078 20130
rect 15486 20066 15538 20078
rect 21534 20066 21586 20078
rect 22766 20066 22818 20078
rect 24334 20066 24386 20078
rect 15374 20018 15426 20030
rect 16270 20018 16322 20030
rect 13794 19966 13806 20018
rect 13858 19966 13870 20018
rect 15922 19966 15934 20018
rect 15986 19966 15998 20018
rect 15374 19954 15426 19966
rect 16270 19954 16322 19966
rect 16494 20018 16546 20030
rect 16494 19954 16546 19966
rect 16830 20018 16882 20030
rect 16830 19954 16882 19966
rect 17614 20018 17666 20030
rect 17614 19954 17666 19966
rect 18062 20018 18114 20030
rect 18062 19954 18114 19966
rect 19182 20018 19234 20030
rect 19182 19954 19234 19966
rect 19518 20018 19570 20030
rect 19518 19954 19570 19966
rect 20638 20018 20690 20030
rect 23886 20018 23938 20030
rect 22082 19966 22094 20018
rect 22146 19966 22158 20018
rect 23426 19966 23438 20018
rect 23490 19966 23502 20018
rect 20638 19954 20690 19966
rect 23886 19954 23938 19966
rect 24110 20018 24162 20030
rect 25330 19966 25342 20018
rect 25394 19966 25406 20018
rect 24110 19954 24162 19966
rect 14478 19906 14530 19918
rect 10882 19854 10894 19906
rect 10946 19854 10958 19906
rect 13010 19854 13022 19906
rect 13074 19854 13086 19906
rect 14478 19842 14530 19854
rect 14702 19906 14754 19918
rect 14702 19842 14754 19854
rect 15598 19906 15650 19918
rect 15598 19842 15650 19854
rect 16382 19906 16434 19918
rect 16382 19842 16434 19854
rect 20974 19906 21026 19918
rect 20974 19842 21026 19854
rect 23998 19906 24050 19918
rect 28130 19854 28142 19906
rect 28194 19854 28206 19906
rect 23998 19842 24050 19854
rect 14142 19794 14194 19806
rect 14142 19730 14194 19742
rect 17502 19794 17554 19806
rect 22542 19794 22594 19806
rect 18946 19742 18958 19794
rect 19010 19742 19022 19794
rect 17502 19730 17554 19742
rect 22542 19730 22594 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 23886 19458 23938 19470
rect 23886 19394 23938 19406
rect 14030 19346 14082 19358
rect 14030 19282 14082 19294
rect 21310 19346 21362 19358
rect 21310 19282 21362 19294
rect 23998 19346 24050 19358
rect 23998 19282 24050 19294
rect 24334 19346 24386 19358
rect 29822 19346 29874 19358
rect 28578 19294 28590 19346
rect 28642 19294 28654 19346
rect 24334 19282 24386 19294
rect 29822 19282 29874 19294
rect 40014 19346 40066 19358
rect 40014 19282 40066 19294
rect 22094 19234 22146 19246
rect 12226 19182 12238 19234
rect 12290 19182 12302 19234
rect 14802 19182 14814 19234
rect 14866 19182 14878 19234
rect 15474 19182 15486 19234
rect 15538 19182 15550 19234
rect 16482 19182 16494 19234
rect 16546 19182 16558 19234
rect 17378 19182 17390 19234
rect 17442 19182 17454 19234
rect 17826 19182 17838 19234
rect 17890 19182 17902 19234
rect 19954 19182 19966 19234
rect 20018 19182 20030 19234
rect 20290 19182 20302 19234
rect 20354 19182 20366 19234
rect 21858 19182 21870 19234
rect 21922 19182 21934 19234
rect 22094 19170 22146 19182
rect 24446 19234 24498 19246
rect 24446 19170 24498 19182
rect 25006 19234 25058 19246
rect 25006 19170 25058 19182
rect 25454 19234 25506 19246
rect 29038 19234 29090 19246
rect 25666 19182 25678 19234
rect 25730 19182 25742 19234
rect 25454 19170 25506 19182
rect 29038 19170 29090 19182
rect 29374 19234 29426 19246
rect 37650 19182 37662 19234
rect 37714 19182 37726 19234
rect 29374 19170 29426 19182
rect 12462 19122 12514 19134
rect 15026 19070 15038 19122
rect 15090 19070 15102 19122
rect 17266 19070 17278 19122
rect 17330 19070 17342 19122
rect 18162 19070 18174 19122
rect 18226 19070 18238 19122
rect 18722 19070 18734 19122
rect 18786 19070 18798 19122
rect 26450 19070 26462 19122
rect 26514 19070 26526 19122
rect 12462 19058 12514 19070
rect 24782 19010 24834 19022
rect 15698 18958 15710 19010
rect 15762 18958 15774 19010
rect 17154 18958 17166 19010
rect 17218 18958 17230 19010
rect 24782 18946 24834 18958
rect 24894 19010 24946 19022
rect 24894 18946 24946 18958
rect 29262 19010 29314 19022
rect 29262 18946 29314 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 16158 18674 16210 18686
rect 16158 18610 16210 18622
rect 25566 18674 25618 18686
rect 25566 18610 25618 18622
rect 25790 18674 25842 18686
rect 25790 18610 25842 18622
rect 20750 18562 20802 18574
rect 18498 18510 18510 18562
rect 18562 18510 18574 18562
rect 19506 18510 19518 18562
rect 19570 18510 19582 18562
rect 20750 18498 20802 18510
rect 25454 18562 25506 18574
rect 25454 18498 25506 18510
rect 14478 18450 14530 18462
rect 4274 18398 4286 18450
rect 4338 18398 4350 18450
rect 13570 18398 13582 18450
rect 13634 18398 13646 18450
rect 14478 18386 14530 18398
rect 14702 18450 14754 18462
rect 14702 18386 14754 18398
rect 15150 18450 15202 18462
rect 15150 18386 15202 18398
rect 16046 18450 16098 18462
rect 16046 18386 16098 18398
rect 16494 18450 16546 18462
rect 17490 18398 17502 18450
rect 17554 18398 17566 18450
rect 18722 18398 18734 18450
rect 18786 18398 18798 18450
rect 19394 18398 19406 18450
rect 19458 18398 19470 18450
rect 26114 18398 26126 18450
rect 26178 18398 26190 18450
rect 26786 18398 26798 18450
rect 26850 18398 26862 18450
rect 16494 18386 16546 18398
rect 24670 18338 24722 18350
rect 10658 18286 10670 18338
rect 10722 18286 10734 18338
rect 12786 18286 12798 18338
rect 12850 18286 12862 18338
rect 19058 18286 19070 18338
rect 19122 18286 19134 18338
rect 28914 18286 28926 18338
rect 28978 18286 28990 18338
rect 24670 18274 24722 18286
rect 1934 18226 1986 18238
rect 1934 18162 1986 18174
rect 13806 18226 13858 18238
rect 13806 18162 13858 18174
rect 14254 18226 14306 18238
rect 14254 18162 14306 18174
rect 20974 18226 21026 18238
rect 20974 18162 21026 18174
rect 21310 18226 21362 18238
rect 21310 18162 21362 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 13806 17890 13858 17902
rect 16046 17890 16098 17902
rect 14130 17838 14142 17890
rect 14194 17838 14206 17890
rect 17154 17838 17166 17890
rect 17218 17838 17230 17890
rect 19506 17838 19518 17890
rect 19570 17838 19582 17890
rect 13806 17826 13858 17838
rect 16046 17826 16098 17838
rect 13582 17778 13634 17790
rect 40014 17778 40066 17790
rect 17490 17726 17502 17778
rect 17554 17726 17566 17778
rect 18386 17726 18398 17778
rect 18450 17726 18462 17778
rect 13582 17714 13634 17726
rect 40014 17714 40066 17726
rect 15486 17666 15538 17678
rect 20302 17666 20354 17678
rect 12226 17614 12238 17666
rect 12290 17614 12302 17666
rect 16034 17614 16046 17666
rect 16098 17614 16110 17666
rect 17042 17614 17054 17666
rect 17106 17614 17118 17666
rect 18274 17614 18286 17666
rect 18338 17614 18350 17666
rect 19058 17614 19070 17666
rect 19122 17614 19134 17666
rect 19506 17614 19518 17666
rect 19570 17614 19582 17666
rect 15486 17602 15538 17614
rect 20302 17602 20354 17614
rect 22878 17666 22930 17678
rect 22878 17602 22930 17614
rect 23550 17666 23602 17678
rect 24670 17666 24722 17678
rect 24434 17614 24446 17666
rect 24498 17614 24510 17666
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 23550 17602 23602 17614
rect 24670 17602 24722 17614
rect 12462 17554 12514 17566
rect 12462 17490 12514 17502
rect 16382 17554 16434 17566
rect 23326 17554 23378 17566
rect 19954 17502 19966 17554
rect 20018 17502 20030 17554
rect 21634 17502 21646 17554
rect 21698 17502 21710 17554
rect 16382 17490 16434 17502
rect 23326 17490 23378 17502
rect 23886 17554 23938 17566
rect 23886 17490 23938 17502
rect 25006 17554 25058 17566
rect 25006 17490 25058 17502
rect 15598 17442 15650 17454
rect 15598 17378 15650 17390
rect 15822 17442 15874 17454
rect 15822 17378 15874 17390
rect 21310 17442 21362 17454
rect 21310 17378 21362 17390
rect 23214 17442 23266 17454
rect 23214 17378 23266 17390
rect 23998 17442 24050 17454
rect 23998 17378 24050 17390
rect 24110 17442 24162 17454
rect 24110 17378 24162 17390
rect 24894 17442 24946 17454
rect 24894 17378 24946 17390
rect 25678 17442 25730 17454
rect 25678 17378 25730 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 17950 17106 18002 17118
rect 17950 17042 18002 17054
rect 25790 17106 25842 17118
rect 25790 17042 25842 17054
rect 15486 16994 15538 17006
rect 26462 16994 26514 17006
rect 16482 16942 16494 16994
rect 16546 16942 16558 16994
rect 20850 16942 20862 16994
rect 20914 16942 20926 16994
rect 15486 16930 15538 16942
rect 26462 16930 26514 16942
rect 26574 16994 26626 17006
rect 26574 16930 26626 16942
rect 18062 16882 18114 16894
rect 25566 16882 25618 16894
rect 15698 16830 15710 16882
rect 15762 16830 15774 16882
rect 16258 16830 16270 16882
rect 16322 16830 16334 16882
rect 24322 16830 24334 16882
rect 24386 16830 24398 16882
rect 18062 16818 18114 16830
rect 25566 16818 25618 16830
rect 26238 16882 26290 16894
rect 37650 16830 37662 16882
rect 37714 16830 37726 16882
rect 26238 16818 26290 16830
rect 25678 16770 25730 16782
rect 39890 16718 39902 16770
rect 39954 16718 39966 16770
rect 25678 16706 25730 16718
rect 26574 16658 26626 16670
rect 26574 16594 26626 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 19966 16322 20018 16334
rect 19966 16258 20018 16270
rect 21422 16322 21474 16334
rect 21422 16258 21474 16270
rect 22542 16322 22594 16334
rect 22542 16258 22594 16270
rect 17726 16210 17778 16222
rect 22094 16210 22146 16222
rect 40014 16210 40066 16222
rect 14242 16158 14254 16210
rect 14306 16158 14318 16210
rect 16370 16158 16382 16210
rect 16434 16158 16446 16210
rect 17154 16158 17166 16210
rect 17218 16158 17230 16210
rect 20290 16158 20302 16210
rect 20354 16158 20366 16210
rect 23762 16158 23774 16210
rect 23826 16158 23838 16210
rect 25890 16158 25902 16210
rect 25954 16158 25966 16210
rect 17726 16146 17778 16158
rect 22094 16146 22146 16158
rect 40014 16146 40066 16158
rect 16718 16098 16770 16110
rect 21310 16098 21362 16110
rect 13458 16046 13470 16098
rect 13522 16046 13534 16098
rect 18050 16046 18062 16098
rect 18114 16046 18126 16098
rect 19170 16046 19182 16098
rect 19234 16046 19246 16098
rect 16718 16034 16770 16046
rect 21310 16034 21362 16046
rect 22430 16098 22482 16110
rect 26238 16098 26290 16110
rect 22978 16046 22990 16098
rect 23042 16046 23054 16098
rect 28018 16046 28030 16098
rect 28082 16046 28094 16098
rect 37650 16046 37662 16098
rect 37714 16046 37726 16098
rect 22430 16034 22482 16046
rect 26238 16034 26290 16046
rect 22542 15986 22594 15998
rect 18162 15934 18174 15986
rect 18226 15934 18238 15986
rect 26562 15934 26574 15986
rect 26626 15934 26638 15986
rect 22542 15922 22594 15934
rect 20190 15874 20242 15886
rect 19058 15822 19070 15874
rect 19122 15822 19134 15874
rect 28242 15822 28254 15874
rect 28306 15822 28318 15874
rect 20190 15810 20242 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 17726 15538 17778 15550
rect 17378 15486 17390 15538
rect 17442 15486 17454 15538
rect 17726 15474 17778 15486
rect 22654 15538 22706 15550
rect 22654 15474 22706 15486
rect 24670 15538 24722 15550
rect 24670 15474 24722 15486
rect 15598 15426 15650 15438
rect 18050 15374 18062 15426
rect 18114 15374 18126 15426
rect 20066 15374 20078 15426
rect 20130 15374 20142 15426
rect 26338 15374 26350 15426
rect 26402 15374 26414 15426
rect 15598 15362 15650 15374
rect 16258 15262 16270 15314
rect 16322 15262 16334 15314
rect 18274 15262 18286 15314
rect 18338 15262 18350 15314
rect 19282 15262 19294 15314
rect 19346 15262 19358 15314
rect 25554 15262 25566 15314
rect 25618 15262 25630 15314
rect 15922 15150 15934 15202
rect 15986 15150 15998 15202
rect 22194 15150 22206 15202
rect 22258 15150 22270 15202
rect 28466 15150 28478 15202
rect 28530 15150 28542 15202
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 21646 14754 21698 14766
rect 23986 14702 23998 14754
rect 24050 14702 24062 14754
rect 21646 14690 21698 14702
rect 18398 14642 18450 14654
rect 15810 14590 15822 14642
rect 15874 14590 15886 14642
rect 17938 14590 17950 14642
rect 18002 14590 18014 14642
rect 18398 14578 18450 14590
rect 24670 14642 24722 14654
rect 24670 14578 24722 14590
rect 22430 14530 22482 14542
rect 15138 14478 15150 14530
rect 15202 14478 15214 14530
rect 22430 14466 22482 14478
rect 23438 14530 23490 14542
rect 23986 14478 23998 14530
rect 24050 14478 24062 14530
rect 23438 14466 23490 14478
rect 21870 14418 21922 14430
rect 21870 14354 21922 14366
rect 22766 14418 22818 14430
rect 24558 14418 24610 14430
rect 23650 14366 23662 14418
rect 23714 14366 23726 14418
rect 22766 14354 22818 14366
rect 24558 14354 24610 14366
rect 24782 14306 24834 14318
rect 21298 14254 21310 14306
rect 21362 14254 21374 14306
rect 23874 14254 23886 14306
rect 23938 14254 23950 14306
rect 24782 14242 24834 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 18286 13858 18338 13870
rect 18286 13794 18338 13806
rect 20190 13858 20242 13870
rect 20190 13794 20242 13806
rect 21086 13858 21138 13870
rect 21086 13794 21138 13806
rect 22766 13858 22818 13870
rect 22766 13794 22818 13806
rect 22990 13858 23042 13870
rect 22990 13794 23042 13806
rect 18498 13694 18510 13746
rect 18562 13694 18574 13746
rect 20738 13694 20750 13746
rect 20802 13694 20814 13746
rect 20078 13522 20130 13534
rect 20078 13458 20130 13470
rect 20414 13522 20466 13534
rect 20414 13458 20466 13470
rect 20750 13522 20802 13534
rect 20750 13458 20802 13470
rect 22654 13522 22706 13534
rect 22654 13458 22706 13470
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 21758 13186 21810 13198
rect 21758 13122 21810 13134
rect 20750 13074 20802 13086
rect 22766 13074 22818 13086
rect 18162 13022 18174 13074
rect 18226 13022 18238 13074
rect 20290 13022 20302 13074
rect 20354 13022 20366 13074
rect 21410 13022 21422 13074
rect 21474 13022 21486 13074
rect 23874 13022 23886 13074
rect 23938 13022 23950 13074
rect 26002 13022 26014 13074
rect 26066 13022 26078 13074
rect 20750 13010 20802 13022
rect 22766 13010 22818 13022
rect 17490 12910 17502 12962
rect 17554 12910 17566 12962
rect 23090 12910 23102 12962
rect 23154 12910 23166 12962
rect 21534 12850 21586 12862
rect 21534 12786 21586 12798
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 23774 12402 23826 12414
rect 18274 12350 18286 12402
rect 18338 12350 18350 12402
rect 23774 12338 23826 12350
rect 18846 12290 18898 12302
rect 21186 12238 21198 12290
rect 21250 12238 21262 12290
rect 18846 12226 18898 12238
rect 18622 12178 18674 12190
rect 20514 12126 20526 12178
rect 20578 12126 20590 12178
rect 18622 12114 18674 12126
rect 23314 12014 23326 12066
rect 23378 12014 23390 12066
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 26798 5234 26850 5246
rect 26798 5170 26850 5182
rect 25778 5070 25790 5122
rect 25842 5070 25854 5122
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 25218 4286 25230 4338
rect 25282 4286 25294 4338
rect 26238 4114 26290 4126
rect 26238 4050 26290 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 20738 3502 20750 3554
rect 20802 3502 20814 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 19070 3330 19122 3342
rect 19070 3266 19122 3278
rect 21758 3330 21810 3342
rect 21758 3266 21810 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 27582 38558 27634 38610
rect 28366 38558 28418 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 18062 38222 18114 38274
rect 22430 38222 22482 38274
rect 26126 38222 26178 38274
rect 17054 37998 17106 38050
rect 21422 37998 21474 38050
rect 25230 37998 25282 38050
rect 28366 37886 28418 37938
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 22094 37438 22146 37490
rect 26798 37438 26850 37490
rect 1710 37326 1762 37378
rect 21086 37214 21138 37266
rect 26014 37214 26066 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 22318 36654 22370 36706
rect 21310 36430 21362 36482
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 21086 29262 21138 29314
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 20750 28702 20802 28754
rect 17950 28590 18002 28642
rect 21646 28590 21698 28642
rect 22094 28590 22146 28642
rect 18622 28478 18674 28530
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 18510 27806 18562 27858
rect 21870 27806 21922 27858
rect 19294 27694 19346 27746
rect 21422 27694 21474 27746
rect 22542 27694 22594 27746
rect 24670 27694 24722 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 19630 27246 19682 27298
rect 21310 27246 21362 27298
rect 16942 27134 16994 27186
rect 17390 27134 17442 27186
rect 26014 27134 26066 27186
rect 14142 27022 14194 27074
rect 20526 27022 20578 27074
rect 20750 27022 20802 27074
rect 22206 27022 22258 27074
rect 22542 27022 22594 27074
rect 23102 27022 23154 27074
rect 14814 26910 14866 26962
rect 19742 26910 19794 26962
rect 20078 26910 20130 26962
rect 20414 26910 20466 26962
rect 21422 26910 21474 26962
rect 22654 26910 22706 26962
rect 23886 26910 23938 26962
rect 20302 26798 20354 26850
rect 22318 26798 22370 26850
rect 22430 26798 22482 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 15710 26462 15762 26514
rect 17838 26462 17890 26514
rect 21646 26462 21698 26514
rect 21870 26462 21922 26514
rect 23662 26462 23714 26514
rect 23886 26462 23938 26514
rect 24446 26462 24498 26514
rect 17390 26350 17442 26402
rect 23102 26350 23154 26402
rect 23438 26350 23490 26402
rect 17614 26238 17666 26290
rect 17950 26238 18002 26290
rect 21422 26238 21474 26290
rect 21982 26238 22034 26290
rect 24110 26238 24162 26290
rect 24558 26238 24610 26290
rect 15822 26126 15874 26178
rect 17726 26126 17778 26178
rect 21534 26126 21586 26178
rect 22654 26126 22706 26178
rect 23998 26126 24050 26178
rect 22990 26014 23042 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 1934 25566 1986 25618
rect 13918 25566 13970 25618
rect 20414 25566 20466 25618
rect 40014 25566 40066 25618
rect 4286 25454 4338 25506
rect 16830 25454 16882 25506
rect 17614 25454 17666 25506
rect 37662 25454 37714 25506
rect 16046 25342 16098 25394
rect 18286 25342 18338 25394
rect 25566 25342 25618 25394
rect 26686 25342 26738 25394
rect 26910 25342 26962 25394
rect 27246 25342 27298 25394
rect 27582 25342 27634 25394
rect 21422 25230 21474 25282
rect 25230 25230 25282 25282
rect 27022 25230 27074 25282
rect 27694 25230 27746 25282
rect 27918 25230 27970 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 16046 24894 16098 24946
rect 17502 24894 17554 24946
rect 18622 24894 18674 24946
rect 28590 24894 28642 24946
rect 15934 24782 15986 24834
rect 28702 24782 28754 24834
rect 17838 24670 17890 24722
rect 18062 24670 18114 24722
rect 18398 24670 18450 24722
rect 18622 24670 18674 24722
rect 23886 24670 23938 24722
rect 25342 24670 25394 24722
rect 37662 24670 37714 24722
rect 18734 24558 18786 24610
rect 19182 24558 19234 24610
rect 22654 24558 22706 24610
rect 26126 24558 26178 24610
rect 28254 24558 28306 24610
rect 16158 24446 16210 24498
rect 40014 24446 40066 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 19966 24110 20018 24162
rect 1934 23998 1986 24050
rect 15150 23998 15202 24050
rect 16830 23998 16882 24050
rect 20078 23998 20130 24050
rect 21646 23998 21698 24050
rect 24894 23998 24946 24050
rect 26462 23998 26514 24050
rect 28590 23998 28642 24050
rect 40014 23998 40066 24050
rect 4286 23886 4338 23938
rect 17726 23886 17778 23938
rect 18174 23886 18226 23938
rect 22094 23886 22146 23938
rect 25678 23886 25730 23938
rect 37662 23886 37714 23938
rect 15822 23774 15874 23826
rect 16830 23774 16882 23826
rect 17278 23774 17330 23826
rect 22766 23774 22818 23826
rect 15598 23662 15650 23714
rect 15710 23662 15762 23714
rect 16718 23662 16770 23714
rect 17054 23662 17106 23714
rect 17838 23662 17890 23714
rect 25342 23662 25394 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 15486 23326 15538 23378
rect 22318 23326 22370 23378
rect 23102 23326 23154 23378
rect 23662 23326 23714 23378
rect 26126 23326 26178 23378
rect 26350 23326 26402 23378
rect 14142 23214 14194 23266
rect 15598 23214 15650 23266
rect 17838 23214 17890 23266
rect 20750 23214 20802 23266
rect 21198 23214 21250 23266
rect 21534 23214 21586 23266
rect 22654 23214 22706 23266
rect 4286 23102 4338 23154
rect 14926 23102 14978 23154
rect 16046 23102 16098 23154
rect 16158 23102 16210 23154
rect 16606 23102 16658 23154
rect 17950 23102 18002 23154
rect 18174 23102 18226 23154
rect 20974 23102 21026 23154
rect 21310 23102 21362 23154
rect 21870 23102 21922 23154
rect 21982 23102 22034 23154
rect 22318 23102 22370 23154
rect 22878 23102 22930 23154
rect 23326 23102 23378 23154
rect 26014 23102 26066 23154
rect 12014 22990 12066 23042
rect 15822 22990 15874 23042
rect 20526 22990 20578 23042
rect 22990 22990 23042 23042
rect 23774 22990 23826 23042
rect 25342 22990 25394 23042
rect 1934 22878 1986 22930
rect 17390 22878 17442 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 13806 22542 13858 22594
rect 20078 22542 20130 22594
rect 21870 22542 21922 22594
rect 21982 22542 22034 22594
rect 16158 22430 16210 22482
rect 16830 22430 16882 22482
rect 15038 22318 15090 22370
rect 15262 22318 15314 22370
rect 15486 22318 15538 22370
rect 15710 22318 15762 22370
rect 16718 22318 16770 22370
rect 20078 22318 20130 22370
rect 20302 22318 20354 22370
rect 21422 22318 21474 22370
rect 21646 22318 21698 22370
rect 17614 22206 17666 22258
rect 18622 22206 18674 22258
rect 22990 22206 23042 22258
rect 13582 22094 13634 22146
rect 13694 22094 13746 22146
rect 15374 22094 15426 22146
rect 16942 22094 16994 22146
rect 17166 22094 17218 22146
rect 17950 22094 18002 22146
rect 18958 22094 19010 22146
rect 23326 22094 23378 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 14814 21758 14866 21810
rect 19182 21758 19234 21810
rect 20526 21758 20578 21810
rect 25342 21758 25394 21810
rect 13582 21646 13634 21698
rect 20190 21646 20242 21698
rect 24110 21646 24162 21698
rect 25566 21646 25618 21698
rect 27022 21646 27074 21698
rect 27470 21646 27522 21698
rect 27582 21646 27634 21698
rect 14366 21534 14418 21586
rect 19518 21534 19570 21586
rect 19854 21534 19906 21586
rect 20862 21534 20914 21586
rect 23774 21534 23826 21586
rect 25230 21534 25282 21586
rect 37662 21534 37714 21586
rect 11454 21422 11506 21474
rect 25902 21422 25954 21474
rect 19854 21310 19906 21362
rect 27470 21310 27522 21362
rect 40014 21310 40066 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 17950 20974 18002 21026
rect 1934 20862 1986 20914
rect 23886 20862 23938 20914
rect 4286 20750 4338 20802
rect 16718 20750 16770 20802
rect 18174 20750 18226 20802
rect 18622 20750 18674 20802
rect 19294 20750 19346 20802
rect 20302 20750 20354 20802
rect 20526 20750 20578 20802
rect 21310 20750 21362 20802
rect 14478 20638 14530 20690
rect 16494 20638 16546 20690
rect 18958 20638 19010 20690
rect 14590 20526 14642 20578
rect 19070 20526 19122 20578
rect 20638 20526 20690 20578
rect 20862 20526 20914 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 15710 20190 15762 20242
rect 22654 20190 22706 20242
rect 15486 20078 15538 20130
rect 19854 20078 19906 20130
rect 20302 20078 20354 20130
rect 21534 20078 21586 20130
rect 21870 20078 21922 20130
rect 22766 20078 22818 20130
rect 23214 20078 23266 20130
rect 24334 20078 24386 20130
rect 26014 20078 26066 20130
rect 13806 19966 13858 20018
rect 15374 19966 15426 20018
rect 15934 19966 15986 20018
rect 16270 19966 16322 20018
rect 16494 19966 16546 20018
rect 16830 19966 16882 20018
rect 17614 19966 17666 20018
rect 18062 19966 18114 20018
rect 19182 19966 19234 20018
rect 19518 19966 19570 20018
rect 20638 19966 20690 20018
rect 22094 19966 22146 20018
rect 23438 19966 23490 20018
rect 23886 19966 23938 20018
rect 24110 19966 24162 20018
rect 25342 19966 25394 20018
rect 10894 19854 10946 19906
rect 13022 19854 13074 19906
rect 14478 19854 14530 19906
rect 14702 19854 14754 19906
rect 15598 19854 15650 19906
rect 16382 19854 16434 19906
rect 20974 19854 21026 19906
rect 23998 19854 24050 19906
rect 28142 19854 28194 19906
rect 14142 19742 14194 19794
rect 17502 19742 17554 19794
rect 18958 19742 19010 19794
rect 22542 19742 22594 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 23886 19406 23938 19458
rect 14030 19294 14082 19346
rect 21310 19294 21362 19346
rect 23998 19294 24050 19346
rect 24334 19294 24386 19346
rect 28590 19294 28642 19346
rect 29822 19294 29874 19346
rect 40014 19294 40066 19346
rect 12238 19182 12290 19234
rect 14814 19182 14866 19234
rect 15486 19182 15538 19234
rect 16494 19182 16546 19234
rect 17390 19182 17442 19234
rect 17838 19182 17890 19234
rect 19966 19182 20018 19234
rect 20302 19182 20354 19234
rect 21870 19182 21922 19234
rect 22094 19182 22146 19234
rect 24446 19182 24498 19234
rect 25006 19182 25058 19234
rect 25454 19182 25506 19234
rect 25678 19182 25730 19234
rect 29038 19182 29090 19234
rect 29374 19182 29426 19234
rect 37662 19182 37714 19234
rect 12462 19070 12514 19122
rect 15038 19070 15090 19122
rect 17278 19070 17330 19122
rect 18174 19070 18226 19122
rect 18734 19070 18786 19122
rect 26462 19070 26514 19122
rect 15710 18958 15762 19010
rect 17166 18958 17218 19010
rect 24782 18958 24834 19010
rect 24894 18958 24946 19010
rect 29262 18958 29314 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 16158 18622 16210 18674
rect 25566 18622 25618 18674
rect 25790 18622 25842 18674
rect 18510 18510 18562 18562
rect 19518 18510 19570 18562
rect 20750 18510 20802 18562
rect 25454 18510 25506 18562
rect 4286 18398 4338 18450
rect 13582 18398 13634 18450
rect 14478 18398 14530 18450
rect 14702 18398 14754 18450
rect 15150 18398 15202 18450
rect 16046 18398 16098 18450
rect 16494 18398 16546 18450
rect 17502 18398 17554 18450
rect 18734 18398 18786 18450
rect 19406 18398 19458 18450
rect 26126 18398 26178 18450
rect 26798 18398 26850 18450
rect 10670 18286 10722 18338
rect 12798 18286 12850 18338
rect 19070 18286 19122 18338
rect 24670 18286 24722 18338
rect 28926 18286 28978 18338
rect 1934 18174 1986 18226
rect 13806 18174 13858 18226
rect 14254 18174 14306 18226
rect 20974 18174 21026 18226
rect 21310 18174 21362 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 13806 17838 13858 17890
rect 14142 17838 14194 17890
rect 16046 17838 16098 17890
rect 17166 17838 17218 17890
rect 19518 17838 19570 17890
rect 13582 17726 13634 17778
rect 17502 17726 17554 17778
rect 18398 17726 18450 17778
rect 40014 17726 40066 17778
rect 12238 17614 12290 17666
rect 15486 17614 15538 17666
rect 16046 17614 16098 17666
rect 17054 17614 17106 17666
rect 18286 17614 18338 17666
rect 19070 17614 19122 17666
rect 19518 17614 19570 17666
rect 20302 17614 20354 17666
rect 22878 17614 22930 17666
rect 23550 17614 23602 17666
rect 24446 17614 24498 17666
rect 24670 17614 24722 17666
rect 37662 17614 37714 17666
rect 12462 17502 12514 17554
rect 16382 17502 16434 17554
rect 19966 17502 20018 17554
rect 21646 17502 21698 17554
rect 23326 17502 23378 17554
rect 23886 17502 23938 17554
rect 25006 17502 25058 17554
rect 15598 17390 15650 17442
rect 15822 17390 15874 17442
rect 21310 17390 21362 17442
rect 23214 17390 23266 17442
rect 23998 17390 24050 17442
rect 24110 17390 24162 17442
rect 24894 17390 24946 17442
rect 25678 17390 25730 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 17950 17054 18002 17106
rect 25790 17054 25842 17106
rect 15486 16942 15538 16994
rect 16494 16942 16546 16994
rect 20862 16942 20914 16994
rect 26462 16942 26514 16994
rect 26574 16942 26626 16994
rect 15710 16830 15762 16882
rect 16270 16830 16322 16882
rect 18062 16830 18114 16882
rect 24334 16830 24386 16882
rect 25566 16830 25618 16882
rect 26238 16830 26290 16882
rect 37662 16830 37714 16882
rect 25678 16718 25730 16770
rect 39902 16718 39954 16770
rect 26574 16606 26626 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 19966 16270 20018 16322
rect 21422 16270 21474 16322
rect 22542 16270 22594 16322
rect 14254 16158 14306 16210
rect 16382 16158 16434 16210
rect 17166 16158 17218 16210
rect 17726 16158 17778 16210
rect 20302 16158 20354 16210
rect 22094 16158 22146 16210
rect 23774 16158 23826 16210
rect 25902 16158 25954 16210
rect 40014 16158 40066 16210
rect 13470 16046 13522 16098
rect 16718 16046 16770 16098
rect 18062 16046 18114 16098
rect 19182 16046 19234 16098
rect 21310 16046 21362 16098
rect 22430 16046 22482 16098
rect 22990 16046 23042 16098
rect 26238 16046 26290 16098
rect 28030 16046 28082 16098
rect 37662 16046 37714 16098
rect 18174 15934 18226 15986
rect 22542 15934 22594 15986
rect 26574 15934 26626 15986
rect 19070 15822 19122 15874
rect 20190 15822 20242 15874
rect 28254 15822 28306 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 17390 15486 17442 15538
rect 17726 15486 17778 15538
rect 22654 15486 22706 15538
rect 24670 15486 24722 15538
rect 15598 15374 15650 15426
rect 18062 15374 18114 15426
rect 20078 15374 20130 15426
rect 26350 15374 26402 15426
rect 16270 15262 16322 15314
rect 18286 15262 18338 15314
rect 19294 15262 19346 15314
rect 25566 15262 25618 15314
rect 15934 15150 15986 15202
rect 22206 15150 22258 15202
rect 28478 15150 28530 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 21646 14702 21698 14754
rect 23998 14702 24050 14754
rect 15822 14590 15874 14642
rect 17950 14590 18002 14642
rect 18398 14590 18450 14642
rect 24670 14590 24722 14642
rect 15150 14478 15202 14530
rect 22430 14478 22482 14530
rect 23438 14478 23490 14530
rect 23998 14478 24050 14530
rect 21870 14366 21922 14418
rect 22766 14366 22818 14418
rect 23662 14366 23714 14418
rect 24558 14366 24610 14418
rect 21310 14254 21362 14306
rect 23886 14254 23938 14306
rect 24782 14254 24834 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 18286 13806 18338 13858
rect 20190 13806 20242 13858
rect 21086 13806 21138 13858
rect 22766 13806 22818 13858
rect 22990 13806 23042 13858
rect 18510 13694 18562 13746
rect 20750 13694 20802 13746
rect 20078 13470 20130 13522
rect 20414 13470 20466 13522
rect 20750 13470 20802 13522
rect 22654 13470 22706 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 21758 13134 21810 13186
rect 18174 13022 18226 13074
rect 20302 13022 20354 13074
rect 20750 13022 20802 13074
rect 21422 13022 21474 13074
rect 22766 13022 22818 13074
rect 23886 13022 23938 13074
rect 26014 13022 26066 13074
rect 17502 12910 17554 12962
rect 23102 12910 23154 12962
rect 21534 12798 21586 12850
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 18286 12350 18338 12402
rect 23774 12350 23826 12402
rect 18846 12238 18898 12290
rect 21198 12238 21250 12290
rect 18622 12126 18674 12178
rect 20526 12126 20578 12178
rect 23326 12014 23378 12066
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 26798 5182 26850 5234
rect 25790 5070 25842 5122
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 25230 4286 25282 4338
rect 26238 4062 26290 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 25566 3614 25618 3666
rect 20750 3502 20802 3554
rect 24558 3502 24610 3554
rect 19070 3278 19122 3330
rect 21758 3278 21810 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 16800 41200 16912 42000
rect 20160 41200 20272 42000
rect 20832 41200 20944 42000
rect 22176 41200 22288 42000
rect 24864 41200 24976 42000
rect 25536 41200 25648 42000
rect 27552 41200 27664 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 16828 38276 16884 41200
rect 16828 38210 16884 38220
rect 18060 38276 18116 38286
rect 18060 38182 18116 38220
rect 17052 38050 17108 38062
rect 17052 37998 17054 38050
rect 17106 37998 17108 38050
rect 1708 37378 1764 37390
rect 1708 37326 1710 37378
rect 1762 37326 1764 37378
rect 1708 37044 1764 37326
rect 1708 36978 1764 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 17052 31948 17108 37998
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20188 36708 20244 41200
rect 20860 37492 20916 41200
rect 22204 38276 22260 41200
rect 22428 38276 22484 38286
rect 22204 38274 22484 38276
rect 22204 38222 22430 38274
rect 22482 38222 22484 38274
rect 22204 38220 22484 38222
rect 22428 38210 22484 38220
rect 24892 38276 24948 41200
rect 24892 38210 24948 38220
rect 20860 37426 20916 37436
rect 21420 38050 21476 38062
rect 21420 37998 21422 38050
rect 21474 37998 21476 38050
rect 20188 36642 20244 36652
rect 21084 37266 21140 37278
rect 21084 37214 21086 37266
rect 21138 37214 21140 37266
rect 20300 36484 20356 36494
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20300 31948 20356 36428
rect 21084 31948 21140 37214
rect 21308 36484 21364 36494
rect 21308 36390 21364 36428
rect 16940 31892 17108 31948
rect 20188 31892 20356 31948
rect 20748 31892 21140 31948
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4172 27636 4228 27646
rect 1932 25618 1988 25630
rect 1932 25566 1934 25618
rect 1986 25566 1988 25618
rect 1932 24948 1988 25566
rect 1932 24882 1988 24892
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 1932 23538 1988 23548
rect 1932 22932 1988 22942
rect 1932 22838 1988 22876
rect 1932 20914 1988 20926
rect 1932 20862 1934 20914
rect 1986 20862 1988 20914
rect 1932 20244 1988 20862
rect 4172 20804 4228 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 14140 27188 14196 27198
rect 14140 27074 14196 27132
rect 16940 27188 16996 31892
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 17948 28642 18004 28654
rect 17948 28590 17950 28642
rect 18002 28590 18004 28642
rect 17388 28532 17444 28542
rect 17388 27188 17444 28476
rect 17948 28532 18004 28590
rect 17948 28466 18004 28476
rect 18508 28532 18564 28542
rect 18508 27858 18564 28476
rect 18620 28532 18676 28542
rect 18620 28530 19684 28532
rect 18620 28478 18622 28530
rect 18674 28478 19684 28530
rect 18620 28476 19684 28478
rect 18620 28466 18676 28476
rect 18508 27806 18510 27858
rect 18562 27806 18564 27858
rect 18508 27794 18564 27806
rect 19292 27748 19348 27758
rect 19292 27654 19348 27692
rect 19628 27298 19684 28476
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19628 27246 19630 27298
rect 19682 27246 19684 27298
rect 19628 27234 19684 27246
rect 16940 27186 17332 27188
rect 16940 27134 16942 27186
rect 16994 27134 17332 27186
rect 16940 27132 17332 27134
rect 16940 27122 16996 27132
rect 14140 27022 14142 27074
rect 14194 27022 14196 27074
rect 14140 27010 14196 27022
rect 14812 26962 14868 26974
rect 14812 26910 14814 26962
rect 14866 26910 14868 26962
rect 14812 26516 14868 26910
rect 17276 26908 17332 27132
rect 17444 27132 17556 27188
rect 17388 27094 17444 27132
rect 17276 26852 17444 26908
rect 14812 26450 14868 26460
rect 15708 26516 15764 26526
rect 15708 26422 15764 26460
rect 17388 26402 17444 26852
rect 17388 26350 17390 26402
rect 17442 26350 17444 26402
rect 17388 26338 17444 26350
rect 15820 26180 15876 26190
rect 15820 26086 15876 26124
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 13916 25618 13972 25630
rect 13916 25566 13918 25618
rect 13970 25566 13972 25618
rect 4284 25508 4340 25518
rect 4284 25414 4340 25452
rect 13916 25508 13972 25566
rect 13916 25442 13972 25452
rect 16828 25508 16884 25518
rect 17500 25508 17556 27132
rect 19740 26964 19796 26974
rect 19740 26870 19796 26908
rect 20076 26962 20132 26974
rect 20076 26910 20078 26962
rect 20130 26910 20132 26962
rect 17836 26852 17892 26862
rect 17836 26514 17892 26796
rect 20076 26852 20132 26910
rect 20076 26786 20132 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 17836 26462 17838 26514
rect 17890 26462 17892 26514
rect 17612 26292 17668 26302
rect 17612 26198 17668 26236
rect 17724 26180 17780 26190
rect 17724 26086 17780 26124
rect 17612 25508 17668 25518
rect 16828 25506 17668 25508
rect 16828 25454 16830 25506
rect 16882 25454 17614 25506
rect 17666 25454 17668 25506
rect 16828 25452 17668 25454
rect 16828 25442 16884 25452
rect 16044 25394 16100 25406
rect 16044 25342 16046 25394
rect 16098 25342 16100 25394
rect 15148 24948 15204 24958
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 15148 24052 15204 24892
rect 16044 24946 16100 25342
rect 16828 25284 16884 25294
rect 16884 25228 16996 25284
rect 16828 25218 16884 25228
rect 16044 24894 16046 24946
rect 16098 24894 16100 24946
rect 16044 24882 16100 24894
rect 15932 24834 15988 24846
rect 15932 24782 15934 24834
rect 15986 24782 15988 24834
rect 15932 24724 15988 24782
rect 15932 24658 15988 24668
rect 16492 24724 16548 24734
rect 14924 24050 15204 24052
rect 14924 23998 15150 24050
rect 15202 23998 15204 24050
rect 14924 23996 15204 23998
rect 4284 23940 4340 23950
rect 4284 23846 4340 23884
rect 11452 23940 11508 23950
rect 4284 23156 4340 23166
rect 4284 23062 4340 23100
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 11452 22372 11508 23884
rect 12012 23492 12068 23502
rect 12012 23156 12068 23436
rect 14140 23380 14196 23390
rect 14140 23266 14196 23324
rect 14140 23214 14142 23266
rect 14194 23214 14196 23266
rect 14140 23202 14196 23214
rect 12012 23042 12068 23100
rect 12012 22990 12014 23042
rect 12066 22990 12068 23042
rect 12012 22978 12068 22990
rect 14924 23154 14980 23996
rect 15148 23958 15204 23996
rect 16156 24498 16212 24510
rect 16156 24446 16158 24498
rect 16210 24446 16212 24498
rect 16156 24052 16212 24446
rect 16156 23986 16212 23996
rect 15820 23828 15876 23838
rect 15820 23826 16212 23828
rect 15820 23774 15822 23826
rect 15874 23774 16212 23826
rect 15820 23772 16212 23774
rect 15820 23762 15876 23772
rect 15596 23714 15652 23726
rect 15596 23662 15598 23714
rect 15650 23662 15652 23714
rect 15596 23492 15652 23662
rect 15596 23426 15652 23436
rect 15708 23714 15764 23726
rect 15708 23662 15710 23714
rect 15762 23662 15764 23714
rect 15484 23380 15540 23390
rect 15708 23380 15764 23662
rect 15708 23324 16100 23380
rect 15484 23286 15540 23324
rect 14924 23102 14926 23154
rect 14978 23102 14980 23154
rect 13804 22932 13860 22942
rect 13804 22594 13860 22876
rect 13804 22542 13806 22594
rect 13858 22542 13860 22594
rect 13804 22530 13860 22542
rect 11452 21474 11508 22316
rect 13580 22148 13636 22158
rect 13580 22054 13636 22092
rect 13692 22146 13748 22158
rect 13692 22094 13694 22146
rect 13746 22094 13748 22146
rect 13580 21700 13636 21710
rect 13692 21700 13748 22094
rect 14812 21812 14868 21822
rect 14924 21812 14980 23102
rect 15596 23268 15652 23278
rect 15036 22932 15092 22942
rect 15036 22596 15092 22876
rect 15260 22820 15316 22830
rect 15036 22540 15204 22596
rect 15036 22372 15092 22382
rect 15036 22278 15092 22316
rect 15148 22148 15204 22540
rect 13580 21698 13748 21700
rect 13580 21646 13582 21698
rect 13634 21646 13748 21698
rect 13580 21644 13748 21646
rect 14364 21810 14980 21812
rect 14364 21758 14814 21810
rect 14866 21758 14980 21810
rect 14364 21756 14980 21758
rect 15036 22092 15204 22148
rect 15260 22370 15316 22764
rect 15260 22318 15262 22370
rect 15314 22318 15316 22370
rect 13580 21634 13636 21644
rect 14364 21586 14420 21756
rect 14812 21746 14868 21756
rect 15036 21700 15092 22092
rect 15260 21924 15316 22318
rect 15484 22372 15540 22382
rect 15596 22372 15652 23212
rect 16044 23154 16100 23324
rect 16044 23102 16046 23154
rect 16098 23102 16100 23154
rect 16044 23090 16100 23102
rect 16156 23156 16212 23772
rect 16156 23062 16212 23100
rect 15820 23044 15876 23054
rect 15484 22370 15652 22372
rect 15484 22318 15486 22370
rect 15538 22318 15652 22370
rect 15484 22316 15652 22318
rect 15708 22372 15764 22382
rect 15820 22372 15876 22988
rect 16156 22820 16212 22830
rect 16156 22482 16212 22764
rect 16156 22430 16158 22482
rect 16210 22430 16212 22482
rect 16156 22418 16212 22430
rect 15708 22370 15876 22372
rect 15708 22318 15710 22370
rect 15762 22318 15876 22370
rect 15708 22316 15876 22318
rect 15484 22306 15540 22316
rect 15708 22306 15764 22316
rect 15372 22148 15428 22158
rect 15372 22054 15428 22092
rect 14364 21534 14366 21586
rect 14418 21534 14420 21586
rect 14364 21522 14420 21534
rect 14924 21644 15092 21700
rect 15148 21868 15316 21924
rect 11452 21422 11454 21474
rect 11506 21422 11508 21474
rect 11452 21410 11508 21422
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4172 20738 4228 20748
rect 4284 20802 4340 20814
rect 4284 20750 4286 20802
rect 4338 20750 4340 20802
rect 4284 20468 4340 20750
rect 4284 20402 4340 20412
rect 10892 20692 10948 20702
rect 1932 20178 1988 20188
rect 10892 19906 10948 20636
rect 14476 20692 14532 20702
rect 14476 20598 14532 20636
rect 14588 20578 14644 20590
rect 14588 20526 14590 20578
rect 14642 20526 14644 20578
rect 14588 20132 14644 20526
rect 14924 20188 14980 21644
rect 15148 21588 15204 21868
rect 14588 20066 14644 20076
rect 14700 20132 14980 20188
rect 15036 21532 15204 21588
rect 13804 20020 13860 20030
rect 13580 20018 14084 20020
rect 13580 19966 13806 20018
rect 13858 19966 14084 20018
rect 13580 19964 14084 19966
rect 13020 19908 13076 19918
rect 10892 19854 10894 19906
rect 10946 19854 10948 19906
rect 10892 19842 10948 19854
rect 12460 19906 13076 19908
rect 12460 19854 13022 19906
rect 13074 19854 13076 19906
rect 12460 19852 13076 19854
rect 12236 19796 12292 19806
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 12236 19234 12292 19740
rect 12236 19182 12238 19234
rect 12290 19182 12292 19234
rect 12236 19170 12292 19182
rect 12460 19122 12516 19852
rect 13020 19842 13076 19852
rect 12460 19070 12462 19122
rect 12514 19070 12516 19122
rect 12460 19058 12516 19070
rect 4284 18452 4340 18462
rect 13580 18452 13636 19964
rect 13804 19954 13860 19964
rect 14028 19346 14084 19964
rect 14476 19908 14532 19918
rect 14700 19908 14756 20132
rect 14476 19814 14532 19852
rect 14588 19906 14756 19908
rect 14588 19854 14702 19906
rect 14754 19854 14756 19906
rect 14588 19852 14756 19854
rect 14140 19796 14196 19806
rect 14140 19702 14196 19740
rect 14028 19294 14030 19346
rect 14082 19294 14084 19346
rect 14028 19282 14084 19294
rect 4284 18358 4340 18396
rect 13468 18396 13580 18452
rect 10668 18340 10724 18350
rect 12796 18340 12852 18350
rect 1932 18228 1988 18238
rect 1932 18134 1988 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 10668 17780 10724 18284
rect 12460 18338 12852 18340
rect 12460 18286 12798 18338
rect 12850 18286 12852 18338
rect 12460 18284 12852 18286
rect 10668 17714 10724 17724
rect 12236 18228 12292 18238
rect 12236 17666 12292 18172
rect 12236 17614 12238 17666
rect 12290 17614 12292 17666
rect 12236 17602 12292 17614
rect 12460 17554 12516 18284
rect 12796 18274 12852 18284
rect 12460 17502 12462 17554
rect 12514 17502 12516 17554
rect 12460 17490 12516 17502
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 13468 16098 13524 18396
rect 13580 18358 13636 18396
rect 14476 19012 14532 19022
rect 14476 18450 14532 18956
rect 14476 18398 14478 18450
rect 14530 18398 14532 18450
rect 14476 18386 14532 18398
rect 14588 18452 14644 19852
rect 14700 19842 14756 19852
rect 14812 19234 14868 19246
rect 14812 19182 14814 19234
rect 14866 19182 14868 19234
rect 14700 18452 14756 18462
rect 14588 18450 14756 18452
rect 14588 18398 14702 18450
rect 14754 18398 14756 18450
rect 14588 18396 14756 18398
rect 14700 18386 14756 18396
rect 13804 18228 13860 18238
rect 13804 18134 13860 18172
rect 14252 18226 14308 18238
rect 14252 18174 14254 18226
rect 14306 18174 14308 18226
rect 13804 17892 13860 17902
rect 13804 17798 13860 17836
rect 14140 17892 14196 17902
rect 14252 17892 14308 18174
rect 14140 17890 14308 17892
rect 14140 17838 14142 17890
rect 14194 17838 14308 17890
rect 14140 17836 14308 17838
rect 14812 17892 14868 19182
rect 15036 19122 15092 21532
rect 16492 20692 16548 24668
rect 16828 24052 16884 24062
rect 16828 23958 16884 23996
rect 16828 23828 16884 23838
rect 16940 23828 16996 25228
rect 17500 24948 17556 24958
rect 17612 24948 17668 25452
rect 17500 24946 17612 24948
rect 17500 24894 17502 24946
rect 17554 24894 17612 24946
rect 17500 24892 17612 24894
rect 17500 24882 17556 24892
rect 17612 24882 17668 24892
rect 17836 24722 17892 26462
rect 17836 24670 17838 24722
rect 17890 24670 17892 24722
rect 17724 23938 17780 23950
rect 17724 23886 17726 23938
rect 17778 23886 17780 23938
rect 16828 23826 16996 23828
rect 16828 23774 16830 23826
rect 16882 23774 16996 23826
rect 16828 23772 16996 23774
rect 17276 23826 17332 23838
rect 17276 23774 17278 23826
rect 17330 23774 17332 23826
rect 16828 23762 16884 23772
rect 16716 23714 16772 23726
rect 16716 23662 16718 23714
rect 16770 23662 16772 23714
rect 16604 23154 16660 23166
rect 16604 23102 16606 23154
rect 16658 23102 16660 23154
rect 16604 21140 16660 23102
rect 16716 22372 16772 23662
rect 17052 23714 17108 23726
rect 17052 23662 17054 23714
rect 17106 23662 17108 23714
rect 17052 23380 17108 23662
rect 17164 23380 17220 23390
rect 17052 23324 17164 23380
rect 16828 23156 16884 23166
rect 16828 22482 16884 23100
rect 16828 22430 16830 22482
rect 16882 22430 16884 22482
rect 16828 22418 16884 22430
rect 17164 22372 17220 23324
rect 17276 23156 17332 23774
rect 17276 23090 17332 23100
rect 17612 23268 17668 23278
rect 17388 22932 17444 22942
rect 17388 22838 17444 22876
rect 17164 22316 17332 22372
rect 16716 22278 16772 22316
rect 16940 22148 16996 22158
rect 16940 22146 17108 22148
rect 16940 22094 16942 22146
rect 16994 22094 17108 22146
rect 16940 22092 17108 22094
rect 16940 22082 16996 22092
rect 16604 21084 16996 21140
rect 15708 20690 16548 20692
rect 15708 20638 16494 20690
rect 16546 20638 16548 20690
rect 15708 20636 16548 20638
rect 15708 20242 15764 20636
rect 16492 20626 16548 20636
rect 16716 20802 16772 20814
rect 16716 20750 16718 20802
rect 16770 20750 16772 20802
rect 15708 20190 15710 20242
rect 15762 20190 15764 20242
rect 15484 20132 15540 20142
rect 15484 20038 15540 20076
rect 15372 20020 15428 20030
rect 15372 19926 15428 19964
rect 15596 19908 15652 19918
rect 15596 19814 15652 19852
rect 15708 19684 15764 20190
rect 15932 20020 15988 20030
rect 16268 20020 16324 20030
rect 15932 20018 16324 20020
rect 15932 19966 15934 20018
rect 15986 19966 16270 20018
rect 16322 19966 16324 20018
rect 15932 19964 16324 19966
rect 15932 19954 15988 19964
rect 16268 19796 16324 19964
rect 16492 20020 16548 20030
rect 16716 20020 16772 20750
rect 16492 20018 16772 20020
rect 16492 19966 16494 20018
rect 16546 19966 16772 20018
rect 16492 19964 16772 19966
rect 16828 20018 16884 20030
rect 16828 19966 16830 20018
rect 16882 19966 16884 20018
rect 16268 19730 16324 19740
rect 16380 19906 16436 19918
rect 16380 19854 16382 19906
rect 16434 19854 16436 19906
rect 15036 19070 15038 19122
rect 15090 19070 15092 19122
rect 15036 19058 15092 19070
rect 15372 19628 15764 19684
rect 15148 18452 15204 18462
rect 14140 17826 14196 17836
rect 14812 17826 14868 17836
rect 15036 18396 15148 18452
rect 13580 17780 13636 17790
rect 13580 17686 13636 17724
rect 15036 16884 15092 18396
rect 15148 18358 15204 18396
rect 15372 17668 15428 19628
rect 15484 19236 15540 19246
rect 15484 19234 16100 19236
rect 15484 19182 15486 19234
rect 15538 19182 16100 19234
rect 15484 19180 16100 19182
rect 15484 19170 15540 19180
rect 15708 19010 15764 19022
rect 15708 18958 15710 19010
rect 15762 18958 15764 19010
rect 15708 18900 15764 18958
rect 15708 18834 15764 18844
rect 16044 18452 16100 19180
rect 16268 19124 16324 19134
rect 16156 19068 16268 19124
rect 16156 18674 16212 19068
rect 16268 19058 16324 19068
rect 16380 19012 16436 19854
rect 16492 19236 16548 19964
rect 16492 19142 16548 19180
rect 16380 18946 16436 18956
rect 16156 18622 16158 18674
rect 16210 18622 16212 18674
rect 16156 18610 16212 18622
rect 16828 18564 16884 19966
rect 16940 19012 16996 21084
rect 17052 19908 17108 22092
rect 17164 22146 17220 22158
rect 17164 22094 17166 22146
rect 17218 22094 17220 22146
rect 17164 20020 17220 22094
rect 17164 19954 17220 19964
rect 17052 19842 17108 19852
rect 17276 19122 17332 22316
rect 17612 22258 17668 23212
rect 17612 22206 17614 22258
rect 17666 22206 17668 22258
rect 17612 22194 17668 22206
rect 17724 22820 17780 23886
rect 17836 23714 17892 24670
rect 17836 23662 17838 23714
rect 17890 23662 17892 23714
rect 17836 23650 17892 23662
rect 17948 26290 18004 26302
rect 17948 26238 17950 26290
rect 18002 26238 18004 26290
rect 17948 23380 18004 26238
rect 18732 26292 18788 26302
rect 18284 25396 18340 25406
rect 18732 25396 18788 26236
rect 20188 25620 20244 31892
rect 20748 28756 20804 31892
rect 20524 28754 20804 28756
rect 20524 28702 20750 28754
rect 20802 28702 20804 28754
rect 20524 28700 20804 28702
rect 20524 27074 20580 28700
rect 20748 28690 20804 28700
rect 21084 29314 21140 29326
rect 21084 29262 21086 29314
rect 21138 29262 21140 29314
rect 21084 28644 21140 29262
rect 21084 28578 21140 28588
rect 21308 27748 21364 27758
rect 21308 27298 21364 27692
rect 21420 27748 21476 37998
rect 25228 38050 25284 38062
rect 25228 37998 25230 38050
rect 25282 37998 25284 38050
rect 22092 37492 22148 37502
rect 22092 37398 22148 37436
rect 22316 36708 22372 36718
rect 22316 36614 22372 36652
rect 21644 28644 21700 28654
rect 22092 28644 22148 28654
rect 21700 28588 21924 28644
rect 21644 28550 21700 28588
rect 21868 27858 21924 28588
rect 22092 28550 22148 28588
rect 25228 28532 25284 37998
rect 25564 37492 25620 41200
rect 27580 38610 27636 41200
rect 27580 38558 27582 38610
rect 27634 38558 27636 38610
rect 27580 38546 27636 38558
rect 28364 38610 28420 38622
rect 28364 38558 28366 38610
rect 28418 38558 28420 38610
rect 26124 38276 26180 38286
rect 26124 38182 26180 38220
rect 28364 37938 28420 38558
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 28364 37886 28366 37938
rect 28418 37886 28420 37938
rect 28364 37874 28420 37886
rect 25564 37426 25620 37436
rect 26796 37492 26852 37502
rect 26796 37398 26852 37436
rect 21868 27806 21870 27858
rect 21922 27806 21924 27858
rect 21868 27794 21924 27806
rect 24668 28476 25284 28532
rect 26012 37266 26068 37278
rect 26012 37214 26014 37266
rect 26066 37214 26068 37266
rect 22540 27748 22596 27758
rect 21420 27746 21700 27748
rect 21420 27694 21422 27746
rect 21474 27694 21700 27746
rect 21420 27692 21700 27694
rect 21420 27682 21476 27692
rect 21308 27246 21310 27298
rect 21362 27246 21364 27298
rect 21308 27234 21364 27246
rect 20524 27022 20526 27074
rect 20578 27022 20580 27074
rect 20524 27010 20580 27022
rect 20748 27074 20804 27086
rect 20748 27022 20750 27074
rect 20802 27022 20804 27074
rect 20412 26964 20468 26974
rect 20412 26870 20468 26908
rect 20748 26964 20804 27022
rect 20748 26898 20804 26908
rect 21308 26964 21364 26974
rect 20300 26850 20356 26862
rect 20300 26798 20302 26850
rect 20354 26798 20356 26850
rect 20300 26628 20356 26798
rect 20300 26562 20356 26572
rect 20748 26628 20804 26638
rect 20524 26516 20580 26526
rect 20412 25620 20468 25630
rect 20188 25618 20468 25620
rect 20188 25566 20414 25618
rect 20466 25566 20468 25618
rect 20188 25564 20468 25566
rect 18284 25394 18452 25396
rect 18284 25342 18286 25394
rect 18338 25342 18452 25394
rect 18284 25340 18452 25342
rect 18284 25330 18340 25340
rect 18396 24948 18452 25340
rect 18620 24948 18676 24958
rect 18396 24946 18676 24948
rect 18396 24894 18622 24946
rect 18674 24894 18676 24946
rect 18396 24892 18676 24894
rect 18620 24882 18676 24892
rect 18060 24724 18116 24734
rect 18060 24630 18116 24668
rect 18396 24724 18452 24734
rect 18620 24724 18676 24734
rect 18396 24722 18564 24724
rect 18396 24670 18398 24722
rect 18450 24670 18564 24722
rect 18396 24668 18564 24670
rect 18396 24658 18452 24668
rect 18508 24612 18564 24668
rect 18620 24630 18676 24668
rect 17836 23324 18004 23380
rect 18172 23938 18228 23950
rect 18172 23886 18174 23938
rect 18226 23886 18228 23938
rect 17836 23266 17892 23324
rect 17836 23214 17838 23266
rect 17890 23214 17892 23266
rect 17836 23044 17892 23214
rect 18172 23268 18228 23886
rect 17836 22978 17892 22988
rect 17948 23154 18004 23166
rect 17948 23102 17950 23154
rect 18002 23102 18004 23154
rect 17948 22820 18004 23102
rect 18172 23154 18228 23212
rect 18172 23102 18174 23154
rect 18226 23102 18228 23154
rect 18172 23090 18228 23102
rect 17724 22764 18004 22820
rect 18060 23044 18116 23054
rect 17612 21252 17668 21262
rect 17612 20580 17668 21196
rect 17612 20018 17668 20524
rect 17612 19966 17614 20018
rect 17666 19966 17668 20018
rect 17500 19796 17556 19806
rect 17276 19070 17278 19122
rect 17330 19070 17332 19122
rect 17164 19012 17220 19022
rect 16940 19010 17220 19012
rect 16940 18958 17166 19010
rect 17218 18958 17220 19010
rect 16940 18956 17220 18958
rect 17164 18946 17220 18956
rect 17276 18676 17332 19070
rect 17388 19234 17444 19246
rect 17388 19182 17390 19234
rect 17442 19182 17444 19234
rect 17388 19124 17444 19182
rect 17388 19058 17444 19068
rect 17276 18610 17332 18620
rect 15932 18450 16100 18452
rect 15932 18398 16046 18450
rect 16098 18398 16100 18450
rect 15932 18396 16100 18398
rect 15484 17668 15540 17678
rect 15372 17666 15540 17668
rect 15372 17614 15486 17666
rect 15538 17614 15540 17666
rect 15372 17612 15540 17614
rect 15484 17602 15540 17612
rect 15596 17442 15652 17454
rect 15596 17390 15598 17442
rect 15650 17390 15652 17442
rect 14252 16212 14308 16222
rect 14252 16118 14308 16156
rect 13468 16046 13470 16098
rect 13522 16046 13524 16098
rect 13468 16034 13524 16046
rect 15036 15204 15092 16828
rect 15484 16996 15540 17006
rect 15596 16996 15652 17390
rect 15484 16994 15652 16996
rect 15484 16942 15486 16994
rect 15538 16942 15652 16994
rect 15484 16940 15652 16942
rect 15820 17442 15876 17454
rect 15820 17390 15822 17442
rect 15874 17390 15876 17442
rect 15820 16996 15876 17390
rect 15484 16212 15540 16940
rect 15820 16930 15876 16940
rect 15708 16884 15764 16894
rect 15484 16146 15540 16156
rect 15596 16882 15764 16884
rect 15596 16830 15710 16882
rect 15762 16830 15764 16882
rect 15596 16828 15764 16830
rect 15596 15426 15652 16828
rect 15708 16818 15764 16828
rect 15932 16212 15988 18396
rect 16044 18386 16100 18396
rect 16492 18450 16548 18462
rect 16492 18398 16494 18450
rect 16546 18398 16548 18450
rect 16044 17892 16100 17902
rect 16044 17798 16100 17836
rect 16044 17668 16100 17678
rect 16044 17574 16100 17612
rect 16380 17554 16436 17566
rect 16380 17502 16382 17554
rect 16434 17502 16436 17554
rect 16380 17108 16436 17502
rect 16492 17220 16548 18398
rect 16828 17892 16884 18508
rect 17500 18450 17556 19740
rect 17500 18398 17502 18450
rect 17554 18398 17556 18450
rect 17500 18386 17556 18398
rect 17164 17892 17220 17902
rect 16828 17890 17220 17892
rect 16828 17838 17166 17890
rect 17218 17838 17220 17890
rect 16828 17836 17220 17838
rect 17164 17826 17220 17836
rect 17500 17778 17556 17790
rect 17500 17726 17502 17778
rect 17554 17726 17556 17778
rect 17052 17668 17108 17678
rect 17052 17574 17108 17612
rect 16492 17154 16548 17164
rect 16604 17444 16660 17454
rect 16380 17042 16436 17052
rect 16492 16996 16548 17006
rect 16604 16996 16660 17388
rect 17500 17108 17556 17726
rect 17500 17042 17556 17052
rect 16492 16994 16660 16996
rect 16492 16942 16494 16994
rect 16546 16942 16660 16994
rect 16492 16940 16660 16942
rect 16492 16930 16548 16940
rect 16268 16884 16324 16894
rect 17612 16884 17668 19966
rect 17724 19908 17780 22764
rect 17948 22146 18004 22158
rect 17948 22094 17950 22146
rect 18002 22094 18004 22146
rect 17948 21252 18004 22094
rect 17948 21186 18004 21196
rect 17948 21028 18004 21038
rect 18060 21028 18116 22988
rect 17948 21026 18116 21028
rect 17948 20974 17950 21026
rect 18002 20974 18116 21026
rect 17948 20972 18116 20974
rect 17948 20962 18004 20972
rect 18172 20802 18228 20814
rect 18172 20750 18174 20802
rect 18226 20750 18228 20802
rect 18060 20020 18116 20030
rect 18172 20020 18228 20750
rect 18060 20018 18228 20020
rect 18060 19966 18062 20018
rect 18114 19966 18228 20018
rect 18060 19964 18228 19966
rect 17836 19908 17892 19918
rect 17724 19852 17836 19908
rect 17836 19234 17892 19852
rect 17836 19182 17838 19234
rect 17890 19182 17892 19234
rect 17836 18900 17892 19182
rect 17836 18834 17892 18844
rect 18060 19908 18116 19964
rect 18060 17668 18116 19852
rect 18508 19796 18564 24556
rect 18732 24610 18788 25340
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 18732 24558 18734 24610
rect 18786 24558 18788 24610
rect 18732 24546 18788 24558
rect 19180 24612 19236 24622
rect 19180 24610 20020 24612
rect 19180 24558 19182 24610
rect 19234 24558 20020 24610
rect 19180 24556 20020 24558
rect 19180 24546 19236 24556
rect 19964 24162 20020 24556
rect 19964 24110 19966 24162
rect 20018 24110 20020 24162
rect 19964 24098 20020 24110
rect 20076 24052 20132 24062
rect 20412 24052 20468 25564
rect 20076 24050 20468 24052
rect 20076 23998 20078 24050
rect 20130 23998 20468 24050
rect 20076 23996 20468 23998
rect 20524 24724 20580 26460
rect 20076 23986 20132 23996
rect 20524 23940 20580 24668
rect 20188 23884 20580 23940
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 18620 23156 18676 23166
rect 18620 22258 18676 23100
rect 20076 22596 20132 22606
rect 20188 22596 20244 23884
rect 20748 23492 20804 26572
rect 21308 26292 21364 26908
rect 21420 26964 21476 26974
rect 21420 26962 21588 26964
rect 21420 26910 21422 26962
rect 21474 26910 21588 26962
rect 21420 26908 21588 26910
rect 21420 26898 21476 26908
rect 21420 26292 21476 26302
rect 21308 26290 21476 26292
rect 21308 26238 21422 26290
rect 21474 26238 21476 26290
rect 21308 26236 21476 26238
rect 21420 26226 21476 26236
rect 21532 26178 21588 26908
rect 21644 26514 21700 27692
rect 22540 27746 23268 27748
rect 22540 27694 22542 27746
rect 22594 27694 23268 27746
rect 22540 27692 23268 27694
rect 22540 27682 22596 27692
rect 22204 27074 22260 27086
rect 22204 27022 22206 27074
rect 22258 27022 22260 27074
rect 21644 26462 21646 26514
rect 21698 26462 21700 26514
rect 21644 26450 21700 26462
rect 21868 26628 21924 26638
rect 21868 26514 21924 26572
rect 21868 26462 21870 26514
rect 21922 26462 21924 26514
rect 21868 26450 21924 26462
rect 22204 26516 22260 27022
rect 22540 27076 22596 27086
rect 23100 27076 23156 27086
rect 22540 26982 22596 27020
rect 22988 27074 23156 27076
rect 22988 27022 23102 27074
rect 23154 27022 23156 27074
rect 22988 27020 23156 27022
rect 22652 26964 22708 26974
rect 22652 26870 22708 26908
rect 22204 26450 22260 26460
rect 22316 26850 22372 26862
rect 22316 26798 22318 26850
rect 22370 26798 22372 26850
rect 21532 26126 21534 26178
rect 21586 26126 21588 26178
rect 21532 26114 21588 26126
rect 21980 26292 22036 26302
rect 22316 26292 22372 26798
rect 22428 26850 22484 26862
rect 22428 26798 22430 26850
rect 22482 26798 22484 26850
rect 22428 26404 22484 26798
rect 22428 26338 22484 26348
rect 22988 26292 23044 27020
rect 23100 27010 23156 27020
rect 23100 26404 23156 26414
rect 23100 26310 23156 26348
rect 21980 26290 22372 26292
rect 21980 26238 21982 26290
rect 22034 26238 22372 26290
rect 21980 26236 22372 26238
rect 22764 26236 23044 26292
rect 21420 25282 21476 25294
rect 21420 25230 21422 25282
rect 21474 25230 21476 25282
rect 21420 24948 21476 25230
rect 21420 24052 21476 24892
rect 21868 24612 21924 24622
rect 21980 24612 22036 26236
rect 22652 26180 22708 26190
rect 22764 26180 22820 26236
rect 22652 26178 22820 26180
rect 22652 26126 22654 26178
rect 22706 26126 22820 26178
rect 22652 26124 22820 26126
rect 21924 24556 22036 24612
rect 22092 24612 22148 24622
rect 21868 24546 21924 24556
rect 21644 24052 21700 24062
rect 22092 24052 22148 24556
rect 22652 24612 22708 26124
rect 22988 26068 23044 26078
rect 23212 26068 23268 27692
rect 24668 27746 24724 28476
rect 24668 27694 24670 27746
rect 24722 27694 24724 27746
rect 24668 27076 24724 27694
rect 24668 27010 24724 27020
rect 26012 27186 26068 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 26012 27134 26014 27186
rect 26066 27134 26068 27186
rect 22988 26066 23268 26068
rect 22988 26014 22990 26066
rect 23042 26014 23268 26066
rect 22988 26012 23268 26014
rect 23324 26964 23380 26974
rect 22988 26002 23044 26012
rect 22652 24518 22708 24556
rect 21420 24050 22148 24052
rect 21420 23998 21646 24050
rect 21698 23998 22148 24050
rect 21420 23996 22148 23998
rect 21644 23986 21700 23996
rect 22092 23938 22148 23996
rect 22092 23886 22094 23938
rect 22146 23886 22148 23938
rect 22092 23874 22148 23886
rect 22316 24388 22372 24398
rect 20748 23436 21588 23492
rect 20748 23268 20804 23436
rect 20636 23266 20804 23268
rect 20636 23214 20750 23266
rect 20802 23214 20804 23266
rect 20636 23212 20804 23214
rect 20524 23044 20580 23054
rect 20524 22950 20580 22988
rect 20076 22594 20244 22596
rect 20076 22542 20078 22594
rect 20130 22542 20244 22594
rect 20076 22540 20244 22542
rect 20076 22530 20132 22540
rect 18620 22206 18622 22258
rect 18674 22206 18676 22258
rect 18620 22194 18676 22206
rect 19180 22372 19236 22382
rect 18956 22146 19012 22158
rect 18956 22094 18958 22146
rect 19010 22094 19012 22146
rect 18620 20916 18676 20926
rect 18620 20802 18676 20860
rect 18620 20750 18622 20802
rect 18674 20750 18676 20802
rect 18620 20132 18676 20750
rect 18956 20690 19012 22094
rect 19180 21810 19236 22316
rect 20076 22372 20132 22382
rect 20076 22278 20132 22316
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19180 21758 19182 21810
rect 19234 21758 19236 21810
rect 19180 21746 19236 21758
rect 20188 21698 20244 22540
rect 20188 21646 20190 21698
rect 20242 21646 20244 21698
rect 20188 21634 20244 21646
rect 20300 22370 20356 22382
rect 20300 22318 20302 22370
rect 20354 22318 20356 22370
rect 19292 21588 19348 21598
rect 19292 20802 19348 21532
rect 19516 21586 19572 21598
rect 19516 21534 19518 21586
rect 19570 21534 19572 21586
rect 19516 20916 19572 21534
rect 19852 21588 19908 21626
rect 19852 21522 19908 21532
rect 19852 21364 19908 21374
rect 19516 20850 19572 20860
rect 19628 21362 19908 21364
rect 19628 21310 19854 21362
rect 19906 21310 19908 21362
rect 19628 21308 19908 21310
rect 19292 20750 19294 20802
rect 19346 20750 19348 20802
rect 19292 20738 19348 20750
rect 18956 20638 18958 20690
rect 19010 20638 19012 20690
rect 18620 20076 18900 20132
rect 18844 19796 18900 20076
rect 18956 20020 19012 20638
rect 19068 20580 19124 20590
rect 19068 20486 19124 20524
rect 19180 20020 19236 20030
rect 18956 20018 19348 20020
rect 18956 19966 19182 20018
rect 19234 19966 19348 20018
rect 18956 19964 19348 19966
rect 19180 19954 19236 19964
rect 18956 19796 19012 19806
rect 18844 19794 19012 19796
rect 18844 19742 18958 19794
rect 19010 19742 19012 19794
rect 18844 19740 19012 19742
rect 18508 19730 18564 19740
rect 18956 19572 19012 19740
rect 18956 19516 19236 19572
rect 18172 19348 18228 19358
rect 18172 19122 18228 19292
rect 18172 19070 18174 19122
rect 18226 19070 18228 19122
rect 18172 19058 18228 19070
rect 18732 19236 18788 19246
rect 18732 19122 18788 19180
rect 18732 19070 18734 19122
rect 18786 19070 18788 19122
rect 18508 18564 18564 18574
rect 18508 18470 18564 18508
rect 18732 18450 18788 19070
rect 18732 18398 18734 18450
rect 18786 18398 18788 18450
rect 18732 18386 18788 18398
rect 19068 18340 19124 18350
rect 18844 18338 19124 18340
rect 18844 18286 19070 18338
rect 19122 18286 19124 18338
rect 18844 18284 19124 18286
rect 18396 17778 18452 17790
rect 18396 17726 18398 17778
rect 18450 17726 18452 17778
rect 18060 17602 18116 17612
rect 18284 17668 18340 17678
rect 18284 17574 18340 17612
rect 17948 17220 18004 17230
rect 17948 17108 18004 17164
rect 17836 17106 18004 17108
rect 17836 17054 17950 17106
rect 18002 17054 18004 17106
rect 17836 17052 18004 17054
rect 16268 16882 16436 16884
rect 16268 16830 16270 16882
rect 16322 16830 16436 16882
rect 16268 16828 16436 16830
rect 16268 16818 16324 16828
rect 15596 15374 15598 15426
rect 15650 15374 15652 15426
rect 15596 15362 15652 15374
rect 15820 15988 15876 15998
rect 15036 15148 15204 15204
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 15148 14530 15204 15148
rect 15820 14642 15876 15932
rect 15932 15202 15988 16156
rect 16380 16212 16436 16828
rect 17500 16828 17668 16884
rect 17724 16884 17780 16894
rect 17164 16212 17220 16222
rect 16380 16210 16772 16212
rect 16380 16158 16382 16210
rect 16434 16158 16772 16210
rect 16380 16156 16772 16158
rect 16380 16146 16436 16156
rect 16716 16098 16772 16156
rect 17164 16118 17220 16156
rect 16716 16046 16718 16098
rect 16770 16046 16772 16098
rect 16716 16034 16772 16046
rect 17388 15988 17444 15998
rect 17388 15538 17444 15932
rect 17388 15486 17390 15538
rect 17442 15486 17444 15538
rect 17388 15474 17444 15486
rect 16268 15316 16324 15326
rect 16268 15222 16324 15260
rect 17500 15316 17556 16828
rect 17724 16212 17780 16828
rect 17500 15250 17556 15260
rect 17612 16210 17780 16212
rect 17612 16158 17726 16210
rect 17778 16158 17780 16210
rect 17612 16156 17780 16158
rect 15932 15150 15934 15202
rect 15986 15150 15988 15202
rect 15932 15138 15988 15150
rect 17612 15148 17668 16156
rect 17724 16146 17780 16156
rect 17724 15540 17780 15550
rect 17836 15540 17892 17052
rect 17948 17042 18004 17052
rect 18060 16884 18116 16894
rect 18060 16882 18228 16884
rect 18060 16830 18062 16882
rect 18114 16830 18228 16882
rect 18060 16828 18228 16830
rect 18060 16818 18116 16828
rect 18060 16212 18116 16222
rect 18060 16098 18116 16156
rect 18060 16046 18062 16098
rect 18114 16046 18116 16098
rect 18060 16034 18116 16046
rect 17724 15538 17892 15540
rect 17724 15486 17726 15538
rect 17778 15486 17892 15538
rect 17724 15484 17892 15486
rect 18172 15986 18228 16828
rect 18172 15934 18174 15986
rect 18226 15934 18228 15986
rect 17724 15474 17780 15484
rect 18060 15426 18116 15438
rect 18060 15374 18062 15426
rect 18114 15374 18116 15426
rect 18060 15316 18116 15374
rect 18060 15250 18116 15260
rect 18172 15316 18228 15934
rect 18396 15988 18452 17726
rect 18396 15922 18452 15932
rect 18284 15316 18340 15326
rect 18172 15314 18340 15316
rect 18172 15262 18286 15314
rect 18338 15262 18340 15314
rect 18172 15260 18340 15262
rect 17612 15092 17780 15148
rect 17724 14644 17780 15092
rect 15820 14590 15822 14642
rect 15874 14590 15876 14642
rect 15820 14578 15876 14590
rect 17500 14588 17724 14644
rect 15148 14478 15150 14530
rect 15202 14478 15204 14530
rect 15148 14466 15204 14478
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 17500 12962 17556 14588
rect 17724 14578 17780 14588
rect 17948 14644 18004 14654
rect 18172 14644 18228 15260
rect 18284 15250 18340 15260
rect 18508 15204 18564 15214
rect 17948 14642 18228 14644
rect 17948 14590 17950 14642
rect 18002 14590 18228 14642
rect 17948 14588 18228 14590
rect 18396 15092 18564 15148
rect 18396 14644 18452 15092
rect 17948 14578 18004 14588
rect 18396 14550 18452 14588
rect 18284 13858 18340 13870
rect 18284 13806 18286 13858
rect 18338 13806 18340 13858
rect 18172 13076 18228 13086
rect 18284 13076 18340 13806
rect 18508 13748 18564 13758
rect 18172 13074 18340 13076
rect 18172 13022 18174 13074
rect 18226 13022 18340 13074
rect 18172 13020 18340 13022
rect 18396 13746 18564 13748
rect 18396 13694 18510 13746
rect 18562 13694 18564 13746
rect 18396 13692 18564 13694
rect 18172 13010 18228 13020
rect 17500 12910 17502 12962
rect 17554 12910 17556 12962
rect 17500 12898 17556 12910
rect 18284 12404 18340 12414
rect 18396 12404 18452 13692
rect 18508 13682 18564 13692
rect 18284 12402 18452 12404
rect 18284 12350 18286 12402
rect 18338 12350 18452 12402
rect 18284 12348 18452 12350
rect 18620 13524 18676 13534
rect 18284 12338 18340 12348
rect 18620 12178 18676 13468
rect 18844 12290 18900 18284
rect 19068 18274 19124 18284
rect 19180 18228 19236 19516
rect 19180 18162 19236 18172
rect 19068 17666 19124 17678
rect 19068 17614 19070 17666
rect 19122 17614 19124 17666
rect 19068 17220 19124 17614
rect 19180 17444 19236 17454
rect 19292 17444 19348 19964
rect 19516 20018 19572 20030
rect 19516 19966 19518 20018
rect 19570 19966 19572 20018
rect 19404 19348 19460 19358
rect 19404 18450 19460 19292
rect 19516 19124 19572 19966
rect 19516 18562 19572 19068
rect 19516 18510 19518 18562
rect 19570 18510 19572 18562
rect 19516 18498 19572 18510
rect 19404 18398 19406 18450
rect 19458 18398 19460 18450
rect 19404 18386 19460 18398
rect 19516 18340 19572 18350
rect 19516 17890 19572 18284
rect 19516 17838 19518 17890
rect 19570 17838 19572 17890
rect 19516 17826 19572 17838
rect 19516 17668 19572 17678
rect 19516 17574 19572 17612
rect 19236 17388 19348 17444
rect 19180 17378 19236 17388
rect 19068 17154 19124 17164
rect 18956 17108 19012 17118
rect 19628 17108 19684 21308
rect 19852 21298 19908 21308
rect 20300 21028 20356 22318
rect 20524 21812 20580 21822
rect 20636 21812 20692 23212
rect 20748 23202 20804 23212
rect 21196 23268 21252 23278
rect 21196 23174 21252 23212
rect 21532 23266 21588 23436
rect 21532 23214 21534 23266
rect 21586 23214 21588 23266
rect 21532 23202 21588 23214
rect 21980 23380 22036 23390
rect 20972 23156 21028 23166
rect 20972 23062 21028 23100
rect 21308 23156 21364 23166
rect 21308 23062 21364 23100
rect 21868 23154 21924 23166
rect 21868 23102 21870 23154
rect 21922 23102 21924 23154
rect 21868 22596 21924 23102
rect 21980 23154 22036 23324
rect 22316 23378 22372 24332
rect 22316 23326 22318 23378
rect 22370 23326 22372 23378
rect 22316 23314 22372 23326
rect 22764 23826 22820 23838
rect 22764 23774 22766 23826
rect 22818 23774 22820 23826
rect 22764 23380 22820 23774
rect 22764 23314 22820 23324
rect 23100 23492 23156 23502
rect 23100 23378 23156 23436
rect 23100 23326 23102 23378
rect 23154 23326 23156 23378
rect 23100 23314 23156 23326
rect 22652 23268 22708 23278
rect 22652 23174 22708 23212
rect 21980 23102 21982 23154
rect 22034 23102 22036 23154
rect 21980 23090 22036 23102
rect 22316 23154 22372 23166
rect 22876 23156 22932 23166
rect 23324 23156 23380 26908
rect 23884 26964 23940 26974
rect 23884 26962 24500 26964
rect 23884 26910 23886 26962
rect 23938 26910 24500 26962
rect 23884 26908 24500 26910
rect 23884 26898 23940 26908
rect 23436 26740 23492 26750
rect 23436 26402 23492 26684
rect 23660 26516 23716 26526
rect 23660 26422 23716 26460
rect 23884 26516 23940 26526
rect 23884 26422 23940 26460
rect 23996 26460 24388 26516
rect 23436 26350 23438 26402
rect 23490 26350 23492 26402
rect 23436 26338 23492 26350
rect 23996 26178 24052 26460
rect 24108 26292 24164 26302
rect 24332 26292 24388 26460
rect 24444 26514 24500 26908
rect 24444 26462 24446 26514
rect 24498 26462 24500 26514
rect 24444 26450 24500 26462
rect 26012 26516 26068 27134
rect 26012 26450 26068 26460
rect 24556 26292 24612 26302
rect 24108 26290 24276 26292
rect 24108 26238 24110 26290
rect 24162 26238 24276 26290
rect 24108 26236 24276 26238
rect 24332 26290 24612 26292
rect 24332 26238 24558 26290
rect 24610 26238 24612 26290
rect 24332 26236 24612 26238
rect 24108 26226 24164 26236
rect 23996 26126 23998 26178
rect 24050 26126 24052 26178
rect 23996 26114 24052 26126
rect 24220 25284 24276 26236
rect 24556 26226 24612 26236
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 40012 25618 40068 25630
rect 40012 25566 40014 25618
rect 40066 25566 40068 25618
rect 37660 25506 37716 25518
rect 37660 25454 37662 25506
rect 37714 25454 37716 25506
rect 25564 25396 25620 25406
rect 25564 25302 25620 25340
rect 26684 25394 26740 25406
rect 26684 25342 26686 25394
rect 26738 25342 26740 25394
rect 23884 24722 23940 24734
rect 23884 24670 23886 24722
rect 23938 24670 23940 24722
rect 23660 23380 23716 23390
rect 23660 23286 23716 23324
rect 22316 23102 22318 23154
rect 22370 23102 22372 23154
rect 22316 22932 22372 23102
rect 22316 22866 22372 22876
rect 22764 23154 22932 23156
rect 22764 23102 22878 23154
rect 22930 23102 22932 23154
rect 22764 23100 22932 23102
rect 22764 22708 22820 23100
rect 22876 23090 22932 23100
rect 23100 23154 23380 23156
rect 23100 23102 23326 23154
rect 23378 23102 23380 23154
rect 23100 23100 23380 23102
rect 22988 23044 23044 23054
rect 22988 22950 23044 22988
rect 21756 22594 21924 22596
rect 21756 22542 21870 22594
rect 21922 22542 21924 22594
rect 21756 22540 21924 22542
rect 21420 22372 21476 22382
rect 21420 22278 21476 22316
rect 21644 22370 21700 22382
rect 21644 22318 21646 22370
rect 21698 22318 21700 22370
rect 20524 21810 20692 21812
rect 20524 21758 20526 21810
rect 20578 21758 20692 21810
rect 20524 21756 20692 21758
rect 20524 21746 20580 21756
rect 20188 20972 20356 21028
rect 20412 21588 20468 21598
rect 20188 20580 20244 20972
rect 20300 20804 20356 20814
rect 20412 20804 20468 21532
rect 20860 21588 20916 21598
rect 20860 21586 21252 21588
rect 20860 21534 20862 21586
rect 20914 21534 21252 21586
rect 20860 21532 21252 21534
rect 20860 21522 20916 21532
rect 20524 20804 20580 20814
rect 20412 20802 20580 20804
rect 20412 20750 20526 20802
rect 20578 20750 20580 20802
rect 20412 20748 20580 20750
rect 20300 20710 20356 20748
rect 20524 20738 20580 20748
rect 20636 20580 20692 20590
rect 20188 20578 20692 20580
rect 20188 20526 20638 20578
rect 20690 20526 20692 20578
rect 20188 20524 20692 20526
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19852 20130 19908 20142
rect 19852 20078 19854 20130
rect 19906 20078 19908 20130
rect 19852 19796 19908 20078
rect 20188 20132 20244 20524
rect 20636 20514 20692 20524
rect 20860 20580 20916 20590
rect 20860 20486 20916 20524
rect 20300 20132 20356 20142
rect 20188 20076 20300 20132
rect 20300 20038 20356 20076
rect 19852 19730 19908 19740
rect 19964 20020 20020 20030
rect 19964 19234 20020 19964
rect 20636 20020 20692 20030
rect 20692 19964 20804 20020
rect 20636 19926 20692 19964
rect 19964 19182 19966 19234
rect 20018 19182 20020 19234
rect 19964 19170 20020 19182
rect 20300 19234 20356 19246
rect 20300 19182 20302 19234
rect 20354 19182 20356 19234
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19964 18228 20020 18238
rect 19964 17554 20020 18172
rect 19964 17502 19966 17554
rect 20018 17502 20020 17554
rect 19964 17490 20020 17502
rect 20300 17666 20356 19182
rect 20748 18562 20804 19964
rect 20972 19908 21028 19918
rect 20972 19814 21028 19852
rect 21196 19348 21252 21532
rect 21308 20804 21364 20814
rect 21308 20710 21364 20748
rect 21644 20244 21700 22318
rect 21644 20178 21700 20188
rect 21532 20132 21588 20142
rect 21532 20038 21588 20076
rect 21308 19348 21364 19358
rect 21252 19346 21364 19348
rect 21252 19294 21310 19346
rect 21362 19294 21364 19346
rect 21252 19292 21364 19294
rect 21196 19254 21252 19292
rect 21308 19282 21364 19292
rect 20748 18510 20750 18562
rect 20802 18510 20804 18562
rect 20748 18498 20804 18510
rect 21420 19236 21476 19246
rect 20972 18228 21028 18238
rect 20972 18134 21028 18172
rect 21308 18226 21364 18238
rect 21308 18174 21310 18226
rect 21362 18174 21364 18226
rect 20300 17614 20302 17666
rect 20354 17614 20356 17666
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 17052 20020 17108
rect 18956 15876 19012 17052
rect 19180 16772 19236 16782
rect 19180 16098 19236 16716
rect 19964 16322 20020 17052
rect 20300 16772 20356 17614
rect 21308 17668 21364 18174
rect 21308 17602 21364 17612
rect 21308 17444 21364 17454
rect 21308 17350 21364 17388
rect 20300 16706 20356 16716
rect 20860 16994 20916 17006
rect 20860 16942 20862 16994
rect 20914 16942 20916 16994
rect 19964 16270 19966 16322
rect 20018 16270 20020 16322
rect 19964 16258 20020 16270
rect 19180 16046 19182 16098
rect 19234 16046 19236 16098
rect 19180 16034 19236 16046
rect 20300 16210 20356 16222
rect 20300 16158 20302 16210
rect 20354 16158 20356 16210
rect 19068 15876 19124 15886
rect 18956 15820 19068 15876
rect 19068 15782 19124 15820
rect 20188 15876 20244 15886
rect 20188 15782 20244 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20076 15428 20132 15438
rect 20300 15428 20356 16158
rect 20076 15426 20356 15428
rect 20076 15374 20078 15426
rect 20130 15374 20356 15426
rect 20076 15372 20356 15374
rect 20860 16212 20916 16942
rect 20076 15362 20132 15372
rect 19292 15314 19348 15326
rect 19292 15262 19294 15314
rect 19346 15262 19348 15314
rect 19292 15204 19348 15262
rect 19292 15138 19348 15148
rect 20860 15204 20916 16156
rect 21308 16772 21364 16782
rect 21308 16100 21364 16716
rect 21308 16006 21364 16044
rect 21420 16322 21476 19180
rect 21756 17668 21812 22540
rect 21868 22530 21924 22540
rect 21980 22652 22820 22708
rect 22876 22932 22932 22942
rect 21980 22594 22036 22652
rect 21980 22542 21982 22594
rect 22034 22542 22036 22594
rect 21980 22530 22036 22542
rect 22876 21812 22932 22876
rect 22988 22260 23044 22270
rect 23100 22260 23156 23100
rect 23324 23090 23380 23100
rect 23772 23044 23828 23054
rect 23772 22950 23828 22988
rect 22988 22258 23156 22260
rect 22988 22206 22990 22258
rect 23042 22206 23156 22258
rect 22988 22204 23156 22206
rect 22988 22194 23044 22204
rect 22876 21746 22932 21756
rect 23324 22146 23380 22158
rect 23324 22094 23326 22146
rect 23378 22094 23380 22146
rect 22652 21588 22708 21598
rect 22652 20242 22708 21532
rect 23324 21588 23380 22094
rect 23324 21522 23380 21532
rect 23772 21588 23828 21598
rect 23772 21494 23828 21532
rect 23884 20916 23940 24670
rect 24108 21700 24164 21710
rect 24220 21700 24276 25228
rect 25228 25284 25284 25294
rect 25228 25190 25284 25228
rect 26460 25284 26516 25294
rect 25340 24722 25396 24734
rect 25340 24670 25342 24722
rect 25394 24670 25396 24722
rect 25340 24612 25396 24670
rect 24892 24052 24948 24062
rect 24892 23492 24948 23996
rect 24892 23426 24948 23436
rect 25340 23716 25396 24556
rect 26124 24612 26180 24622
rect 26124 24610 26404 24612
rect 26124 24558 26126 24610
rect 26178 24558 26404 24610
rect 26124 24556 26404 24558
rect 26124 24546 26180 24556
rect 26124 24276 26180 24286
rect 25676 23938 25732 23950
rect 25676 23886 25678 23938
rect 25730 23886 25732 23938
rect 25676 23716 25732 23886
rect 25340 23714 25732 23716
rect 25340 23662 25342 23714
rect 25394 23662 25732 23714
rect 25340 23660 25732 23662
rect 25228 23156 25284 23166
rect 25228 21812 25284 23100
rect 25340 23044 25396 23660
rect 26124 23378 26180 24220
rect 26124 23326 26126 23378
rect 26178 23326 26180 23378
rect 26124 23314 26180 23326
rect 26348 23378 26404 24556
rect 26460 24050 26516 25228
rect 26684 24388 26740 25342
rect 26908 25394 26964 25406
rect 26908 25342 26910 25394
rect 26962 25342 26964 25394
rect 26908 24948 26964 25342
rect 27244 25396 27300 25406
rect 27580 25396 27636 25406
rect 27300 25394 27636 25396
rect 27300 25342 27582 25394
rect 27634 25342 27636 25394
rect 27300 25340 27636 25342
rect 27244 25302 27300 25340
rect 27580 25330 27636 25340
rect 27020 25284 27076 25294
rect 27020 25190 27076 25228
rect 27692 25282 27748 25294
rect 27692 25230 27694 25282
rect 27746 25230 27748 25282
rect 26908 24882 26964 24892
rect 27692 24612 27748 25230
rect 27692 24546 27748 24556
rect 27916 25282 27972 25294
rect 27916 25230 27918 25282
rect 27970 25230 27972 25282
rect 26684 24322 26740 24332
rect 27916 24276 27972 25230
rect 28588 24948 28644 24958
rect 28588 24854 28644 24892
rect 37660 24948 37716 25454
rect 37660 24882 37716 24892
rect 40012 24948 40068 25566
rect 40012 24882 40068 24892
rect 28700 24836 28756 24846
rect 28252 24612 28308 24622
rect 28252 24518 28308 24556
rect 27916 24210 27972 24220
rect 26460 23998 26462 24050
rect 26514 23998 26516 24050
rect 26460 23986 26516 23998
rect 28588 24052 28644 24062
rect 28700 24052 28756 24780
rect 37660 24724 37716 24734
rect 37660 24630 37716 24668
rect 40012 24498 40068 24510
rect 40012 24446 40014 24498
rect 40066 24446 40068 24498
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 40012 24276 40068 24446
rect 40012 24210 40068 24220
rect 28588 24050 28756 24052
rect 28588 23998 28590 24050
rect 28642 23998 28756 24050
rect 28588 23996 28756 23998
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 28588 23986 28644 23996
rect 37660 23940 37716 23950
rect 37660 23846 37716 23884
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 26348 23326 26350 23378
rect 26402 23326 26404 23378
rect 26348 23314 26404 23326
rect 26012 23156 26068 23166
rect 26012 23062 26068 23100
rect 25340 23042 25508 23044
rect 25340 22990 25342 23042
rect 25394 22990 25508 23042
rect 25340 22988 25508 22990
rect 25340 22978 25396 22988
rect 25340 21812 25396 21822
rect 25228 21810 25396 21812
rect 25228 21758 25342 21810
rect 25394 21758 25396 21810
rect 25228 21756 25396 21758
rect 25340 21746 25396 21756
rect 24108 21698 24276 21700
rect 24108 21646 24110 21698
rect 24162 21646 24276 21698
rect 24108 21644 24276 21646
rect 24108 21634 24164 21644
rect 23772 20914 23940 20916
rect 23772 20862 23886 20914
rect 23938 20862 23940 20914
rect 23772 20860 23940 20862
rect 22652 20190 22654 20242
rect 22706 20190 22708 20242
rect 22652 20178 22708 20190
rect 23100 20244 23156 20254
rect 21868 20130 21924 20142
rect 21868 20078 21870 20130
rect 21922 20078 21924 20130
rect 21868 20020 21924 20078
rect 22764 20132 22820 20142
rect 22764 20038 22820 20076
rect 23100 20132 23156 20188
rect 23212 20132 23268 20142
rect 23100 20130 23268 20132
rect 23100 20078 23214 20130
rect 23266 20078 23268 20130
rect 23100 20076 23268 20078
rect 22092 20020 22148 20030
rect 21868 19234 21924 19964
rect 21980 20018 22148 20020
rect 21980 19966 22094 20018
rect 22146 19966 22148 20018
rect 21980 19964 22148 19966
rect 21980 19348 22036 19964
rect 22092 19954 22148 19964
rect 22540 19796 22596 19806
rect 21980 19282 22036 19292
rect 22092 19794 22596 19796
rect 22092 19742 22542 19794
rect 22594 19742 22596 19794
rect 22092 19740 22596 19742
rect 21868 19182 21870 19234
rect 21922 19182 21924 19234
rect 21868 19170 21924 19182
rect 22092 19236 22148 19740
rect 22540 19730 22596 19740
rect 22092 19142 22148 19180
rect 21644 17556 21700 17566
rect 21756 17556 21812 17612
rect 21644 17554 21812 17556
rect 21644 17502 21646 17554
rect 21698 17502 21812 17554
rect 21644 17500 21812 17502
rect 22428 17668 22484 17678
rect 21644 17490 21700 17500
rect 21420 16270 21422 16322
rect 21474 16270 21476 16322
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20188 13860 20244 13870
rect 20188 13766 20244 13804
rect 20748 13748 20804 13758
rect 20300 13746 20804 13748
rect 20300 13694 20750 13746
rect 20802 13694 20804 13746
rect 20300 13692 20804 13694
rect 20076 13524 20132 13534
rect 20076 13430 20132 13468
rect 20300 13074 20356 13692
rect 20748 13682 20804 13692
rect 20412 13524 20468 13534
rect 20748 13524 20804 13534
rect 20412 13522 20804 13524
rect 20412 13470 20414 13522
rect 20466 13470 20750 13522
rect 20802 13470 20804 13522
rect 20412 13468 20804 13470
rect 20412 13458 20468 13468
rect 20748 13458 20804 13468
rect 20748 13076 20804 13086
rect 20860 13076 20916 15148
rect 21420 14532 21476 16270
rect 22092 16212 22148 16222
rect 22092 16118 22148 16156
rect 22204 16100 22260 16110
rect 21644 15876 21700 15886
rect 21644 14754 21700 15820
rect 22204 15202 22260 16044
rect 22428 16098 22484 17612
rect 22876 17668 22932 17678
rect 22876 17574 22932 17612
rect 22540 17444 22596 17454
rect 22540 16322 22596 17388
rect 22540 16270 22542 16322
rect 22594 16270 22596 16322
rect 22540 16258 22596 16270
rect 22428 16046 22430 16098
rect 22482 16046 22484 16098
rect 22428 16034 22484 16046
rect 22652 16212 22708 16222
rect 22652 16100 22708 16156
rect 22988 16100 23044 16110
rect 22652 16098 23044 16100
rect 22652 16046 22990 16098
rect 23042 16046 23044 16098
rect 22652 16044 23044 16046
rect 22540 15988 22596 15998
rect 22540 15894 22596 15932
rect 22652 15540 22708 16044
rect 22988 16034 23044 16044
rect 22652 15446 22708 15484
rect 22204 15150 22206 15202
rect 22258 15150 22260 15202
rect 22204 15138 22260 15150
rect 23100 15148 23156 20076
rect 23212 20066 23268 20076
rect 23436 20132 23492 20142
rect 23436 20018 23492 20076
rect 23436 19966 23438 20018
rect 23490 19966 23492 20018
rect 23436 19460 23492 19966
rect 23436 19394 23492 19404
rect 23772 19124 23828 20860
rect 23884 20850 23940 20860
rect 23884 20018 23940 20030
rect 23884 19966 23886 20018
rect 23938 19966 23940 20018
rect 23884 19796 23940 19966
rect 24108 20018 24164 20030
rect 24108 19966 24110 20018
rect 24162 19966 24164 20018
rect 23996 19908 24052 19918
rect 23996 19814 24052 19852
rect 23884 19730 23940 19740
rect 23884 19460 23940 19470
rect 23884 19366 23940 19404
rect 23996 19348 24052 19358
rect 23996 19254 24052 19292
rect 23772 19058 23828 19068
rect 24108 18004 24164 19966
rect 23548 17948 24164 18004
rect 23548 17666 23604 17948
rect 23548 17614 23550 17666
rect 23602 17614 23604 17666
rect 23324 17554 23380 17566
rect 23324 17502 23326 17554
rect 23378 17502 23380 17554
rect 23212 17442 23268 17454
rect 23212 17390 23214 17442
rect 23266 17390 23268 17442
rect 23212 17108 23268 17390
rect 23212 17042 23268 17052
rect 23324 15988 23380 17502
rect 23324 15922 23380 15932
rect 23436 17444 23492 17454
rect 23100 15092 23380 15148
rect 21644 14702 21646 14754
rect 21698 14702 21700 14754
rect 21644 14690 21700 14702
rect 22764 14644 22820 14654
rect 21084 14476 21420 14532
rect 21084 13858 21140 14476
rect 21420 14466 21476 14476
rect 22428 14532 22484 14542
rect 22428 14438 22484 14476
rect 21868 14420 21924 14430
rect 21868 14326 21924 14364
rect 22764 14420 22820 14588
rect 22764 14418 23044 14420
rect 22764 14366 22766 14418
rect 22818 14366 23044 14418
rect 22764 14364 23044 14366
rect 22764 14354 22820 14364
rect 21308 14308 21364 14318
rect 21308 14306 21588 14308
rect 21308 14254 21310 14306
rect 21362 14254 21588 14306
rect 21308 14252 21588 14254
rect 21308 14242 21364 14252
rect 21084 13806 21086 13858
rect 21138 13806 21140 13858
rect 21084 13794 21140 13806
rect 21532 13860 21588 14252
rect 21420 13076 21476 13086
rect 20300 13022 20302 13074
rect 20354 13022 20356 13074
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 18844 12238 18846 12290
rect 18898 12238 18900 12290
rect 18844 12226 18900 12238
rect 18620 12126 18622 12178
rect 18674 12126 18676 12178
rect 18620 12114 18676 12126
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 20300 8428 20356 13022
rect 20524 13074 20860 13076
rect 20524 13022 20750 13074
rect 20802 13022 20860 13074
rect 20524 13020 20860 13022
rect 20524 12178 20580 13020
rect 20748 13010 20804 13020
rect 20860 12982 20916 13020
rect 21196 13074 21476 13076
rect 21196 13022 21422 13074
rect 21474 13022 21476 13074
rect 21196 13020 21476 13022
rect 21196 12290 21252 13020
rect 21420 13010 21476 13020
rect 21532 12850 21588 13804
rect 22764 13860 22820 13870
rect 22764 13858 22932 13860
rect 22764 13806 22766 13858
rect 22818 13806 22932 13858
rect 22764 13804 22932 13806
rect 22764 13794 22820 13804
rect 21756 13524 21812 13534
rect 21756 13186 21812 13468
rect 22652 13524 22708 13534
rect 22652 13430 22708 13468
rect 21756 13134 21758 13186
rect 21810 13134 21812 13186
rect 21756 13122 21812 13134
rect 22764 13076 22820 13086
rect 22764 12982 22820 13020
rect 21532 12798 21534 12850
rect 21586 12798 21588 12850
rect 21532 12786 21588 12798
rect 21196 12238 21198 12290
rect 21250 12238 21252 12290
rect 21196 12226 21252 12238
rect 20524 12126 20526 12178
rect 20578 12126 20580 12178
rect 20524 12114 20580 12126
rect 22876 12068 22932 13804
rect 22988 13858 23044 14364
rect 23324 14308 23380 15092
rect 23436 14530 23492 17388
rect 23548 14644 23604 17614
rect 23884 17556 23940 17566
rect 23884 17462 23940 17500
rect 23996 17442 24052 17454
rect 23996 17390 23998 17442
rect 24050 17390 24052 17442
rect 23772 16212 23828 16222
rect 23996 16212 24052 17390
rect 24108 17444 24164 17454
rect 24108 17350 24164 17388
rect 24220 17332 24276 21644
rect 25228 21586 25284 21598
rect 25228 21534 25230 21586
rect 25282 21534 25284 21586
rect 24332 20580 24388 20590
rect 24332 20130 24388 20524
rect 25228 20580 25284 21534
rect 25452 21476 25508 22988
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 25564 21700 25620 21710
rect 27020 21700 27076 21710
rect 25564 21698 26068 21700
rect 25564 21646 25566 21698
rect 25618 21646 26068 21698
rect 25564 21644 26068 21646
rect 25564 21634 25620 21644
rect 25900 21476 25956 21486
rect 25452 21474 25956 21476
rect 25452 21422 25902 21474
rect 25954 21422 25956 21474
rect 25452 21420 25956 21422
rect 25228 20514 25284 20524
rect 24332 20078 24334 20130
rect 24386 20078 24388 20130
rect 24332 19346 24388 20078
rect 25340 20020 25396 20030
rect 25900 20020 25956 21420
rect 26012 20130 26068 21644
rect 27020 21606 27076 21644
rect 27468 21698 27524 21710
rect 27468 21646 27470 21698
rect 27522 21646 27524 21698
rect 27468 21588 27524 21646
rect 27580 21700 27636 21710
rect 27580 21588 27636 21644
rect 27692 21588 27748 21598
rect 27580 21532 27692 21588
rect 27468 21522 27524 21532
rect 27692 21522 27748 21532
rect 29372 21588 29428 21598
rect 28588 21476 28644 21486
rect 26236 21364 26292 21374
rect 26012 20078 26014 20130
rect 26066 20078 26068 20130
rect 26012 20066 26068 20078
rect 26124 21308 26236 21364
rect 25340 20018 25956 20020
rect 25340 19966 25342 20018
rect 25394 19966 25956 20018
rect 25340 19964 25956 19966
rect 25340 19954 25396 19964
rect 24332 19294 24334 19346
rect 24386 19294 24388 19346
rect 24332 19282 24388 19294
rect 25228 19908 25284 19918
rect 26124 19908 26180 21308
rect 26236 21298 26292 21308
rect 27468 21364 27524 21374
rect 27468 21270 27524 21308
rect 24444 19236 24500 19246
rect 25004 19236 25060 19246
rect 24444 19234 25060 19236
rect 24444 19182 24446 19234
rect 24498 19182 25006 19234
rect 25058 19182 25060 19234
rect 24444 19180 25060 19182
rect 24444 19170 24500 19180
rect 25004 19170 25060 19180
rect 24220 17266 24276 17276
rect 24332 19124 24388 19134
rect 24332 16882 24388 19068
rect 24780 19010 24836 19022
rect 24780 18958 24782 19010
rect 24834 18958 24836 19010
rect 24668 18340 24724 18350
rect 24668 18246 24724 18284
rect 24444 17668 24500 17678
rect 24668 17668 24724 17678
rect 24444 17666 24724 17668
rect 24444 17614 24446 17666
rect 24498 17614 24670 17666
rect 24722 17614 24724 17666
rect 24444 17612 24724 17614
rect 24444 17602 24500 17612
rect 24668 17602 24724 17612
rect 24780 17108 24836 18958
rect 24892 19010 24948 19022
rect 24892 18958 24894 19010
rect 24946 18958 24948 19010
rect 24892 18452 24948 18958
rect 25228 18564 25284 19852
rect 25564 19852 26180 19908
rect 28140 19906 28196 19918
rect 28140 19854 28142 19906
rect 28194 19854 28196 19906
rect 25452 19236 25508 19246
rect 25452 19142 25508 19180
rect 25564 18674 25620 19852
rect 28140 19348 28196 19854
rect 28140 19282 28196 19292
rect 28588 19346 28644 21420
rect 28588 19294 28590 19346
rect 28642 19294 28644 19346
rect 28588 19282 28644 19294
rect 29372 19348 29428 21532
rect 37660 21588 37716 21598
rect 37660 21494 37716 21532
rect 40012 21362 40068 21374
rect 40012 21310 40014 21362
rect 40066 21310 40068 21362
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 40012 20916 40068 21310
rect 40012 20850 40068 20860
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 29820 19348 29876 19358
rect 29372 19346 29876 19348
rect 29372 19294 29822 19346
rect 29874 19294 29876 19346
rect 29372 19292 29876 19294
rect 25564 18622 25566 18674
rect 25618 18622 25620 18674
rect 25564 18610 25620 18622
rect 25676 19234 25732 19246
rect 25676 19182 25678 19234
rect 25730 19182 25732 19234
rect 25452 18564 25508 18574
rect 25228 18562 25508 18564
rect 25228 18510 25454 18562
rect 25506 18510 25508 18562
rect 25228 18508 25508 18510
rect 25452 18498 25508 18508
rect 24892 18386 24948 18396
rect 25676 18340 25732 19182
rect 29036 19236 29092 19246
rect 29036 19142 29092 19180
rect 29372 19234 29428 19292
rect 29820 19282 29876 19292
rect 40012 19346 40068 19358
rect 40012 19294 40014 19346
rect 40066 19294 40068 19346
rect 29372 19182 29374 19234
rect 29426 19182 29428 19234
rect 29372 19170 29428 19182
rect 37660 19236 37716 19246
rect 37660 19142 37716 19180
rect 26460 19124 26516 19134
rect 25788 19122 26516 19124
rect 25788 19070 26462 19122
rect 26514 19070 26516 19122
rect 25788 19068 26516 19070
rect 25788 18674 25844 19068
rect 26460 19058 26516 19068
rect 29260 19012 29316 19022
rect 25788 18622 25790 18674
rect 25842 18622 25844 18674
rect 25788 18610 25844 18622
rect 28924 18956 29260 19012
rect 25004 17554 25060 17566
rect 25004 17502 25006 17554
rect 25058 17502 25060 17554
rect 24780 17042 24836 17052
rect 24892 17442 24948 17454
rect 24892 17390 24894 17442
rect 24946 17390 24948 17442
rect 24332 16830 24334 16882
rect 24386 16830 24388 16882
rect 24332 16818 24388 16830
rect 24892 16884 24948 17390
rect 25004 17332 25060 17502
rect 25004 17266 25060 17276
rect 25676 17442 25732 18284
rect 26124 18450 26180 18462
rect 26124 18398 26126 18450
rect 26178 18398 26180 18450
rect 26124 18340 26180 18398
rect 26796 18452 26852 18462
rect 26796 18358 26852 18396
rect 26124 18274 26180 18284
rect 28924 18338 28980 18956
rect 29260 18918 29316 18956
rect 40012 18900 40068 19294
rect 40012 18834 40068 18844
rect 28924 18286 28926 18338
rect 28978 18286 28980 18338
rect 28924 18274 28980 18286
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 25676 17390 25678 17442
rect 25730 17390 25732 17442
rect 25676 17108 25732 17390
rect 28028 17668 28084 17678
rect 26460 17332 26516 17342
rect 24892 16818 24948 16828
rect 25452 17052 25732 17108
rect 25788 17108 25844 17118
rect 23772 16210 24052 16212
rect 23772 16158 23774 16210
rect 23826 16158 24052 16210
rect 23772 16156 24052 16158
rect 23772 16146 23828 16156
rect 24668 15540 24724 15550
rect 25452 15540 25508 17052
rect 25788 17014 25844 17052
rect 26460 16994 26516 17276
rect 26460 16942 26462 16994
rect 26514 16942 26516 16994
rect 26460 16930 26516 16942
rect 26572 16996 26628 17006
rect 26572 16902 26628 16940
rect 28028 16996 28084 17612
rect 37660 17668 37716 17678
rect 37660 17574 37716 17612
rect 25564 16884 25620 16894
rect 25564 16790 25620 16828
rect 26236 16884 26292 16894
rect 26236 16882 26404 16884
rect 26236 16830 26238 16882
rect 26290 16830 26404 16882
rect 26236 16828 26404 16830
rect 26236 16818 26292 16828
rect 25676 16772 25732 16782
rect 25676 16770 26180 16772
rect 25676 16718 25678 16770
rect 25730 16718 26180 16770
rect 25676 16716 26180 16718
rect 25676 16706 25732 16716
rect 25564 16660 25620 16670
rect 25564 16324 25620 16604
rect 26124 16436 26180 16716
rect 26348 16660 26404 16828
rect 26572 16660 26628 16670
rect 26348 16658 26628 16660
rect 26348 16606 26574 16658
rect 26626 16606 26628 16658
rect 26348 16604 26628 16606
rect 26572 16594 26628 16604
rect 26124 16380 26404 16436
rect 25564 16268 25956 16324
rect 25900 16212 25956 16268
rect 25900 16210 26292 16212
rect 25900 16158 25902 16210
rect 25954 16158 26292 16210
rect 25900 16156 26292 16158
rect 25564 15540 25620 15550
rect 25452 15484 25564 15540
rect 24668 15446 24724 15484
rect 25564 15314 25620 15484
rect 25564 15262 25566 15314
rect 25618 15262 25620 15314
rect 25564 15250 25620 15262
rect 25900 15148 25956 16156
rect 26236 16098 26292 16156
rect 26236 16046 26238 16098
rect 26290 16046 26292 16098
rect 26236 16034 26292 16046
rect 26348 15426 26404 16380
rect 28028 16100 28084 16940
rect 37660 16884 37716 16894
rect 37436 16882 37716 16884
rect 37436 16830 37662 16882
rect 37714 16830 37716 16882
rect 37436 16828 37716 16830
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 28028 16098 28532 16100
rect 28028 16046 28030 16098
rect 28082 16046 28532 16098
rect 28028 16044 28532 16046
rect 28028 16034 28084 16044
rect 26572 15988 26628 15998
rect 26572 15894 26628 15932
rect 28252 15876 28308 15886
rect 28252 15782 28308 15820
rect 26348 15374 26350 15426
rect 26402 15374 26404 15426
rect 26348 15362 26404 15374
rect 25788 15092 25956 15148
rect 28476 15202 28532 16044
rect 37436 15988 37492 16828
rect 37660 16818 37716 16828
rect 40012 16884 40068 17726
rect 40012 16818 40068 16828
rect 39900 16770 39956 16782
rect 39900 16718 39902 16770
rect 39954 16718 39956 16770
rect 39900 16212 39956 16718
rect 39900 16146 39956 16156
rect 40012 16210 40068 16222
rect 40012 16158 40014 16210
rect 40066 16158 40068 16210
rect 37660 16100 37716 16110
rect 37660 16006 37716 16044
rect 37436 15922 37492 15932
rect 40012 15540 40068 16158
rect 40012 15474 40068 15484
rect 28476 15150 28478 15202
rect 28530 15150 28532 15202
rect 28476 15138 28532 15150
rect 23996 14756 24052 14766
rect 23996 14754 24724 14756
rect 23996 14702 23998 14754
rect 24050 14702 24724 14754
rect 23996 14700 24724 14702
rect 23996 14690 24052 14700
rect 23604 14588 23940 14644
rect 23548 14550 23604 14588
rect 23436 14478 23438 14530
rect 23490 14478 23492 14530
rect 23436 14466 23492 14478
rect 23884 14532 23940 14588
rect 24668 14642 24724 14700
rect 24668 14590 24670 14642
rect 24722 14590 24724 14642
rect 24668 14578 24724 14590
rect 23996 14532 24052 14542
rect 23884 14530 24052 14532
rect 23884 14478 23998 14530
rect 24050 14478 24052 14530
rect 23884 14476 24052 14478
rect 23996 14466 24052 14476
rect 23660 14420 23716 14430
rect 23660 14308 23716 14364
rect 24556 14420 24612 14430
rect 24556 14326 24612 14364
rect 23324 14252 23716 14308
rect 23884 14306 23940 14318
rect 23884 14254 23886 14306
rect 23938 14254 23940 14306
rect 22988 13806 22990 13858
rect 23042 13806 23044 13858
rect 22988 13794 23044 13806
rect 23100 13076 23156 13086
rect 23100 12962 23156 13020
rect 23100 12910 23102 12962
rect 23154 12910 23156 12962
rect 23100 12898 23156 12910
rect 23772 13076 23828 13086
rect 23772 12402 23828 13020
rect 23884 13074 23940 14254
rect 23884 13022 23886 13074
rect 23938 13022 23940 13074
rect 23884 13010 23940 13022
rect 24780 14306 24836 14318
rect 24780 14254 24782 14306
rect 24834 14254 24836 14306
rect 24780 13076 24836 14254
rect 24780 13010 24836 13020
rect 25228 13076 25284 13086
rect 23772 12350 23774 12402
rect 23826 12350 23828 12402
rect 23772 12338 23828 12350
rect 23324 12068 23380 12078
rect 22876 12066 23380 12068
rect 22876 12014 23326 12066
rect 23378 12014 23380 12066
rect 22876 12012 23380 12014
rect 23324 11508 23380 12012
rect 23324 11442 23380 11452
rect 24556 11508 24612 11518
rect 20300 8372 20804 8428
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 20748 3554 20804 8372
rect 20748 3502 20750 3554
rect 20802 3502 20804 3554
rect 20748 3490 20804 3502
rect 22876 3668 22932 3678
rect 20188 3444 20244 3454
rect 19068 3332 19124 3342
rect 18844 3330 19124 3332
rect 18844 3278 19070 3330
rect 19122 3278 19124 3330
rect 18844 3276 19124 3278
rect 18844 800 18900 3276
rect 19068 3266 19124 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 800 20244 3388
rect 21756 3444 21812 3454
rect 21756 3330 21812 3388
rect 21756 3278 21758 3330
rect 21810 3278 21812 3330
rect 21756 3266 21812 3278
rect 22876 800 22932 3612
rect 24556 3554 24612 11452
rect 25228 4338 25284 13020
rect 25228 4286 25230 4338
rect 25282 4286 25284 4338
rect 25228 4274 25284 4286
rect 25676 5236 25732 5246
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 24892 4116 24948 4126
rect 24892 800 24948 4060
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 25676 2436 25732 5180
rect 25788 5122 25844 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 26012 13076 26068 13086
rect 26012 12982 26068 13020
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 26796 5236 26852 5246
rect 26796 5142 26852 5180
rect 25788 5070 25790 5122
rect 25842 5070 25844 5122
rect 25788 5058 25844 5070
rect 26236 4116 26292 4126
rect 26236 4022 26292 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 25564 2380 25732 2436
rect 25564 800 25620 2380
rect 18816 0 18928 800
rect 20160 0 20272 800
rect 22848 0 22960 800
rect 24864 0 24976 800
rect 25536 0 25648 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 16828 38220 16884 38276
rect 18060 38274 18116 38276
rect 18060 38222 18062 38274
rect 18062 38222 18114 38274
rect 18114 38222 18116 38274
rect 18060 38220 18116 38222
rect 1708 36988 1764 37044
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 24892 38220 24948 38276
rect 20860 37436 20916 37492
rect 20188 36652 20244 36708
rect 20300 36428 20356 36484
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 21308 36482 21364 36484
rect 21308 36430 21310 36482
rect 21310 36430 21362 36482
rect 21362 36430 21364 36482
rect 21308 36428 21364 36430
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4172 27580 4228 27636
rect 1932 24892 1988 24948
rect 1932 23548 1988 23604
rect 1932 22930 1988 22932
rect 1932 22878 1934 22930
rect 1934 22878 1986 22930
rect 1986 22878 1988 22930
rect 1932 22876 1988 22878
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 14140 27132 14196 27188
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 17388 28476 17444 28532
rect 17948 28476 18004 28532
rect 18508 28476 18564 28532
rect 19292 27746 19348 27748
rect 19292 27694 19294 27746
rect 19294 27694 19346 27746
rect 19346 27694 19348 27746
rect 19292 27692 19348 27694
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 17388 27186 17444 27188
rect 17388 27134 17390 27186
rect 17390 27134 17442 27186
rect 17442 27134 17444 27186
rect 17388 27132 17444 27134
rect 14812 26460 14868 26516
rect 15708 26514 15764 26516
rect 15708 26462 15710 26514
rect 15710 26462 15762 26514
rect 15762 26462 15764 26514
rect 15708 26460 15764 26462
rect 15820 26178 15876 26180
rect 15820 26126 15822 26178
rect 15822 26126 15874 26178
rect 15874 26126 15876 26178
rect 15820 26124 15876 26126
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4284 25506 4340 25508
rect 4284 25454 4286 25506
rect 4286 25454 4338 25506
rect 4338 25454 4340 25506
rect 4284 25452 4340 25454
rect 13916 25452 13972 25508
rect 19740 26962 19796 26964
rect 19740 26910 19742 26962
rect 19742 26910 19794 26962
rect 19794 26910 19796 26962
rect 19740 26908 19796 26910
rect 17836 26796 17892 26852
rect 20076 26796 20132 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 17612 26290 17668 26292
rect 17612 26238 17614 26290
rect 17614 26238 17666 26290
rect 17666 26238 17668 26290
rect 17612 26236 17668 26238
rect 17724 26178 17780 26180
rect 17724 26126 17726 26178
rect 17726 26126 17778 26178
rect 17778 26126 17780 26178
rect 17724 26124 17780 26126
rect 15148 24892 15204 24948
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 16828 25228 16884 25284
rect 15932 24668 15988 24724
rect 16492 24668 16548 24724
rect 4284 23938 4340 23940
rect 4284 23886 4286 23938
rect 4286 23886 4338 23938
rect 4338 23886 4340 23938
rect 4284 23884 4340 23886
rect 11452 23884 11508 23940
rect 4284 23154 4340 23156
rect 4284 23102 4286 23154
rect 4286 23102 4338 23154
rect 4338 23102 4340 23154
rect 4284 23100 4340 23102
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 12012 23436 12068 23492
rect 14140 23324 14196 23380
rect 12012 23100 12068 23156
rect 16156 23996 16212 24052
rect 15596 23436 15652 23492
rect 15484 23378 15540 23380
rect 15484 23326 15486 23378
rect 15486 23326 15538 23378
rect 15538 23326 15540 23378
rect 15484 23324 15540 23326
rect 13804 22876 13860 22932
rect 11452 22316 11508 22372
rect 13580 22146 13636 22148
rect 13580 22094 13582 22146
rect 13582 22094 13634 22146
rect 13634 22094 13636 22146
rect 13580 22092 13636 22094
rect 15596 23266 15652 23268
rect 15596 23214 15598 23266
rect 15598 23214 15650 23266
rect 15650 23214 15652 23266
rect 15596 23212 15652 23214
rect 15036 22876 15092 22932
rect 15260 22764 15316 22820
rect 15036 22370 15092 22372
rect 15036 22318 15038 22370
rect 15038 22318 15090 22370
rect 15090 22318 15092 22370
rect 15036 22316 15092 22318
rect 16156 23154 16212 23156
rect 16156 23102 16158 23154
rect 16158 23102 16210 23154
rect 16210 23102 16212 23154
rect 16156 23100 16212 23102
rect 15820 23042 15876 23044
rect 15820 22990 15822 23042
rect 15822 22990 15874 23042
rect 15874 22990 15876 23042
rect 15820 22988 15876 22990
rect 16156 22764 16212 22820
rect 15372 22146 15428 22148
rect 15372 22094 15374 22146
rect 15374 22094 15426 22146
rect 15426 22094 15428 22146
rect 15372 22092 15428 22094
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4172 20748 4228 20804
rect 4284 20412 4340 20468
rect 10892 20636 10948 20692
rect 1932 20188 1988 20244
rect 14476 20690 14532 20692
rect 14476 20638 14478 20690
rect 14478 20638 14530 20690
rect 14530 20638 14532 20690
rect 14476 20636 14532 20638
rect 14588 20076 14644 20132
rect 12236 19740 12292 19796
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 14476 19906 14532 19908
rect 14476 19854 14478 19906
rect 14478 19854 14530 19906
rect 14530 19854 14532 19906
rect 14476 19852 14532 19854
rect 14140 19794 14196 19796
rect 14140 19742 14142 19794
rect 14142 19742 14194 19794
rect 14194 19742 14196 19794
rect 14140 19740 14196 19742
rect 4284 18450 4340 18452
rect 4284 18398 4286 18450
rect 4286 18398 4338 18450
rect 4338 18398 4340 18450
rect 4284 18396 4340 18398
rect 13580 18450 13636 18452
rect 13580 18398 13582 18450
rect 13582 18398 13634 18450
rect 13634 18398 13636 18450
rect 13580 18396 13636 18398
rect 10668 18338 10724 18340
rect 10668 18286 10670 18338
rect 10670 18286 10722 18338
rect 10722 18286 10724 18338
rect 10668 18284 10724 18286
rect 1932 18226 1988 18228
rect 1932 18174 1934 18226
rect 1934 18174 1986 18226
rect 1986 18174 1988 18226
rect 1932 18172 1988 18174
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 10668 17724 10724 17780
rect 12236 18172 12292 18228
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 14476 18956 14532 19012
rect 13804 18226 13860 18228
rect 13804 18174 13806 18226
rect 13806 18174 13858 18226
rect 13858 18174 13860 18226
rect 13804 18172 13860 18174
rect 13804 17890 13860 17892
rect 13804 17838 13806 17890
rect 13806 17838 13858 17890
rect 13858 17838 13860 17890
rect 13804 17836 13860 17838
rect 16828 24050 16884 24052
rect 16828 23998 16830 24050
rect 16830 23998 16882 24050
rect 16882 23998 16884 24050
rect 16828 23996 16884 23998
rect 17612 24892 17668 24948
rect 17164 23324 17220 23380
rect 16828 23100 16884 23156
rect 16716 22370 16772 22372
rect 16716 22318 16718 22370
rect 16718 22318 16770 22370
rect 16770 22318 16772 22370
rect 16716 22316 16772 22318
rect 17276 23100 17332 23156
rect 17612 23212 17668 23268
rect 17388 22930 17444 22932
rect 17388 22878 17390 22930
rect 17390 22878 17442 22930
rect 17442 22878 17444 22930
rect 17388 22876 17444 22878
rect 15484 20130 15540 20132
rect 15484 20078 15486 20130
rect 15486 20078 15538 20130
rect 15538 20078 15540 20130
rect 15484 20076 15540 20078
rect 15372 20018 15428 20020
rect 15372 19966 15374 20018
rect 15374 19966 15426 20018
rect 15426 19966 15428 20018
rect 15372 19964 15428 19966
rect 15596 19906 15652 19908
rect 15596 19854 15598 19906
rect 15598 19854 15650 19906
rect 15650 19854 15652 19906
rect 15596 19852 15652 19854
rect 16268 19740 16324 19796
rect 14812 17836 14868 17892
rect 15148 18450 15204 18452
rect 15148 18398 15150 18450
rect 15150 18398 15202 18450
rect 15202 18398 15204 18450
rect 15148 18396 15204 18398
rect 13580 17778 13636 17780
rect 13580 17726 13582 17778
rect 13582 17726 13634 17778
rect 13634 17726 13636 17778
rect 13580 17724 13636 17726
rect 15708 18844 15764 18900
rect 16268 19068 16324 19124
rect 16492 19234 16548 19236
rect 16492 19182 16494 19234
rect 16494 19182 16546 19234
rect 16546 19182 16548 19234
rect 16492 19180 16548 19182
rect 16380 18956 16436 19012
rect 17164 19964 17220 20020
rect 17052 19852 17108 19908
rect 18732 26236 18788 26292
rect 21084 28588 21140 28644
rect 21308 27692 21364 27748
rect 22092 37490 22148 37492
rect 22092 37438 22094 37490
rect 22094 37438 22146 37490
rect 22146 37438 22148 37490
rect 22092 37436 22148 37438
rect 22316 36706 22372 36708
rect 22316 36654 22318 36706
rect 22318 36654 22370 36706
rect 22370 36654 22372 36706
rect 22316 36652 22372 36654
rect 21644 28642 21700 28644
rect 21644 28590 21646 28642
rect 21646 28590 21698 28642
rect 21698 28590 21700 28642
rect 21644 28588 21700 28590
rect 22092 28642 22148 28644
rect 22092 28590 22094 28642
rect 22094 28590 22146 28642
rect 22146 28590 22148 28642
rect 22092 28588 22148 28590
rect 26124 38274 26180 38276
rect 26124 38222 26126 38274
rect 26126 38222 26178 38274
rect 26178 38222 26180 38274
rect 26124 38220 26180 38222
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 25564 37436 25620 37492
rect 26796 37490 26852 37492
rect 26796 37438 26798 37490
rect 26798 37438 26850 37490
rect 26850 37438 26852 37490
rect 26796 37436 26852 37438
rect 20412 26962 20468 26964
rect 20412 26910 20414 26962
rect 20414 26910 20466 26962
rect 20466 26910 20468 26962
rect 20412 26908 20468 26910
rect 20748 26908 20804 26964
rect 21308 26908 21364 26964
rect 20300 26572 20356 26628
rect 20748 26572 20804 26628
rect 20524 26460 20580 26516
rect 18732 25340 18788 25396
rect 18060 24722 18116 24724
rect 18060 24670 18062 24722
rect 18062 24670 18114 24722
rect 18114 24670 18116 24722
rect 18060 24668 18116 24670
rect 18620 24722 18676 24724
rect 18620 24670 18622 24722
rect 18622 24670 18674 24722
rect 18674 24670 18676 24722
rect 18620 24668 18676 24670
rect 18508 24556 18564 24612
rect 18172 23212 18228 23268
rect 17836 22988 17892 23044
rect 18060 22988 18116 23044
rect 17612 21196 17668 21252
rect 17612 20524 17668 20580
rect 17500 19794 17556 19796
rect 17500 19742 17502 19794
rect 17502 19742 17554 19794
rect 17554 19742 17556 19794
rect 17500 19740 17556 19742
rect 17388 19068 17444 19124
rect 17276 18620 17332 18676
rect 16828 18508 16884 18564
rect 15036 16828 15092 16884
rect 14252 16210 14308 16212
rect 14252 16158 14254 16210
rect 14254 16158 14306 16210
rect 14306 16158 14308 16210
rect 14252 16156 14308 16158
rect 15820 16940 15876 16996
rect 15484 16156 15540 16212
rect 16044 17890 16100 17892
rect 16044 17838 16046 17890
rect 16046 17838 16098 17890
rect 16098 17838 16100 17890
rect 16044 17836 16100 17838
rect 16044 17666 16100 17668
rect 16044 17614 16046 17666
rect 16046 17614 16098 17666
rect 16098 17614 16100 17666
rect 16044 17612 16100 17614
rect 17052 17666 17108 17668
rect 17052 17614 17054 17666
rect 17054 17614 17106 17666
rect 17106 17614 17108 17666
rect 17052 17612 17108 17614
rect 16492 17164 16548 17220
rect 16604 17388 16660 17444
rect 16380 17052 16436 17108
rect 17500 17052 17556 17108
rect 17948 21196 18004 21252
rect 17836 19852 17892 19908
rect 17836 18844 17892 18900
rect 18060 19852 18116 19908
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20524 24668 20580 24724
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 18620 23100 18676 23156
rect 21868 26572 21924 26628
rect 22540 27074 22596 27076
rect 22540 27022 22542 27074
rect 22542 27022 22594 27074
rect 22594 27022 22596 27074
rect 22540 27020 22596 27022
rect 22652 26962 22708 26964
rect 22652 26910 22654 26962
rect 22654 26910 22706 26962
rect 22706 26910 22708 26962
rect 22652 26908 22708 26910
rect 22204 26460 22260 26516
rect 22428 26348 22484 26404
rect 23100 26402 23156 26404
rect 23100 26350 23102 26402
rect 23102 26350 23154 26402
rect 23154 26350 23156 26402
rect 23100 26348 23156 26350
rect 21420 24892 21476 24948
rect 21868 24556 21924 24612
rect 22092 24556 22148 24612
rect 24668 27020 24724 27076
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 23324 26908 23380 26964
rect 22652 24610 22708 24612
rect 22652 24558 22654 24610
rect 22654 24558 22706 24610
rect 22706 24558 22708 24610
rect 22652 24556 22708 24558
rect 22316 24332 22372 24388
rect 20524 23042 20580 23044
rect 20524 22990 20526 23042
rect 20526 22990 20578 23042
rect 20578 22990 20580 23042
rect 20524 22988 20580 22990
rect 19180 22316 19236 22372
rect 18620 20860 18676 20916
rect 20076 22370 20132 22372
rect 20076 22318 20078 22370
rect 20078 22318 20130 22370
rect 20130 22318 20132 22370
rect 20076 22316 20132 22318
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19292 21532 19348 21588
rect 19852 21586 19908 21588
rect 19852 21534 19854 21586
rect 19854 21534 19906 21586
rect 19906 21534 19908 21586
rect 19852 21532 19908 21534
rect 19516 20860 19572 20916
rect 18508 19740 18564 19796
rect 19068 20578 19124 20580
rect 19068 20526 19070 20578
rect 19070 20526 19122 20578
rect 19122 20526 19124 20578
rect 19068 20524 19124 20526
rect 18172 19292 18228 19348
rect 18732 19180 18788 19236
rect 18508 18562 18564 18564
rect 18508 18510 18510 18562
rect 18510 18510 18562 18562
rect 18562 18510 18564 18562
rect 18508 18508 18564 18510
rect 18060 17612 18116 17668
rect 18284 17666 18340 17668
rect 18284 17614 18286 17666
rect 18286 17614 18338 17666
rect 18338 17614 18340 17666
rect 18284 17612 18340 17614
rect 17948 17164 18004 17220
rect 15932 16156 15988 16212
rect 15820 15932 15876 15988
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 17724 16828 17780 16884
rect 17164 16210 17220 16212
rect 17164 16158 17166 16210
rect 17166 16158 17218 16210
rect 17218 16158 17220 16210
rect 17164 16156 17220 16158
rect 17388 15932 17444 15988
rect 16268 15314 16324 15316
rect 16268 15262 16270 15314
rect 16270 15262 16322 15314
rect 16322 15262 16324 15314
rect 16268 15260 16324 15262
rect 17500 15260 17556 15316
rect 18060 16156 18116 16212
rect 18060 15260 18116 15316
rect 18396 15932 18452 15988
rect 17724 14588 17780 14644
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 18508 15148 18564 15204
rect 18396 14642 18452 14644
rect 18396 14590 18398 14642
rect 18398 14590 18450 14642
rect 18450 14590 18452 14642
rect 18396 14588 18452 14590
rect 18620 13468 18676 13524
rect 19180 18172 19236 18228
rect 19404 19292 19460 19348
rect 19516 19068 19572 19124
rect 19516 18284 19572 18340
rect 19516 17666 19572 17668
rect 19516 17614 19518 17666
rect 19518 17614 19570 17666
rect 19570 17614 19572 17666
rect 19516 17612 19572 17614
rect 19180 17388 19236 17444
rect 19068 17164 19124 17220
rect 18956 17052 19012 17108
rect 21196 23266 21252 23268
rect 21196 23214 21198 23266
rect 21198 23214 21250 23266
rect 21250 23214 21252 23266
rect 21196 23212 21252 23214
rect 21980 23324 22036 23380
rect 20972 23154 21028 23156
rect 20972 23102 20974 23154
rect 20974 23102 21026 23154
rect 21026 23102 21028 23154
rect 20972 23100 21028 23102
rect 21308 23154 21364 23156
rect 21308 23102 21310 23154
rect 21310 23102 21362 23154
rect 21362 23102 21364 23154
rect 21308 23100 21364 23102
rect 22764 23324 22820 23380
rect 23100 23436 23156 23492
rect 22652 23266 22708 23268
rect 22652 23214 22654 23266
rect 22654 23214 22706 23266
rect 22706 23214 22708 23266
rect 22652 23212 22708 23214
rect 23436 26684 23492 26740
rect 23660 26514 23716 26516
rect 23660 26462 23662 26514
rect 23662 26462 23714 26514
rect 23714 26462 23716 26514
rect 23660 26460 23716 26462
rect 23884 26514 23940 26516
rect 23884 26462 23886 26514
rect 23886 26462 23938 26514
rect 23938 26462 23940 26514
rect 23884 26460 23940 26462
rect 26012 26460 26068 26516
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 25564 25394 25620 25396
rect 25564 25342 25566 25394
rect 25566 25342 25618 25394
rect 25618 25342 25620 25394
rect 25564 25340 25620 25342
rect 24220 25228 24276 25284
rect 23660 23378 23716 23380
rect 23660 23326 23662 23378
rect 23662 23326 23714 23378
rect 23714 23326 23716 23378
rect 23660 23324 23716 23326
rect 22316 22876 22372 22932
rect 22988 23042 23044 23044
rect 22988 22990 22990 23042
rect 22990 22990 23042 23042
rect 23042 22990 23044 23042
rect 22988 22988 23044 22990
rect 21420 22370 21476 22372
rect 21420 22318 21422 22370
rect 21422 22318 21474 22370
rect 21474 22318 21476 22370
rect 21420 22316 21476 22318
rect 20412 21532 20468 21588
rect 20300 20802 20356 20804
rect 20300 20750 20302 20802
rect 20302 20750 20354 20802
rect 20354 20750 20356 20802
rect 20300 20748 20356 20750
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20860 20578 20916 20580
rect 20860 20526 20862 20578
rect 20862 20526 20914 20578
rect 20914 20526 20916 20578
rect 20860 20524 20916 20526
rect 20300 20130 20356 20132
rect 20300 20078 20302 20130
rect 20302 20078 20354 20130
rect 20354 20078 20356 20130
rect 20300 20076 20356 20078
rect 19852 19740 19908 19796
rect 19964 19964 20020 20020
rect 20636 20018 20692 20020
rect 20636 19966 20638 20018
rect 20638 19966 20690 20018
rect 20690 19966 20692 20018
rect 20636 19964 20692 19966
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19964 18172 20020 18228
rect 20972 19906 21028 19908
rect 20972 19854 20974 19906
rect 20974 19854 21026 19906
rect 21026 19854 21028 19906
rect 20972 19852 21028 19854
rect 21308 20802 21364 20804
rect 21308 20750 21310 20802
rect 21310 20750 21362 20802
rect 21362 20750 21364 20802
rect 21308 20748 21364 20750
rect 21644 20188 21700 20244
rect 21532 20130 21588 20132
rect 21532 20078 21534 20130
rect 21534 20078 21586 20130
rect 21586 20078 21588 20130
rect 21532 20076 21588 20078
rect 21196 19292 21252 19348
rect 21420 19180 21476 19236
rect 20972 18226 21028 18228
rect 20972 18174 20974 18226
rect 20974 18174 21026 18226
rect 21026 18174 21028 18226
rect 20972 18172 21028 18174
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19180 16716 19236 16772
rect 21308 17612 21364 17668
rect 21308 17442 21364 17444
rect 21308 17390 21310 17442
rect 21310 17390 21362 17442
rect 21362 17390 21364 17442
rect 21308 17388 21364 17390
rect 20300 16716 20356 16772
rect 19068 15874 19124 15876
rect 19068 15822 19070 15874
rect 19070 15822 19122 15874
rect 19122 15822 19124 15874
rect 19068 15820 19124 15822
rect 20188 15874 20244 15876
rect 20188 15822 20190 15874
rect 20190 15822 20242 15874
rect 20242 15822 20244 15874
rect 20188 15820 20244 15822
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20860 16156 20916 16212
rect 19292 15148 19348 15204
rect 21308 16716 21364 16772
rect 21308 16098 21364 16100
rect 21308 16046 21310 16098
rect 21310 16046 21362 16098
rect 21362 16046 21364 16098
rect 21308 16044 21364 16046
rect 22876 22876 22932 22932
rect 23772 23042 23828 23044
rect 23772 22990 23774 23042
rect 23774 22990 23826 23042
rect 23826 22990 23828 23042
rect 23772 22988 23828 22990
rect 22876 21756 22932 21812
rect 22652 21532 22708 21588
rect 23324 21532 23380 21588
rect 23772 21586 23828 21588
rect 23772 21534 23774 21586
rect 23774 21534 23826 21586
rect 23826 21534 23828 21586
rect 23772 21532 23828 21534
rect 25228 25282 25284 25284
rect 25228 25230 25230 25282
rect 25230 25230 25282 25282
rect 25282 25230 25284 25282
rect 25228 25228 25284 25230
rect 26460 25228 26516 25284
rect 25340 24556 25396 24612
rect 24892 24050 24948 24052
rect 24892 23998 24894 24050
rect 24894 23998 24946 24050
rect 24946 23998 24948 24050
rect 24892 23996 24948 23998
rect 24892 23436 24948 23492
rect 26124 24220 26180 24276
rect 25228 23100 25284 23156
rect 27244 25394 27300 25396
rect 27244 25342 27246 25394
rect 27246 25342 27298 25394
rect 27298 25342 27300 25394
rect 27244 25340 27300 25342
rect 27020 25282 27076 25284
rect 27020 25230 27022 25282
rect 27022 25230 27074 25282
rect 27074 25230 27076 25282
rect 27020 25228 27076 25230
rect 26908 24892 26964 24948
rect 27692 24556 27748 24612
rect 26684 24332 26740 24388
rect 28588 24946 28644 24948
rect 28588 24894 28590 24946
rect 28590 24894 28642 24946
rect 28642 24894 28644 24946
rect 28588 24892 28644 24894
rect 37660 24892 37716 24948
rect 40012 24892 40068 24948
rect 28700 24834 28756 24836
rect 28700 24782 28702 24834
rect 28702 24782 28754 24834
rect 28754 24782 28756 24834
rect 28700 24780 28756 24782
rect 28252 24610 28308 24612
rect 28252 24558 28254 24610
rect 28254 24558 28306 24610
rect 28306 24558 28308 24610
rect 28252 24556 28308 24558
rect 27916 24220 27972 24276
rect 37660 24722 37716 24724
rect 37660 24670 37662 24722
rect 37662 24670 37714 24722
rect 37714 24670 37716 24722
rect 37660 24668 37716 24670
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 40012 24220 40068 24276
rect 37660 23938 37716 23940
rect 37660 23886 37662 23938
rect 37662 23886 37714 23938
rect 37714 23886 37716 23938
rect 37660 23884 37716 23886
rect 40012 23548 40068 23604
rect 26012 23154 26068 23156
rect 26012 23102 26014 23154
rect 26014 23102 26066 23154
rect 26066 23102 26068 23154
rect 26012 23100 26068 23102
rect 23100 20188 23156 20244
rect 22764 20130 22820 20132
rect 22764 20078 22766 20130
rect 22766 20078 22818 20130
rect 22818 20078 22820 20130
rect 22764 20076 22820 20078
rect 21868 19964 21924 20020
rect 21980 19292 22036 19348
rect 22092 19234 22148 19236
rect 22092 19182 22094 19234
rect 22094 19182 22146 19234
rect 22146 19182 22148 19234
rect 22092 19180 22148 19182
rect 21756 17612 21812 17668
rect 22428 17612 22484 17668
rect 20860 15148 20916 15204
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20188 13858 20244 13860
rect 20188 13806 20190 13858
rect 20190 13806 20242 13858
rect 20242 13806 20244 13858
rect 20188 13804 20244 13806
rect 20076 13522 20132 13524
rect 20076 13470 20078 13522
rect 20078 13470 20130 13522
rect 20130 13470 20132 13522
rect 20076 13468 20132 13470
rect 22092 16210 22148 16212
rect 22092 16158 22094 16210
rect 22094 16158 22146 16210
rect 22146 16158 22148 16210
rect 22092 16156 22148 16158
rect 22204 16044 22260 16100
rect 21644 15820 21700 15876
rect 22876 17666 22932 17668
rect 22876 17614 22878 17666
rect 22878 17614 22930 17666
rect 22930 17614 22932 17666
rect 22876 17612 22932 17614
rect 22540 17388 22596 17444
rect 22652 16156 22708 16212
rect 22540 15986 22596 15988
rect 22540 15934 22542 15986
rect 22542 15934 22594 15986
rect 22594 15934 22596 15986
rect 22540 15932 22596 15934
rect 22652 15538 22708 15540
rect 22652 15486 22654 15538
rect 22654 15486 22706 15538
rect 22706 15486 22708 15538
rect 22652 15484 22708 15486
rect 23436 20076 23492 20132
rect 23436 19404 23492 19460
rect 23996 19906 24052 19908
rect 23996 19854 23998 19906
rect 23998 19854 24050 19906
rect 24050 19854 24052 19906
rect 23996 19852 24052 19854
rect 23884 19740 23940 19796
rect 23884 19458 23940 19460
rect 23884 19406 23886 19458
rect 23886 19406 23938 19458
rect 23938 19406 23940 19458
rect 23884 19404 23940 19406
rect 23996 19346 24052 19348
rect 23996 19294 23998 19346
rect 23998 19294 24050 19346
rect 24050 19294 24052 19346
rect 23996 19292 24052 19294
rect 23772 19068 23828 19124
rect 23212 17052 23268 17108
rect 23324 15932 23380 15988
rect 23436 17388 23492 17444
rect 22764 14588 22820 14644
rect 21420 14476 21476 14532
rect 22428 14530 22484 14532
rect 22428 14478 22430 14530
rect 22430 14478 22482 14530
rect 22482 14478 22484 14530
rect 22428 14476 22484 14478
rect 21868 14418 21924 14420
rect 21868 14366 21870 14418
rect 21870 14366 21922 14418
rect 21922 14366 21924 14418
rect 21868 14364 21924 14366
rect 21532 13804 21588 13860
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 20860 13020 20916 13076
rect 21756 13468 21812 13524
rect 22652 13522 22708 13524
rect 22652 13470 22654 13522
rect 22654 13470 22706 13522
rect 22706 13470 22708 13522
rect 22652 13468 22708 13470
rect 22764 13074 22820 13076
rect 22764 13022 22766 13074
rect 22766 13022 22818 13074
rect 22818 13022 22820 13074
rect 22764 13020 22820 13022
rect 23884 17554 23940 17556
rect 23884 17502 23886 17554
rect 23886 17502 23938 17554
rect 23938 17502 23940 17554
rect 23884 17500 23940 17502
rect 24108 17442 24164 17444
rect 24108 17390 24110 17442
rect 24110 17390 24162 17442
rect 24162 17390 24164 17442
rect 24108 17388 24164 17390
rect 24332 20524 24388 20580
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 25228 20524 25284 20580
rect 27020 21698 27076 21700
rect 27020 21646 27022 21698
rect 27022 21646 27074 21698
rect 27074 21646 27076 21698
rect 27020 21644 27076 21646
rect 27468 21532 27524 21588
rect 27580 21698 27636 21700
rect 27580 21646 27582 21698
rect 27582 21646 27634 21698
rect 27634 21646 27636 21698
rect 27580 21644 27636 21646
rect 27692 21532 27748 21588
rect 29372 21532 29428 21588
rect 28588 21420 28644 21476
rect 26236 21308 26292 21364
rect 27468 21362 27524 21364
rect 27468 21310 27470 21362
rect 27470 21310 27522 21362
rect 27522 21310 27524 21362
rect 27468 21308 27524 21310
rect 25228 19852 25284 19908
rect 24220 17276 24276 17332
rect 24332 19068 24388 19124
rect 24668 18338 24724 18340
rect 24668 18286 24670 18338
rect 24670 18286 24722 18338
rect 24722 18286 24724 18338
rect 24668 18284 24724 18286
rect 25452 19234 25508 19236
rect 25452 19182 25454 19234
rect 25454 19182 25506 19234
rect 25506 19182 25508 19234
rect 25452 19180 25508 19182
rect 28140 19292 28196 19348
rect 37660 21586 37716 21588
rect 37660 21534 37662 21586
rect 37662 21534 37714 21586
rect 37714 21534 37716 21586
rect 37660 21532 37716 21534
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 40012 20860 40068 20916
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 24892 18396 24948 18452
rect 29036 19234 29092 19236
rect 29036 19182 29038 19234
rect 29038 19182 29090 19234
rect 29090 19182 29092 19234
rect 29036 19180 29092 19182
rect 37660 19234 37716 19236
rect 37660 19182 37662 19234
rect 37662 19182 37714 19234
rect 37714 19182 37716 19234
rect 37660 19180 37716 19182
rect 29260 19010 29316 19012
rect 29260 18958 29262 19010
rect 29262 18958 29314 19010
rect 29314 18958 29316 19010
rect 29260 18956 29316 18958
rect 25676 18284 25732 18340
rect 24780 17052 24836 17108
rect 25004 17276 25060 17332
rect 26796 18450 26852 18452
rect 26796 18398 26798 18450
rect 26798 18398 26850 18450
rect 26850 18398 26852 18450
rect 26796 18396 26852 18398
rect 26124 18284 26180 18340
rect 40012 18844 40068 18900
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 28028 17612 28084 17668
rect 26460 17276 26516 17332
rect 24892 16828 24948 16884
rect 25788 17106 25844 17108
rect 25788 17054 25790 17106
rect 25790 17054 25842 17106
rect 25842 17054 25844 17106
rect 25788 17052 25844 17054
rect 24668 15538 24724 15540
rect 24668 15486 24670 15538
rect 24670 15486 24722 15538
rect 24722 15486 24724 15538
rect 24668 15484 24724 15486
rect 26572 16994 26628 16996
rect 26572 16942 26574 16994
rect 26574 16942 26626 16994
rect 26626 16942 26628 16994
rect 26572 16940 26628 16942
rect 37660 17666 37716 17668
rect 37660 17614 37662 17666
rect 37662 17614 37714 17666
rect 37714 17614 37716 17666
rect 37660 17612 37716 17614
rect 28028 16940 28084 16996
rect 25564 16882 25620 16884
rect 25564 16830 25566 16882
rect 25566 16830 25618 16882
rect 25618 16830 25620 16882
rect 25564 16828 25620 16830
rect 25564 16604 25620 16660
rect 25564 15484 25620 15540
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 26572 15986 26628 15988
rect 26572 15934 26574 15986
rect 26574 15934 26626 15986
rect 26626 15934 26628 15986
rect 26572 15932 26628 15934
rect 28252 15874 28308 15876
rect 28252 15822 28254 15874
rect 28254 15822 28306 15874
rect 28306 15822 28308 15874
rect 28252 15820 28308 15822
rect 40012 16828 40068 16884
rect 39900 16156 39956 16212
rect 37660 16098 37716 16100
rect 37660 16046 37662 16098
rect 37662 16046 37714 16098
rect 37714 16046 37716 16098
rect 37660 16044 37716 16046
rect 37436 15932 37492 15988
rect 40012 15484 40068 15540
rect 23548 14588 23604 14644
rect 23660 14418 23716 14420
rect 23660 14366 23662 14418
rect 23662 14366 23714 14418
rect 23714 14366 23716 14418
rect 23660 14364 23716 14366
rect 24556 14418 24612 14420
rect 24556 14366 24558 14418
rect 24558 14366 24610 14418
rect 24610 14366 24612 14418
rect 24556 14364 24612 14366
rect 23100 13020 23156 13076
rect 23772 13020 23828 13076
rect 24780 13020 24836 13076
rect 25228 13020 25284 13076
rect 23324 11452 23380 11508
rect 24556 11452 24612 11508
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 22876 3612 22932 3668
rect 20188 3388 20244 3444
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 21756 3388 21812 3444
rect 25676 5180 25732 5236
rect 24892 4060 24948 4116
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 26012 13074 26068 13076
rect 26012 13022 26014 13074
rect 26014 13022 26066 13074
rect 26066 13022 26068 13074
rect 26012 13020 26068 13022
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 26796 5234 26852 5236
rect 26796 5182 26798 5234
rect 26798 5182 26850 5234
rect 26850 5182 26852 5234
rect 26796 5180 26852 5182
rect 26236 4114 26292 4116
rect 26236 4062 26238 4114
rect 26238 4062 26290 4114
rect 26290 4062 26292 4114
rect 26236 4060 26292 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 16818 38220 16828 38276
rect 16884 38220 18060 38276
rect 18116 38220 18126 38276
rect 24882 38220 24892 38276
rect 24948 38220 26124 38276
rect 26180 38220 26190 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 20850 37436 20860 37492
rect 20916 37436 22092 37492
rect 22148 37436 22158 37492
rect 25554 37436 25564 37492
rect 25620 37436 26796 37492
rect 26852 37436 26862 37492
rect 0 37044 800 37072
rect 0 36988 1708 37044
rect 1764 36988 1774 37044
rect 0 36960 800 36988
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 20178 36652 20188 36708
rect 20244 36652 22316 36708
rect 22372 36652 22382 36708
rect 20290 36428 20300 36484
rect 20356 36428 21308 36484
rect 21364 36428 21374 36484
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 20132 28588 21084 28644
rect 21140 28588 21644 28644
rect 21700 28588 22092 28644
rect 22148 28588 22158 28644
rect 20132 28532 20188 28588
rect 17378 28476 17388 28532
rect 17444 28476 17948 28532
rect 18004 28476 18508 28532
rect 18564 28476 20188 28532
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 19282 27692 19292 27748
rect 19348 27692 21308 27748
rect 21364 27692 21374 27748
rect 0 27636 800 27664
rect 0 27580 4172 27636
rect 4228 27580 4238 27636
rect 0 27552 800 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 14130 27132 14140 27188
rect 14196 27132 17388 27188
rect 17444 27132 17454 27188
rect 22530 27020 22540 27076
rect 22596 27020 24668 27076
rect 24724 27020 24734 27076
rect 19730 26908 19740 26964
rect 19796 26908 20412 26964
rect 20468 26908 20478 26964
rect 20738 26908 20748 26964
rect 20804 26908 21308 26964
rect 21364 26908 22652 26964
rect 22708 26908 23324 26964
rect 23380 26908 23390 26964
rect 17826 26796 17836 26852
rect 17892 26796 20076 26852
rect 20132 26796 20244 26852
rect 20188 26740 20244 26796
rect 20188 26684 23436 26740
rect 23492 26684 23502 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 20290 26572 20300 26628
rect 20356 26572 20748 26628
rect 20804 26572 21868 26628
rect 21924 26572 21934 26628
rect 14802 26460 14812 26516
rect 14868 26460 15708 26516
rect 15764 26460 15774 26516
rect 20514 26460 20524 26516
rect 20580 26460 22204 26516
rect 22260 26460 23660 26516
rect 23716 26460 23726 26516
rect 23874 26460 23884 26516
rect 23940 26460 26012 26516
rect 26068 26460 26078 26516
rect 22418 26348 22428 26404
rect 22484 26348 23100 26404
rect 23156 26348 23166 26404
rect 17602 26236 17612 26292
rect 17668 26236 18732 26292
rect 18788 26236 18798 26292
rect 15810 26124 15820 26180
rect 15876 26124 17724 26180
rect 17780 26124 17790 26180
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 4274 25452 4284 25508
rect 4340 25452 13916 25508
rect 13972 25452 13982 25508
rect 13916 25284 13972 25452
rect 18722 25340 18732 25396
rect 18788 25340 25564 25396
rect 25620 25340 27244 25396
rect 27300 25340 27310 25396
rect 13916 25228 16828 25284
rect 16884 25228 16894 25284
rect 24210 25228 24220 25284
rect 24276 25228 25228 25284
rect 25284 25228 25294 25284
rect 26450 25228 26460 25284
rect 26516 25228 27020 25284
rect 27076 25228 27086 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 0 24948 800 24976
rect 41200 24948 42000 24976
rect 0 24892 1932 24948
rect 1988 24892 1998 24948
rect 15138 24892 15148 24948
rect 15204 24892 17612 24948
rect 17668 24892 21420 24948
rect 21476 24892 21486 24948
rect 26898 24892 26908 24948
rect 26964 24892 28588 24948
rect 28644 24892 28654 24948
rect 31892 24892 37660 24948
rect 37716 24892 37726 24948
rect 40002 24892 40012 24948
rect 40068 24892 42000 24948
rect 0 24864 800 24892
rect 31892 24836 31948 24892
rect 41200 24864 42000 24892
rect 28690 24780 28700 24836
rect 28756 24780 31948 24836
rect 15922 24668 15932 24724
rect 15988 24668 16492 24724
rect 16548 24668 18060 24724
rect 18116 24668 18126 24724
rect 18610 24668 18620 24724
rect 18676 24668 20524 24724
rect 20580 24668 20590 24724
rect 31892 24668 37660 24724
rect 37716 24668 37726 24724
rect 31892 24612 31948 24668
rect 18498 24556 18508 24612
rect 18564 24556 21868 24612
rect 21924 24556 21934 24612
rect 22082 24556 22092 24612
rect 22148 24556 22652 24612
rect 22708 24556 25340 24612
rect 25396 24556 25406 24612
rect 27682 24556 27692 24612
rect 27748 24556 28252 24612
rect 28308 24556 31948 24612
rect 22306 24332 22316 24388
rect 22372 24332 26684 24388
rect 26740 24332 26750 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 41200 24276 42000 24304
rect 26114 24220 26124 24276
rect 26180 24220 27916 24276
rect 27972 24220 27982 24276
rect 40002 24220 40012 24276
rect 40068 24220 42000 24276
rect 41200 24192 42000 24220
rect 16146 23996 16156 24052
rect 16212 23996 16828 24052
rect 16884 23996 16894 24052
rect 24882 23996 24892 24052
rect 24948 23996 31948 24052
rect 31892 23940 31948 23996
rect 4274 23884 4284 23940
rect 4340 23884 11452 23940
rect 11508 23884 11518 23940
rect 31892 23884 37660 23940
rect 37716 23884 37726 23940
rect 0 23604 800 23632
rect 41200 23604 42000 23632
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 41200 23520 42000 23548
rect 12002 23436 12012 23492
rect 12068 23436 15596 23492
rect 15652 23436 15662 23492
rect 23090 23436 23100 23492
rect 23156 23436 24892 23492
rect 24948 23436 24958 23492
rect 14130 23324 14140 23380
rect 14196 23324 15484 23380
rect 15540 23324 15550 23380
rect 17154 23324 17164 23380
rect 17220 23324 21980 23380
rect 22036 23324 22046 23380
rect 22754 23324 22764 23380
rect 22820 23324 23660 23380
rect 23716 23324 23726 23380
rect 15586 23212 15596 23268
rect 15652 23212 17332 23268
rect 17602 23212 17612 23268
rect 17668 23212 18172 23268
rect 18228 23212 21196 23268
rect 21252 23212 22652 23268
rect 22708 23212 22718 23268
rect 17276 23156 17332 23212
rect 4274 23100 4284 23156
rect 4340 23100 12012 23156
rect 12068 23100 12078 23156
rect 16146 23100 16156 23156
rect 16212 23100 16828 23156
rect 16884 23100 16894 23156
rect 17266 23100 17276 23156
rect 17332 23100 18620 23156
rect 18676 23100 20972 23156
rect 21028 23100 21038 23156
rect 21298 23100 21308 23156
rect 21364 23100 25228 23156
rect 25284 23100 26012 23156
rect 26068 23100 26078 23156
rect 15810 22988 15820 23044
rect 15876 22988 17836 23044
rect 17892 22988 18060 23044
rect 18116 22988 18126 23044
rect 20514 22988 20524 23044
rect 20580 22988 22372 23044
rect 22978 22988 22988 23044
rect 23044 22988 23772 23044
rect 23828 22988 23838 23044
rect 0 22932 800 22960
rect 0 22876 1932 22932
rect 1988 22876 1998 22932
rect 13794 22876 13804 22932
rect 13860 22876 15036 22932
rect 15092 22876 17388 22932
rect 17444 22876 17454 22932
rect 0 22848 800 22876
rect 20524 22820 20580 22988
rect 22316 22932 22372 22988
rect 22306 22876 22316 22932
rect 22372 22876 22876 22932
rect 22932 22876 22942 22932
rect 15250 22764 15260 22820
rect 15316 22764 16156 22820
rect 16212 22764 20580 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 11442 22316 11452 22372
rect 11508 22316 15036 22372
rect 15092 22316 15102 22372
rect 16706 22316 16716 22372
rect 16772 22316 19180 22372
rect 19236 22316 20076 22372
rect 20132 22316 21420 22372
rect 21476 22316 21486 22372
rect 13570 22092 13580 22148
rect 13636 22092 15372 22148
rect 15428 22092 15438 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 22866 21756 22876 21812
rect 22932 21756 27076 21812
rect 27020 21700 27076 21756
rect 27010 21644 27020 21700
rect 27076 21644 27580 21700
rect 27636 21644 27646 21700
rect 19282 21532 19292 21588
rect 19348 21532 19852 21588
rect 19908 21532 20412 21588
rect 20468 21532 20478 21588
rect 22642 21532 22652 21588
rect 22708 21532 23324 21588
rect 23380 21532 23772 21588
rect 23828 21532 23838 21588
rect 27458 21532 27468 21588
rect 27524 21532 27534 21588
rect 27682 21532 27692 21588
rect 27748 21532 29372 21588
rect 29428 21532 29438 21588
rect 31892 21532 37660 21588
rect 37716 21532 37726 21588
rect 27468 21476 27524 21532
rect 31892 21476 31948 21532
rect 27468 21420 28588 21476
rect 28644 21420 31948 21476
rect 26226 21308 26236 21364
rect 26292 21308 27468 21364
rect 27524 21308 27534 21364
rect 17602 21196 17612 21252
rect 17668 21196 17948 21252
rect 18004 21196 18014 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 41200 20916 42000 20944
rect 18610 20860 18620 20916
rect 18676 20860 19516 20916
rect 19572 20860 19582 20916
rect 40002 20860 40012 20916
rect 40068 20860 42000 20916
rect 41200 20832 42000 20860
rect 4162 20748 4172 20804
rect 4228 20748 20300 20804
rect 20356 20748 21308 20804
rect 21364 20748 21374 20804
rect 8372 20636 10892 20692
rect 10948 20636 14476 20692
rect 14532 20636 14542 20692
rect 8372 20468 8428 20636
rect 17602 20524 17612 20580
rect 17668 20524 19068 20580
rect 19124 20524 19134 20580
rect 20850 20524 20860 20580
rect 20916 20524 24332 20580
rect 24388 20524 25228 20580
rect 25284 20524 25294 20580
rect 4274 20412 4284 20468
rect 4340 20412 8428 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 0 20244 800 20272
rect 0 20188 1932 20244
rect 1988 20188 1998 20244
rect 21634 20188 21644 20244
rect 21700 20188 23100 20244
rect 23156 20188 23166 20244
rect 0 20160 800 20188
rect 14578 20076 14588 20132
rect 14644 20076 15484 20132
rect 15540 20076 15550 20132
rect 17164 20076 20300 20132
rect 20356 20076 20366 20132
rect 21522 20076 21532 20132
rect 21588 20076 22764 20132
rect 22820 20076 23436 20132
rect 23492 20076 23502 20132
rect 17164 20020 17220 20076
rect 15362 19964 15372 20020
rect 15428 19964 17164 20020
rect 17220 19964 17230 20020
rect 19954 19964 19964 20020
rect 20020 19964 20636 20020
rect 20692 19964 21868 20020
rect 21924 19964 21934 20020
rect 14466 19852 14476 19908
rect 14532 19852 15596 19908
rect 15652 19852 15662 19908
rect 17042 19852 17052 19908
rect 17108 19852 17836 19908
rect 17892 19852 17902 19908
rect 18050 19852 18060 19908
rect 18116 19852 20972 19908
rect 21028 19852 21038 19908
rect 23986 19852 23996 19908
rect 24052 19852 25228 19908
rect 25284 19852 25294 19908
rect 12226 19740 12236 19796
rect 12292 19740 14140 19796
rect 14196 19740 14206 19796
rect 16258 19740 16268 19796
rect 16324 19740 17500 19796
rect 17556 19740 17566 19796
rect 18498 19740 18508 19796
rect 18564 19740 19852 19796
rect 19908 19740 23884 19796
rect 23940 19740 23950 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 23426 19404 23436 19460
rect 23492 19404 23884 19460
rect 23940 19404 23950 19460
rect 18162 19292 18172 19348
rect 18228 19292 19404 19348
rect 19460 19292 21196 19348
rect 21252 19292 21262 19348
rect 21970 19292 21980 19348
rect 22036 19292 23996 19348
rect 24052 19292 28140 19348
rect 28196 19292 28206 19348
rect 16482 19180 16492 19236
rect 16548 19180 18732 19236
rect 18788 19180 18798 19236
rect 21410 19180 21420 19236
rect 21476 19180 22092 19236
rect 22148 19180 22158 19236
rect 25442 19180 25452 19236
rect 25508 19180 29036 19236
rect 29092 19180 29102 19236
rect 31892 19180 37660 19236
rect 37716 19180 37726 19236
rect 16258 19068 16268 19124
rect 16324 19068 17388 19124
rect 17444 19068 19516 19124
rect 19572 19068 19582 19124
rect 23762 19068 23772 19124
rect 23828 19068 24332 19124
rect 24388 19068 24398 19124
rect 31892 19012 31948 19180
rect 14466 18956 14476 19012
rect 14532 18956 16380 19012
rect 16436 18956 16446 19012
rect 29250 18956 29260 19012
rect 29316 18956 31948 19012
rect 41200 18900 42000 18928
rect 15698 18844 15708 18900
rect 15764 18844 17836 18900
rect 17892 18844 17902 18900
rect 40002 18844 40012 18900
rect 40068 18844 42000 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 41200 18816 42000 18844
rect 17266 18620 17276 18676
rect 17332 18620 19572 18676
rect 16818 18508 16828 18564
rect 16884 18508 18508 18564
rect 18564 18508 18574 18564
rect 4274 18396 4284 18452
rect 4340 18396 8428 18452
rect 13570 18396 13580 18452
rect 13636 18396 15148 18452
rect 15204 18396 15214 18452
rect 8372 18340 8428 18396
rect 19516 18340 19572 18620
rect 24882 18396 24892 18452
rect 24948 18396 26796 18452
rect 26852 18396 26862 18452
rect 8372 18284 10668 18340
rect 10724 18284 10734 18340
rect 19506 18284 19516 18340
rect 19572 18284 19582 18340
rect 24658 18284 24668 18340
rect 24724 18284 25676 18340
rect 25732 18284 26124 18340
rect 26180 18284 26190 18340
rect 0 18228 800 18256
rect 0 18172 1932 18228
rect 1988 18172 1998 18228
rect 12226 18172 12236 18228
rect 12292 18172 13804 18228
rect 13860 18172 13870 18228
rect 19170 18172 19180 18228
rect 19236 18172 19964 18228
rect 20020 18172 20972 18228
rect 21028 18172 21038 18228
rect 0 18144 800 18172
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 13794 17836 13804 17892
rect 13860 17836 14812 17892
rect 14868 17836 16044 17892
rect 16100 17836 16110 17892
rect 10658 17724 10668 17780
rect 10724 17724 13580 17780
rect 13636 17724 13646 17780
rect 16034 17612 16044 17668
rect 16100 17612 17052 17668
rect 17108 17612 18060 17668
rect 18116 17612 18126 17668
rect 18274 17612 18284 17668
rect 18340 17612 19516 17668
rect 19572 17612 21308 17668
rect 21364 17612 21374 17668
rect 21746 17612 21756 17668
rect 21812 17612 22428 17668
rect 22484 17612 22876 17668
rect 22932 17612 22942 17668
rect 28018 17612 28028 17668
rect 28084 17612 37660 17668
rect 37716 17612 37726 17668
rect 21308 17556 21364 17612
rect 21308 17500 23884 17556
rect 23940 17500 23950 17556
rect 16594 17388 16604 17444
rect 16660 17388 19180 17444
rect 19236 17388 21308 17444
rect 21364 17388 21374 17444
rect 22530 17388 22540 17444
rect 22596 17388 23436 17444
rect 23492 17388 24108 17444
rect 24164 17388 24174 17444
rect 24210 17276 24220 17332
rect 24276 17276 25004 17332
rect 25060 17276 26460 17332
rect 26516 17276 26526 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 16482 17164 16492 17220
rect 16548 17164 17948 17220
rect 18004 17164 19068 17220
rect 19124 17164 19134 17220
rect 16370 17052 16380 17108
rect 16436 17052 17500 17108
rect 17556 17052 18956 17108
rect 19012 17052 19022 17108
rect 23202 17052 23212 17108
rect 23268 17052 24780 17108
rect 24836 17052 25788 17108
rect 25844 17052 25854 17108
rect 15810 16940 15820 16996
rect 15876 16940 25620 16996
rect 26562 16940 26572 16996
rect 26628 16940 28028 16996
rect 28084 16940 28094 16996
rect 25564 16884 25620 16940
rect 41200 16884 42000 16912
rect 15026 16828 15036 16884
rect 15092 16828 17724 16884
rect 17780 16828 17790 16884
rect 24882 16828 24892 16884
rect 24948 16828 25396 16884
rect 25554 16828 25564 16884
rect 25620 16828 25630 16884
rect 40002 16828 40012 16884
rect 40068 16828 42000 16884
rect 19170 16716 19180 16772
rect 19236 16716 20300 16772
rect 20356 16716 21308 16772
rect 21364 16716 21374 16772
rect 25340 16660 25396 16828
rect 41200 16800 42000 16828
rect 25340 16604 25564 16660
rect 25620 16604 25630 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 41200 16212 42000 16240
rect 14242 16156 14252 16212
rect 14308 16156 15484 16212
rect 15540 16156 15550 16212
rect 15922 16156 15932 16212
rect 15988 16156 17164 16212
rect 17220 16156 18060 16212
rect 18116 16156 18126 16212
rect 20850 16156 20860 16212
rect 20916 16156 22092 16212
rect 22148 16156 22652 16212
rect 22708 16156 22718 16212
rect 39890 16156 39900 16212
rect 39956 16156 42000 16212
rect 41200 16128 42000 16156
rect 21298 16044 21308 16100
rect 21364 16044 22204 16100
rect 22260 16044 22270 16100
rect 37650 16044 37660 16100
rect 37716 16044 37726 16100
rect 15810 15932 15820 15988
rect 15876 15932 17388 15988
rect 17444 15932 18396 15988
rect 18452 15932 22540 15988
rect 22596 15932 23324 15988
rect 23380 15932 23390 15988
rect 26562 15932 26572 15988
rect 26628 15932 37436 15988
rect 37492 15932 37502 15988
rect 37660 15876 37716 16044
rect 19058 15820 19068 15876
rect 19124 15820 20188 15876
rect 20244 15820 21644 15876
rect 21700 15820 21710 15876
rect 28242 15820 28252 15876
rect 28308 15820 37716 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 41200 15540 42000 15568
rect 22642 15484 22652 15540
rect 22708 15484 24668 15540
rect 24724 15484 25564 15540
rect 25620 15484 25630 15540
rect 40002 15484 40012 15540
rect 40068 15484 42000 15540
rect 41200 15456 42000 15484
rect 16258 15260 16268 15316
rect 16324 15260 17500 15316
rect 17556 15260 18060 15316
rect 18116 15260 18126 15316
rect 18498 15148 18508 15204
rect 18564 15148 19292 15204
rect 19348 15148 20860 15204
rect 20916 15148 20926 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 17714 14588 17724 14644
rect 17780 14588 18396 14644
rect 18452 14588 18462 14644
rect 22754 14588 22764 14644
rect 22820 14588 23548 14644
rect 23604 14588 23614 14644
rect 21410 14476 21420 14532
rect 21476 14476 22428 14532
rect 22484 14476 22494 14532
rect 21858 14364 21868 14420
rect 21924 14364 23660 14420
rect 23716 14364 24556 14420
rect 24612 14364 24622 14420
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 20178 13804 20188 13860
rect 20244 13804 21532 13860
rect 21588 13804 21598 13860
rect 18610 13468 18620 13524
rect 18676 13468 20076 13524
rect 20132 13468 20142 13524
rect 21746 13468 21756 13524
rect 21812 13468 22652 13524
rect 22708 13468 22718 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 20850 13020 20860 13076
rect 20916 13020 22764 13076
rect 22820 13020 23100 13076
rect 23156 13020 23772 13076
rect 23828 13020 23838 13076
rect 24770 13020 24780 13076
rect 24836 13020 25228 13076
rect 25284 13020 26012 13076
rect 26068 13020 26078 13076
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 23314 11452 23324 11508
rect 23380 11452 24556 11508
rect 24612 11452 24622 11508
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 25666 5180 25676 5236
rect 25732 5180 26796 5236
rect 26852 5180 26862 5236
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 24882 4060 24892 4116
rect 24948 4060 26236 4116
rect 26292 4060 26302 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 22866 3612 22876 3668
rect 22932 3612 25564 3668
rect 25620 3612 25630 3668
rect 20178 3388 20188 3444
rect 20244 3388 21756 3444
rect 21812 3388 21822 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18592 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _107_
timestamp 1698175906
transform -1 0 18144 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16576 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_
timestamp 1698175906
transform 1 0 15232 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17584 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24192 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _112_
timestamp 1698175906
transform -1 0 21728 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_
timestamp 1698175906
transform -1 0 20496 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _114_
timestamp 1698175906
transform -1 0 18816 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22400 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform 1 0 23632 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698175906
transform 1 0 25088 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _119_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _120_
timestamp 1698175906
transform -1 0 16016 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform -1 0 23520 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _122_
timestamp 1698175906
transform 1 0 16016 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1698175906
transform -1 0 23744 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform -1 0 19712 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21280 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _127_
timestamp 1698175906
transform 1 0 22512 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _128_
timestamp 1698175906
transform -1 0 23968 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27440 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _130_
timestamp 1698175906
transform -1 0 19152 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform -1 0 22400 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _132_
timestamp 1698175906
transform -1 0 22288 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _133_
timestamp 1698175906
transform -1 0 21056 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _134_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20608 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _135_
timestamp 1698175906
transform 1 0 25872 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _136_
timestamp 1698175906
transform -1 0 18256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1698175906
transform -1 0 17920 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform 1 0 22288 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _139_
timestamp 1698175906
transform 1 0 24416 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _140_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22288 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _141_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23296 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _142_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16800 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _143_
timestamp 1698175906
transform -1 0 16016 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _144_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19376 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform 1 0 18816 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _146_
timestamp 1698175906
transform -1 0 20832 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _147_
timestamp 1698175906
transform -1 0 20944 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _148_
timestamp 1698175906
transform -1 0 20384 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _149_
timestamp 1698175906
transform 1 0 19824 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _150_
timestamp 1698175906
transform 1 0 20384 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _151_
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _152_
timestamp 1698175906
transform 1 0 15904 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _153_
timestamp 1698175906
transform 1 0 19376 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _154_
timestamp 1698175906
transform -1 0 22288 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _155_
timestamp 1698175906
transform -1 0 21616 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _156_
timestamp 1698175906
transform 1 0 19936 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _157_
timestamp 1698175906
transform -1 0 19936 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _158_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20608 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _159_
timestamp 1698175906
transform -1 0 17024 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _160_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20608 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _161_
timestamp 1698175906
transform 1 0 18704 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _162_
timestamp 1698175906
transform -1 0 17472 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _163_
timestamp 1698175906
transform -1 0 16352 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _164_
timestamp 1698175906
transform -1 0 25200 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _165_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23744 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _166_
timestamp 1698175906
transform 1 0 21952 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _167_
timestamp 1698175906
transform -1 0 23296 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _168_
timestamp 1698175906
transform 1 0 23296 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _169_
timestamp 1698175906
transform -1 0 24752 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _170_
timestamp 1698175906
transform 1 0 16576 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _171_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _172_
timestamp 1698175906
transform -1 0 16016 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _173_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16688 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _174_
timestamp 1698175906
transform -1 0 20272 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _175_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17696 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _176_
timestamp 1698175906
transform -1 0 16576 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _177_
timestamp 1698175906
transform 1 0 14560 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _178_
timestamp 1698175906
transform 1 0 14896 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _179_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18368 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _180_
timestamp 1698175906
transform -1 0 14000 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _181_
timestamp 1698175906
transform -1 0 22064 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _182_
timestamp 1698175906
transform -1 0 23184 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _183_
timestamp 1698175906
transform -1 0 21952 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _184_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22848 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _185_
timestamp 1698175906
transform 1 0 15344 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _186_
timestamp 1698175906
transform 1 0 26320 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _187_
timestamp 1698175906
transform 1 0 25424 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _188_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _189_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18704 0 1 17248
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _190_
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _191_
timestamp 1698175906
transform -1 0 21280 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _192_
timestamp 1698175906
transform -1 0 20608 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _193_
timestamp 1698175906
transform -1 0 19040 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _194_
timestamp 1698175906
transform -1 0 18816 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _195_
timestamp 1698175906
transform 1 0 16128 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _196_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13440 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _197_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14896 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _198_
timestamp 1698175906
transform 1 0 11984 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _199_
timestamp 1698175906
transform 1 0 14336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _200_
timestamp 1698175906
transform -1 0 16128 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _201_
timestamp 1698175906
transform -1 0 14896 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _202_
timestamp 1698175906
transform 1 0 11984 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _203_
timestamp 1698175906
transform -1 0 27776 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _204_
timestamp 1698175906
transform 1 0 23744 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _205_
timestamp 1698175906
transform 1 0 25312 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _206_
timestamp 1698175906
transform -1 0 28896 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _207_
timestamp 1698175906
transform 1 0 21392 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _208_
timestamp 1698175906
transform -1 0 27440 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _209_
timestamp 1698175906
transform 1 0 24192 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _210_
timestamp 1698175906
transform -1 0 29568 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _211_
timestamp 1698175906
transform 1 0 24640 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13888 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 21840 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 25200 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 22960 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 14896 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 19152 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 18368 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 17696 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform -1 0 17024 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 22848 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 21616 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 22960 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform -1 0 15120 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform 1 0 17360 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform -1 0 14560 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 20272 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 25424 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 17248 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform -1 0 13776 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform -1 0 14000 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 25536 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform 1 0 25536 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform 1 0 25872 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _240_
timestamp 1698175906
transform 1 0 27776 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _241_
timestamp 1698175906
transform 1 0 26096 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__B1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16128 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__A2
timestamp 1698175906
transform 1 0 26992 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__C
timestamp 1698175906
transform -1 0 20608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__A2
timestamp 1698175906
transform 1 0 29792 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 17360 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 21616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 25312 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 22736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 18368 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 17696 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 22624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 25872 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 21616 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform -1 0 21168 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 22064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 22064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 22624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 15120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 21392 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 14784 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 23744 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 15120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform 1 0 25648 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 20384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 24864 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform -1 0 24864 0 -1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_154 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_156 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18816 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_161 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19376 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698175906
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_198 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_202
timestamp 1698175906
transform 1 0 23968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 28000 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 31584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_209
timestamp 1698175906
transform 1 0 24752 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_243
timestamp 1698175906
transform 1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_158
timestamp 1698175906
transform 1 0 19040 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_166
timestamp 1698175906
transform 1 0 19936 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_168
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_198
timestamp 1698175906
transform 1 0 23520 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_202
timestamp 1698175906
transform 1 0 23968 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_139
timestamp 1698175906
transform 1 0 16912 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_141
timestamp 1698175906
transform 1 0 17136 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_184
timestamp 1698175906
transform 1 0 21952 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_188
timestamp 1698175906
transform 1 0 22400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_190
timestamp 1698175906
transform 1 0 22624 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_222
timestamp 1698175906
transform 1 0 26208 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_238
timestamp 1698175906
transform 1 0 28000 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_242
timestamp 1698175906
transform 1 0 28448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698175906
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_156
timestamp 1698175906
transform 1 0 18816 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_164
timestamp 1698175906
transform 1 0 19712 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_178
timestamp 1698175906
transform 1 0 21280 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_186
timestamp 1698175906
transform 1 0 22176 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_188
timestamp 1698175906
transform 1 0 22400 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_195
timestamp 1698175906
transform 1 0 23184 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_203
timestamp 1698175906
transform 1 0 24080 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1698175906
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_115
timestamp 1698175906
transform 1 0 14224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_119
timestamp 1698175906
transform 1 0 14672 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_150
timestamp 1698175906
transform 1 0 18144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_154
timestamp 1698175906
transform 1 0 18592 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_170
timestamp 1698175906
transform 1 0 20384 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_185
timestamp 1698175906
transform 1 0 22064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_193
timestamp 1698175906
transform 1 0 22960 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_195
timestamp 1698175906
transform 1 0 23184 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_212
timestamp 1698175906
transform 1 0 25088 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_104
timestamp 1698175906
transform 1 0 12992 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_120
timestamp 1698175906
transform 1 0 14784 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_124
timestamp 1698175906
transform 1 0 15232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698175906
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_154
timestamp 1698175906
transform 1 0 18592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_158
timestamp 1698175906
transform 1 0 19040 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_188
timestamp 1698175906
transform 1 0 22400 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_192
timestamp 1698175906
transform 1 0 22848 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_214
timestamp 1698175906
transform 1 0 25312 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_244
timestamp 1698175906
transform 1 0 28672 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_144
timestamp 1698175906
transform 1 0 17472 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_161
timestamp 1698175906
transform 1 0 19376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698175906
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_181
timestamp 1698175906
transform 1 0 21616 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_227
timestamp 1698175906
transform 1 0 26768 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_235
timestamp 1698175906
transform 1 0 27664 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698175906
transform 1 0 28448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 37296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_104
timestamp 1698175906
transform 1 0 12992 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_120
timestamp 1698175906
transform 1 0 14784 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_124
timestamp 1698175906
transform 1 0 15232 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698175906
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_146
timestamp 1698175906
transform 1 0 17696 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_151
timestamp 1698175906
transform 1 0 18256 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_159
timestamp 1698175906
transform 1 0 19152 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_214
timestamp 1698175906
transform 1 0 25312 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_228
timestamp 1698175906
transform 1 0 26880 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_260
timestamp 1698175906
transform 1 0 30464 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 36512 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 37408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_69
timestamp 1698175906
transform 1 0 9072 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_85
timestamp 1698175906
transform 1 0 10864 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_93
timestamp 1698175906
transform 1 0 11760 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_116
timestamp 1698175906
transform 1 0 14336 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_124
timestamp 1698175906
transform 1 0 15232 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698175906
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_183
timestamp 1698175906
transform 1 0 21840 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_191
timestamp 1698175906
transform 1 0 22736 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_213
timestamp 1698175906
transform 1 0 25200 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_219
timestamp 1698175906
transform 1 0 25872 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_235
timestamp 1698175906
transform 1 0 27664 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698175906
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 4480 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 8064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_80
timestamp 1698175906
transform 1 0 10304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_121
timestamp 1698175906
transform 1 0 14896 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_125
timestamp 1698175906
transform 1 0 15344 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_129
timestamp 1698175906
transform 1 0 15792 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_165
timestamp 1698175906
transform 1 0 19824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_169
timestamp 1698175906
transform 1 0 20272 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_171
timestamp 1698175906
transform 1 0 20496 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_180
timestamp 1698175906
transform 1 0 21504 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_196
timestamp 1698175906
transform 1 0 23296 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_204
timestamp 1698175906
transform 1 0 24192 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_248
timestamp 1698175906
transform 1 0 29120 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 40320 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_69
timestamp 1698175906
transform 1 0 9072 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_85
timestamp 1698175906
transform 1 0 10864 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_93
timestamp 1698175906
transform 1 0 11760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_111
timestamp 1698175906
transform 1 0 13776 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_115
timestamp 1698175906
transform 1 0 14224 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_117
timestamp 1698175906
transform 1 0 14448 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_153
timestamp 1698175906
transform 1 0 18480 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_172
timestamp 1698175906
transform 1 0 20608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698175906
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_187
timestamp 1698175906
transform 1 0 22288 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_195
timestamp 1698175906
transform 1 0 23184 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_199
timestamp 1698175906
transform 1 0 23632 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_252
timestamp 1698175906
transform 1 0 29568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_256
timestamp 1698175906
transform 1 0 30016 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_288
timestamp 1698175906
transform 1 0 33600 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_304
timestamp 1698175906
transform 1 0 35392 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698175906
transform 1 0 36288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698175906
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_80
timestamp 1698175906
transform 1 0 10304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_121
timestamp 1698175906
transform 1 0 14896 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_167
timestamp 1698175906
transform 1 0 20048 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_208
timestamp 1698175906
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_241
timestamp 1698175906
transform 1 0 28336 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_273
timestamp 1698175906
transform 1 0 31920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698175906
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 40320 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698175906
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698175906
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_115
timestamp 1698175906
transform 1 0 14224 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_120
timestamp 1698175906
transform 1 0 14784 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_128
timestamp 1698175906
transform 1 0 15680 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_132
timestamp 1698175906
transform 1 0 16128 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_140
timestamp 1698175906
transform 1 0 17024 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_144
timestamp 1698175906
transform 1 0 17472 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_161
timestamp 1698175906
transform 1 0 19376 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_165
timestamp 1698175906
transform 1 0 19824 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_167
timestamp 1698175906
transform 1 0 20048 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_227
timestamp 1698175906
transform 1 0 26768 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698175906
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_88
timestamp 1698175906
transform 1 0 11200 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_118
timestamp 1698175906
transform 1 0 14560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_122
timestamp 1698175906
transform 1 0 15008 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_138
timestamp 1698175906
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_176
timestamp 1698175906
transform 1 0 21056 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_192
timestamp 1698175906
transform 1 0 22848 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_196
timestamp 1698175906
transform 1 0 23296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_198
timestamp 1698175906
transform 1 0 23520 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_205
timestamp 1698175906
transform 1 0 24304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_217
timestamp 1698175906
transform 1 0 25648 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_221
timestamp 1698175906
transform 1 0 26096 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_236
timestamp 1698175906
transform 1 0 27776 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_268
timestamp 1698175906
transform 1 0 31360 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698175906
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_113
timestamp 1698175906
transform 1 0 14000 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_130
timestamp 1698175906
transform 1 0 15904 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_134
timestamp 1698175906
transform 1 0 16352 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_150
timestamp 1698175906
transform 1 0 18144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_152
timestamp 1698175906
transform 1 0 18368 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_159
timestamp 1698175906
transform 1 0 19152 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_163
timestamp 1698175906
transform 1 0 19600 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_177
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_186
timestamp 1698175906
transform 1 0 22176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_190
timestamp 1698175906
transform 1 0 22624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_198
timestamp 1698175906
transform 1 0 23520 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_230
timestamp 1698175906
transform 1 0 27104 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_238
timestamp 1698175906
transform 1 0 28000 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_242
timestamp 1698175906
transform 1 0 28448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 4480 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_88
timestamp 1698175906
transform 1 0 11200 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_92
timestamp 1698175906
transform 1 0 11648 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_123
timestamp 1698175906
transform 1 0 15120 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_125
timestamp 1698175906
transform 1 0 15344 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698175906
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_152
timestamp 1698175906
transform 1 0 18368 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_168
timestamp 1698175906
transform 1 0 20160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_202
timestamp 1698175906
transform 1 0 23968 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_216
timestamp 1698175906
transform 1 0 25536 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_218
timestamp 1698175906
transform 1 0 25760 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_224
timestamp 1698175906
transform 1 0 26432 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_256
timestamp 1698175906
transform 1 0 30016 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_272
timestamp 1698175906
transform 1 0 31808 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 40320 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_131
timestamp 1698175906
transform 1 0 16016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_144
timestamp 1698175906
transform 1 0 17472 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_155
timestamp 1698175906
transform 1 0 18704 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_163
timestamp 1698175906
transform 1 0 19600 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_169
timestamp 1698175906
transform 1 0 20272 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_173
timestamp 1698175906
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_212
timestamp 1698175906
transform 1 0 25088 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_104
timestamp 1698175906
transform 1 0 12992 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_120
timestamp 1698175906
transform 1 0 14784 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_134
timestamp 1698175906
transform 1 0 16352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_246
timestamp 1698175906
transform 1 0 28896 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698175906
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 36512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 37408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_140
timestamp 1698175906
transform 1 0 17024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_142
timestamp 1698175906
transform 1 0 17248 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698175906
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_181
timestamp 1698175906
transform 1 0 21616 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_197
timestamp 1698175906
transform 1 0 23408 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_205
timestamp 1698175906
transform 1 0 24304 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_209
timestamp 1698175906
transform 1 0 24752 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_211
timestamp 1698175906
transform 1 0 24976 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_218
timestamp 1698175906
transform 1 0 25760 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_222
timestamp 1698175906
transform 1 0 26208 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_224
timestamp 1698175906
transform 1 0 26432 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_238
timestamp 1698175906
transform 1 0 28000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698175906
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_104
timestamp 1698175906
transform 1 0 12992 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_120
timestamp 1698175906
transform 1 0 14784 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_124
timestamp 1698175906
transform 1 0 15232 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_126
timestamp 1698175906
transform 1 0 15456 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_131
timestamp 1698175906
transform 1 0 16016 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_151
timestamp 1698175906
transform 1 0 18256 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_167
timestamp 1698175906
transform 1 0 20048 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_175
timestamp 1698175906
transform 1 0 20944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_177
timestamp 1698175906
transform 1 0 21168 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_187
timestamp 1698175906
transform 1 0 22288 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_189
timestamp 1698175906
transform 1 0 22512 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_111
timestamp 1698175906
transform 1 0 13776 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_141
timestamp 1698175906
transform 1 0 17136 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_145
timestamp 1698175906
transform 1 0 17584 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_161
timestamp 1698175906
transform 1 0 19376 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_181
timestamp 1698175906
transform 1 0 21616 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_183
timestamp 1698175906
transform 1 0 21840 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_222
timestamp 1698175906
transform 1 0 26208 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698175906
transform 1 0 28000 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_150
timestamp 1698175906
transform 1 0 18144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_139
timestamp 1698175906
transform 1 0 16912 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_143
timestamp 1698175906
transform 1 0 17360 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_145
timestamp 1698175906
transform 1 0 17584 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_183
timestamp 1698175906
transform 1 0 21840 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_187
timestamp 1698175906
transform 1 0 22288 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_219
timestamp 1698175906
transform 1 0 25872 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_235
timestamp 1698175906
transform 1 0 27664 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_243
timestamp 1698175906
transform 1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_174
timestamp 1698175906
transform 1 0 20832 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_177
timestamp 1698175906
transform 1 0 21168 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_209
timestamp 1698175906
transform 1 0 24752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_203
timestamp 1698175906
transform 1 0 24080 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_235
timestamp 1698175906
transform 1 0 27664 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_243
timestamp 1698175906
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_6
timestamp 1698175906
transform 1 0 2016 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_174
timestamp 1698175906
transform 1 0 20832 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_201
timestamp 1698175906
transform 1 0 23856 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 25536 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_243
timestamp 1698175906
transform 1 0 28560 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698175906
transform 1 0 32144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_165
timestamp 1698175906
transform 1 0 19824 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_169
timestamp 1698175906
transform 1 0 20272 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_206
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_210
timestamp 1698175906
transform 1 0 24864 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_237
timestamp 1698175906
transform 1 0 27888 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_244
timestamp 1698175906
transform 1 0 28672 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_260
timestamp 1698175906
transform 1 0 30464 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_268
timestamp 1698175906
transform 1 0 31360 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita5_24 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita5_25
timestamp 1698175906
transform -1 0 28672 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita5_26
timestamp 1698175906
transform -1 0 2016 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 4480 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 37520 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 37520 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 25648 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform -1 0 4480 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform -1 0 4480 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 25648 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 24976 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 37520 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 20944 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 21280 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 37520 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 16912 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 41200 24864 42000 24976 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 41200 18816 42000 18928 0 FreeSans 448 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 20160 41200 20272 42000 0 FreeSans 448 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 41200 15456 42000 15568 0 FreeSans 448 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 27552 41200 27664 42000 0 FreeSans 448 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 41200 16800 42000 16912 0 FreeSans 448 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 0 36960 800 37072 0 FreeSans 448 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 25536 41200 25648 42000 0 FreeSans 448 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 24864 41200 24976 42000 0 FreeSans 448 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 41200 16128 42000 16240 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 20832 41200 20944 42000 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 41200 24192 42000 24304 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 16800 41200 16912 42000 0 FreeSans 448 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 23912 13664 23912 13664 0 _000_
rlabel metal3 22960 15960 22960 15960 0 _001_
rlabel metal2 15512 16576 15512 16576 0 _002_
rlabel metal2 20216 15400 20216 15400 0 _003_
rlabel metal2 26040 20888 26040 20888 0 _004_
rlabel metal2 21336 27496 21336 27496 0 _005_
rlabel metal2 19656 27888 19656 27888 0 _006_
rlabel metal2 16072 25144 16072 25144 0 _007_
rlabel metal2 23912 16184 23912 16184 0 _008_
rlabel metal2 22904 27720 22904 27720 0 _009_
rlabel metal2 24192 26936 24192 26936 0 _010_
rlabel metal2 14168 23296 14168 23296 0 _011_
rlabel metal2 18536 24920 18536 24920 0 _012_
rlabel metal2 13664 21672 13664 21672 0 _013_
rlabel metal2 21224 12656 21224 12656 0 _014_
rlabel metal2 26376 15904 26376 15904 0 _015_
rlabel metal2 18256 13048 18256 13048 0 _016_
rlabel metal2 12488 17920 12488 17920 0 _017_
rlabel metal2 12488 19488 12488 19488 0 _018_
rlabel metal2 25816 18872 25816 18872 0 _019_
rlabel metal2 26488 24640 26488 24640 0 _020_
rlabel metal3 25872 18424 25872 18424 0 _021_
rlabel metal2 14840 26712 14840 26712 0 _022_
rlabel metal3 23240 23352 23240 23352 0 _023_
rlabel metal2 26376 23968 26376 23968 0 _024_
rlabel metal3 20104 26936 20104 26936 0 _025_
rlabel metal2 18760 18760 18760 18760 0 _026_
rlabel metal2 15960 24752 15960 24752 0 _027_
rlabel metal2 21336 17920 21336 17920 0 _028_
rlabel metal2 17080 23520 17080 23520 0 _029_
rlabel metal3 16520 24024 16520 24024 0 _030_
rlabel metal2 24584 17640 24584 17640 0 _031_
rlabel metal3 22792 26376 22792 26376 0 _032_
rlabel metal2 24472 26264 24472 26264 0 _033_
rlabel metal2 16184 23464 16184 23464 0 _034_
rlabel metal2 16632 22120 16632 22120 0 _035_
rlabel metal2 16072 23240 16072 23240 0 _036_
rlabel metal2 19992 24360 19992 24360 0 _037_
rlabel metal2 14840 18536 14840 18536 0 _038_
rlabel metal2 27608 21616 27608 21616 0 _039_
rlabel metal3 14504 22120 14504 22120 0 _040_
rlabel metal2 13832 22736 13832 22736 0 _041_
rlabel metal2 21448 14280 21448 14280 0 _042_
rlabel metal2 21784 13328 21784 13328 0 _043_
rlabel metal2 23240 17248 23240 17248 0 _044_
rlabel metal3 25592 16912 25592 16912 0 _045_
rlabel metal2 26320 16856 26320 16856 0 _046_
rlabel metal2 17528 19096 17528 19096 0 _047_
rlabel metal2 17024 17864 17024 17864 0 _048_
rlabel metal2 18984 18312 18984 18312 0 _049_
rlabel metal2 20608 13496 20608 13496 0 _050_
rlabel metal2 18648 12824 18648 12824 0 _051_
rlabel metal2 18368 12376 18368 12376 0 _052_
rlabel metal2 14504 18704 14504 18704 0 _053_
rlabel metal2 14224 17864 14224 17864 0 _054_
rlabel metal2 12264 17920 12264 17920 0 _055_
rlabel metal2 14616 20328 14616 20328 0 _056_
rlabel metal3 15064 19880 15064 19880 0 _057_
rlabel metal2 12264 19488 12264 19488 0 _058_
rlabel metal2 25592 19264 25592 19264 0 _059_
rlabel metal2 25368 18536 25368 18536 0 _060_
rlabel metal3 27776 24920 27776 24920 0 _061_
rlabel metal2 26712 24864 26712 24864 0 _062_
rlabel metal2 24752 19208 24752 19208 0 _063_
rlabel metal3 27272 19208 27272 19208 0 _064_
rlabel metal2 18088 15344 18088 15344 0 _065_
rlabel metal3 21952 23240 21952 23240 0 _066_
rlabel metal2 16072 18816 16072 18816 0 _067_
rlabel metal2 17864 19040 17864 19040 0 _068_
rlabel metal3 20160 26824 20160 26824 0 _069_
rlabel metal3 22176 20104 22176 20104 0 _070_
rlabel metal3 16576 17640 16576 17640 0 _071_
rlabel metal2 19992 17864 19992 17864 0 _072_
rlabel metal2 17864 23296 17864 23296 0 _073_
rlabel metal3 21952 14504 21952 14504 0 _074_
rlabel metal3 23240 21560 23240 21560 0 _075_
rlabel metal2 25032 17416 25032 17416 0 _076_
rlabel metal2 27440 25368 27440 25368 0 _077_
rlabel metal3 16800 26152 16800 26152 0 _078_
rlabel metal3 23016 26936 23016 26936 0 _079_
rlabel metal3 18984 17416 18984 17416 0 _080_
rlabel metal2 21896 22848 21896 22848 0 _081_
rlabel metal2 23688 14336 23688 14336 0 _082_
rlabel metal2 16744 23016 16744 23016 0 _083_
rlabel metal2 22008 22624 22008 22624 0 _084_
rlabel metal3 23408 23016 23408 23016 0 _085_
rlabel metal2 27944 24752 27944 24752 0 _086_
rlabel metal2 18648 22680 18648 22680 0 _087_
rlabel metal2 21896 19656 21896 19656 0 _088_
rlabel metal2 21280 19320 21280 19320 0 _089_
rlabel metal2 21896 26544 21896 26544 0 _090_
rlabel metal3 23688 23128 23688 23128 0 _091_
rlabel metal2 17976 17136 17976 17136 0 _092_
rlabel metal2 22568 16856 22568 16856 0 _093_
rlabel metal2 24360 14728 24360 14728 0 _094_
rlabel metal2 23968 14504 23968 14504 0 _095_
rlabel metal2 15624 16128 15624 16128 0 _096_
rlabel metal3 20944 15848 20944 15848 0 _097_
rlabel metal3 19600 21560 19600 21560 0 _098_
rlabel metal2 17192 21056 17192 21056 0 _099_
rlabel metal3 22960 26488 22960 26488 0 _100_
rlabel metal2 19992 16688 19992 16688 0 _101_
rlabel metal2 24360 20328 24360 20328 0 _102_
rlabel metal2 19544 19264 19544 19264 0 _103_
rlabel metal2 19880 19936 19880 19936 0 _104_
rlabel metal2 21504 26936 21504 26936 0 _105_
rlabel metal3 2478 27608 2478 27608 0 clk
rlabel metal2 23912 22792 23912 22792 0 clknet_0_clk
rlabel metal2 20832 13048 20832 13048 0 clknet_1_0__leaf_clk
rlabel metal2 23072 27048 23072 27048 0 clknet_1_1__leaf_clk
rlabel metal2 18088 14616 18088 14616 0 dut5.count\[0\]
rlabel metal2 16408 16520 16408 16520 0 dut5.count\[1\]
rlabel metal2 20328 18424 20328 18424 0 dut5.count\[2\]
rlabel metal2 28168 19600 28168 19600 0 dut5.count\[3\]
rlabel metal2 12040 23240 12040 23240 0 net1
rlabel metal2 4312 20608 4312 20608 0 net10
rlabel metal2 27496 21616 27496 21616 0 net11
rlabel metal2 26040 32200 26040 32200 0 net12
rlabel metal2 11480 22680 11480 22680 0 net13
rlabel metal2 23352 11760 23352 11760 0 net14
rlabel metal2 24696 28112 24696 28112 0 net15
rlabel metal2 37464 16408 37464 16408 0 net16
rlabel metal2 13944 25536 13944 25536 0 net17
rlabel metal2 20552 27888 20552 27888 0 net18
rlabel metal2 21560 27720 21560 27720 0 net19
rlabel metal2 28672 24024 28672 24024 0 net2
rlabel metal3 25648 13048 25648 13048 0 net20
rlabel metal2 27720 24920 27720 24920 0 net21
rlabel metal2 17136 27160 17136 27160 0 net22
rlabel metal3 31920 23968 31920 23968 0 net23
rlabel metal2 18872 2030 18872 2030 0 net24
rlabel metal2 28392 38248 28392 38248 0 net25
rlabel metal3 1246 37016 1246 37016 0 net26
rlabel metal2 28952 18648 28952 18648 0 net3
rlabel metal2 20272 31920 20272 31920 0 net4
rlabel metal3 37688 15960 37688 15960 0 net5
rlabel metal2 25816 10108 25816 10108 0 net6
rlabel metal2 28056 16856 28056 16856 0 net7
rlabel metal2 20776 5964 20776 5964 0 net8
rlabel metal3 6356 18424 6356 18424 0 net9
rlabel metal3 1358 22904 1358 22904 0 segm[10]
rlabel metal2 40040 25256 40040 25256 0 segm[11]
rlabel metal2 40040 19096 40040 19096 0 segm[12]
rlabel metal2 20216 38962 20216 38962 0 segm[13]
rlabel metal2 40040 15848 40040 15848 0 segm[1]
rlabel metal2 25592 1582 25592 1582 0 segm[2]
rlabel metal2 40040 17304 40040 17304 0 segm[4]
rlabel metal2 20216 2086 20216 2086 0 segm[6]
rlabel metal3 1358 18200 1358 18200 0 segm[7]
rlabel metal3 1358 20216 1358 20216 0 segm[8]
rlabel metal2 40040 21112 40040 21112 0 segm[9]
rlabel metal2 25592 39354 25592 39354 0 sel[0]
rlabel metal3 1358 23576 1358 23576 0 sel[10]
rlabel metal2 22904 2198 22904 2198 0 sel[11]
rlabel metal2 24920 39746 24920 39746 0 sel[1]
rlabel metal2 39928 16464 39928 16464 0 sel[2]
rlabel metal3 1358 24920 1358 24920 0 sel[3]
rlabel metal2 20888 39354 20888 39354 0 sel[4]
rlabel metal2 22232 39746 22232 39746 0 sel[5]
rlabel metal2 24920 2422 24920 2422 0 sel[6]
rlabel metal2 40040 24360 40040 24360 0 sel[7]
rlabel metal2 16856 39746 16856 39746 0 sel[8]
rlabel metal2 40040 23800 40040 23800 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
