magic
tech gf180mcuD
magscale 1 10
timestamp 1699643462
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 19182 38274 19234 38286
rect 19182 38210 19234 38222
rect 26126 38274 26178 38286
rect 26126 38210 26178 38222
rect 22194 38110 22206 38162
rect 22258 38110 22270 38162
rect 19730 37998 19742 38050
rect 19794 37998 19806 38050
rect 23762 37998 23774 38050
rect 23826 37998 23838 38050
rect 25554 37998 25566 38050
rect 25618 37998 25630 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 18398 37490 18450 37502
rect 18398 37426 18450 37438
rect 21422 37490 21474 37502
rect 21422 37426 21474 37438
rect 26798 37490 26850 37502
rect 26798 37426 26850 37438
rect 17378 37214 17390 37266
rect 17442 37214 17454 37266
rect 20402 37214 20414 37266
rect 20466 37214 20478 37266
rect 25890 37214 25902 37266
rect 25954 37214 25966 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 25666 28702 25678 28754
rect 25730 28702 25742 28754
rect 22754 28590 22766 28642
rect 22818 28590 22830 28642
rect 23538 28478 23550 28530
rect 23602 28478 23614 28530
rect 22430 28418 22482 28430
rect 22430 28354 22482 28366
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 19518 28082 19570 28094
rect 19518 28018 19570 28030
rect 25342 28082 25394 28094
rect 25342 28018 25394 28030
rect 18958 27970 19010 27982
rect 18958 27906 19010 27918
rect 19070 27858 19122 27870
rect 19070 27794 19122 27806
rect 19294 27858 19346 27870
rect 19294 27794 19346 27806
rect 19630 27858 19682 27870
rect 23326 27858 23378 27870
rect 20066 27806 20078 27858
rect 20130 27806 20142 27858
rect 19630 27794 19682 27806
rect 23326 27794 23378 27806
rect 23550 27858 23602 27870
rect 23550 27794 23602 27806
rect 23998 27858 24050 27870
rect 23998 27794 24050 27806
rect 25118 27858 25170 27870
rect 25118 27794 25170 27806
rect 25454 27858 25506 27870
rect 25454 27794 25506 27806
rect 23438 27746 23490 27758
rect 20738 27694 20750 27746
rect 20802 27694 20814 27746
rect 22866 27694 22878 27746
rect 22930 27694 22942 27746
rect 23438 27682 23490 27694
rect 24334 27746 24386 27758
rect 24334 27682 24386 27694
rect 18958 27634 19010 27646
rect 18958 27570 19010 27582
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 1934 27186 1986 27198
rect 18050 27134 18062 27186
rect 18114 27134 18126 27186
rect 20178 27134 20190 27186
rect 20242 27134 20254 27186
rect 23762 27134 23774 27186
rect 23826 27134 23838 27186
rect 25890 27134 25902 27186
rect 25954 27134 25966 27186
rect 1934 27122 1986 27134
rect 20638 27074 20690 27086
rect 4274 27022 4286 27074
rect 4338 27022 4350 27074
rect 17378 27022 17390 27074
rect 17442 27022 17454 27074
rect 20638 27010 20690 27022
rect 21198 27074 21250 27086
rect 21198 27010 21250 27022
rect 22654 27074 22706 27086
rect 23090 27022 23102 27074
rect 23154 27022 23166 27074
rect 22654 27010 22706 27022
rect 21422 26962 21474 26974
rect 21422 26898 21474 26910
rect 21534 26962 21586 26974
rect 21534 26898 21586 26910
rect 21758 26962 21810 26974
rect 21758 26898 21810 26910
rect 21982 26962 22034 26974
rect 21982 26898 22034 26910
rect 22094 26962 22146 26974
rect 22094 26898 22146 26910
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 20750 26514 20802 26526
rect 20750 26450 20802 26462
rect 22430 26514 22482 26526
rect 22430 26450 22482 26462
rect 23102 26514 23154 26526
rect 23102 26450 23154 26462
rect 25118 26514 25170 26526
rect 25118 26450 25170 26462
rect 25342 26514 25394 26526
rect 25342 26450 25394 26462
rect 22206 26402 22258 26414
rect 22206 26338 22258 26350
rect 22094 26290 22146 26302
rect 4274 26238 4286 26290
rect 4338 26238 4350 26290
rect 13906 26238 13918 26290
rect 13970 26238 13982 26290
rect 17490 26238 17502 26290
rect 17554 26238 17566 26290
rect 22094 26226 22146 26238
rect 23326 26290 23378 26302
rect 23326 26226 23378 26238
rect 23774 26290 23826 26302
rect 23774 26226 23826 26238
rect 25454 26290 25506 26302
rect 25454 26226 25506 26238
rect 23214 26178 23266 26190
rect 14690 26126 14702 26178
rect 14754 26126 14766 26178
rect 16818 26126 16830 26178
rect 16882 26126 16894 26178
rect 18162 26126 18174 26178
rect 18226 26126 18238 26178
rect 20290 26126 20302 26178
rect 20354 26126 20366 26178
rect 23214 26114 23266 26126
rect 1934 26066 1986 26078
rect 1934 26002 1986 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 15822 25730 15874 25742
rect 22430 25730 22482 25742
rect 17490 25678 17502 25730
rect 17554 25727 17566 25730
rect 18050 25727 18062 25730
rect 17554 25681 18062 25727
rect 17554 25678 17566 25681
rect 18050 25678 18062 25681
rect 18114 25678 18126 25730
rect 15822 25666 15874 25678
rect 22430 25666 22482 25678
rect 2034 25566 2046 25618
rect 2098 25566 2110 25618
rect 13682 25566 13694 25618
rect 13746 25566 13758 25618
rect 16606 25506 16658 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 12786 25454 12798 25506
rect 12850 25454 12862 25506
rect 14578 25454 14590 25506
rect 14642 25454 14654 25506
rect 16606 25442 16658 25454
rect 16942 25506 16994 25518
rect 18286 25506 18338 25518
rect 17154 25454 17166 25506
rect 17218 25454 17230 25506
rect 16942 25442 16994 25454
rect 18286 25442 18338 25454
rect 19518 25506 19570 25518
rect 19518 25442 19570 25454
rect 14030 25394 14082 25406
rect 15934 25394 15986 25406
rect 12562 25342 12574 25394
rect 12626 25342 12638 25394
rect 14354 25342 14366 25394
rect 14418 25342 14430 25394
rect 14030 25330 14082 25342
rect 15934 25330 15986 25342
rect 16830 25394 16882 25406
rect 16830 25330 16882 25342
rect 17726 25394 17778 25406
rect 17726 25330 17778 25342
rect 18622 25394 18674 25406
rect 18622 25330 18674 25342
rect 19182 25394 19234 25406
rect 19182 25330 19234 25342
rect 19406 25394 19458 25406
rect 22318 25394 22370 25406
rect 21634 25342 21646 25394
rect 21698 25342 21710 25394
rect 19406 25330 19458 25342
rect 22318 25330 22370 25342
rect 13806 25282 13858 25294
rect 13806 25218 13858 25230
rect 16718 25282 16770 25294
rect 16718 25218 16770 25230
rect 18062 25282 18114 25294
rect 18062 25218 18114 25230
rect 18510 25282 18562 25294
rect 18510 25218 18562 25230
rect 21982 25282 22034 25294
rect 21982 25218 22034 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 14814 24946 14866 24958
rect 14814 24882 14866 24894
rect 24110 24834 24162 24846
rect 13570 24782 13582 24834
rect 13634 24782 13646 24834
rect 23650 24782 23662 24834
rect 23714 24782 23726 24834
rect 24110 24770 24162 24782
rect 23326 24722 23378 24734
rect 14242 24670 14254 24722
rect 14306 24670 14318 24722
rect 21858 24670 21870 24722
rect 21922 24670 21934 24722
rect 23326 24658 23378 24670
rect 24222 24722 24274 24734
rect 37650 24670 37662 24722
rect 37714 24670 37726 24722
rect 24222 24658 24274 24670
rect 15486 24610 15538 24622
rect 11442 24558 11454 24610
rect 11506 24558 11518 24610
rect 14690 24558 14702 24610
rect 14754 24558 14766 24610
rect 15486 24546 15538 24558
rect 22318 24610 22370 24622
rect 22318 24546 22370 24558
rect 24670 24610 24722 24622
rect 24670 24546 24722 24558
rect 15038 24498 15090 24510
rect 15038 24434 15090 24446
rect 24110 24498 24162 24510
rect 24110 24434 24162 24446
rect 40014 24498 40066 24510
rect 40014 24434 40066 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 40014 24050 40066 24062
rect 24770 23998 24782 24050
rect 24834 23998 24846 24050
rect 28354 23998 28366 24050
rect 28418 23998 28430 24050
rect 40014 23986 40066 23998
rect 20526 23938 20578 23950
rect 20526 23874 20578 23886
rect 21534 23938 21586 23950
rect 21858 23886 21870 23938
rect 21922 23886 21934 23938
rect 25442 23886 25454 23938
rect 25506 23886 25518 23938
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 21534 23874 21586 23886
rect 22642 23774 22654 23826
rect 22706 23774 22718 23826
rect 26226 23774 26238 23826
rect 26290 23774 26302 23826
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 14366 23378 14418 23390
rect 14366 23314 14418 23326
rect 25790 23378 25842 23390
rect 25790 23314 25842 23326
rect 26686 23378 26738 23390
rect 26686 23314 26738 23326
rect 16606 23266 16658 23278
rect 16606 23202 16658 23214
rect 17950 23266 18002 23278
rect 17950 23202 18002 23214
rect 26574 23266 26626 23278
rect 26574 23202 26626 23214
rect 14814 23154 14866 23166
rect 4274 23102 4286 23154
rect 4338 23102 4350 23154
rect 13906 23102 13918 23154
rect 13970 23102 13982 23154
rect 14814 23090 14866 23102
rect 15150 23154 15202 23166
rect 15150 23090 15202 23102
rect 15374 23154 15426 23166
rect 15374 23090 15426 23102
rect 16494 23154 16546 23166
rect 16494 23090 16546 23102
rect 16830 23154 16882 23166
rect 16830 23090 16882 23102
rect 17838 23154 17890 23166
rect 17838 23090 17890 23102
rect 18174 23154 18226 23166
rect 25678 23154 25730 23166
rect 22978 23102 22990 23154
rect 23042 23102 23054 23154
rect 18174 23090 18226 23102
rect 25678 23090 25730 23102
rect 25902 23154 25954 23166
rect 25902 23090 25954 23102
rect 26350 23154 26402 23166
rect 26350 23090 26402 23102
rect 14926 23042 14978 23054
rect 10994 22990 11006 23042
rect 11058 22990 11070 23042
rect 13122 22990 13134 23042
rect 13186 22990 13198 23042
rect 14926 22978 14978 22990
rect 17502 23042 17554 23054
rect 25342 23042 25394 23054
rect 21746 22990 21758 23042
rect 21810 22990 21822 23042
rect 17502 22978 17554 22990
rect 25342 22978 25394 22990
rect 1934 22930 1986 22942
rect 1934 22866 1986 22878
rect 26686 22930 26738 22942
rect 26686 22866 26738 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 13694 22482 13746 22494
rect 22766 22482 22818 22494
rect 14914 22430 14926 22482
rect 14978 22430 14990 22482
rect 17042 22430 17054 22482
rect 17106 22430 17118 22482
rect 18162 22430 18174 22482
rect 18226 22430 18238 22482
rect 20290 22430 20302 22482
rect 20354 22430 20366 22482
rect 13694 22418 13746 22430
rect 22766 22418 22818 22430
rect 24334 22482 24386 22494
rect 40014 22482 40066 22494
rect 28242 22430 28254 22482
rect 28306 22430 28318 22482
rect 24334 22418 24386 22430
rect 40014 22418 40066 22430
rect 23326 22370 23378 22382
rect 14130 22318 14142 22370
rect 14194 22318 14206 22370
rect 17490 22318 17502 22370
rect 17554 22318 17566 22370
rect 21522 22318 21534 22370
rect 21586 22318 21598 22370
rect 23326 22306 23378 22318
rect 23550 22370 23602 22382
rect 23550 22306 23602 22318
rect 23886 22370 23938 22382
rect 24658 22318 24670 22370
rect 24722 22318 24734 22370
rect 25330 22318 25342 22370
rect 25394 22318 25406 22370
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 23886 22306 23938 22318
rect 20750 22258 20802 22270
rect 20750 22194 20802 22206
rect 22654 22258 22706 22270
rect 22654 22194 22706 22206
rect 23662 22258 23714 22270
rect 23662 22194 23714 22206
rect 24894 22258 24946 22270
rect 24894 22194 24946 22206
rect 25006 22258 25058 22270
rect 26114 22206 26126 22258
rect 26178 22206 26190 22258
rect 25006 22194 25058 22206
rect 20638 22146 20690 22158
rect 21982 22146 22034 22158
rect 22878 22146 22930 22158
rect 21298 22094 21310 22146
rect 21362 22094 21374 22146
rect 22306 22094 22318 22146
rect 22370 22094 22382 22146
rect 20638 22082 20690 22094
rect 21982 22082 22034 22094
rect 22878 22082 22930 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 14142 21810 14194 21822
rect 14142 21746 14194 21758
rect 14814 21810 14866 21822
rect 14814 21746 14866 21758
rect 15486 21810 15538 21822
rect 26126 21810 26178 21822
rect 16482 21758 16494 21810
rect 16546 21758 16558 21810
rect 15486 21746 15538 21758
rect 26126 21746 26178 21758
rect 14590 21698 14642 21710
rect 14590 21634 14642 21646
rect 15934 21698 15986 21710
rect 18174 21698 18226 21710
rect 26238 21698 26290 21710
rect 17378 21646 17390 21698
rect 17442 21646 17454 21698
rect 22978 21646 22990 21698
rect 23042 21646 23054 21698
rect 15934 21634 15986 21646
rect 18174 21634 18226 21646
rect 26238 21634 26290 21646
rect 13918 21586 13970 21598
rect 4274 21534 4286 21586
rect 4338 21534 4350 21586
rect 13458 21534 13470 21586
rect 13522 21534 13534 21586
rect 13918 21522 13970 21534
rect 14142 21586 14194 21598
rect 14142 21522 14194 21534
rect 14478 21586 14530 21598
rect 14478 21522 14530 21534
rect 14926 21586 14978 21598
rect 14926 21522 14978 21534
rect 15374 21586 15426 21598
rect 15374 21522 15426 21534
rect 15710 21586 15762 21598
rect 17726 21586 17778 21598
rect 16706 21534 16718 21586
rect 16770 21534 16782 21586
rect 15710 21522 15762 21534
rect 17726 21522 17778 21534
rect 19070 21586 19122 21598
rect 25678 21586 25730 21598
rect 19394 21534 19406 21586
rect 19458 21534 19470 21586
rect 19070 21522 19122 21534
rect 25678 21522 25730 21534
rect 26014 21586 26066 21598
rect 26014 21522 26066 21534
rect 10546 21422 10558 21474
rect 10610 21422 10622 21474
rect 12674 21422 12686 21474
rect 12738 21422 12750 21474
rect 18610 21422 18622 21474
rect 18674 21422 18686 21474
rect 1934 21362 1986 21374
rect 1934 21298 1986 21310
rect 18062 21362 18114 21374
rect 18062 21298 18114 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 12350 21026 12402 21038
rect 12350 20962 12402 20974
rect 20750 21026 20802 21038
rect 24222 21026 24274 21038
rect 22194 20974 22206 21026
rect 22258 20974 22270 21026
rect 20750 20962 20802 20974
rect 24222 20962 24274 20974
rect 12238 20914 12290 20926
rect 19182 20914 19234 20926
rect 23886 20914 23938 20926
rect 14130 20862 14142 20914
rect 14194 20862 14206 20914
rect 21858 20862 21870 20914
rect 21922 20862 21934 20914
rect 12238 20850 12290 20862
rect 19182 20850 19234 20862
rect 23886 20850 23938 20862
rect 14478 20802 14530 20814
rect 14478 20738 14530 20750
rect 20078 20802 20130 20814
rect 21410 20750 21422 20802
rect 21474 20750 21486 20802
rect 22306 20750 22318 20802
rect 22370 20750 22382 20802
rect 23202 20750 23214 20802
rect 23266 20750 23278 20802
rect 20078 20738 20130 20750
rect 14142 20690 14194 20702
rect 14018 20638 14030 20690
rect 14082 20638 14094 20690
rect 14142 20626 14194 20638
rect 14254 20690 14306 20702
rect 14254 20626 14306 20638
rect 20414 20690 20466 20702
rect 20414 20626 20466 20638
rect 20638 20690 20690 20702
rect 22978 20638 22990 20690
rect 23042 20638 23054 20690
rect 20638 20626 20690 20638
rect 24110 20578 24162 20590
rect 19730 20526 19742 20578
rect 19794 20526 19806 20578
rect 24110 20514 24162 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 14254 20242 14306 20254
rect 14254 20178 14306 20190
rect 18062 20242 18114 20254
rect 23202 20190 23214 20242
rect 23266 20190 23278 20242
rect 18062 20178 18114 20190
rect 18734 20130 18786 20142
rect 15698 20078 15710 20130
rect 15762 20078 15774 20130
rect 17714 20078 17726 20130
rect 17778 20078 17790 20130
rect 18386 20078 18398 20130
rect 18450 20078 18462 20130
rect 18734 20066 18786 20078
rect 20414 20130 20466 20142
rect 20414 20066 20466 20078
rect 20862 20130 20914 20142
rect 20862 20066 20914 20078
rect 21198 20130 21250 20142
rect 21198 20066 21250 20078
rect 21646 20130 21698 20142
rect 27694 20130 27746 20142
rect 23762 20078 23774 20130
rect 23826 20078 23838 20130
rect 26338 20078 26350 20130
rect 26402 20078 26414 20130
rect 21646 20066 21698 20078
rect 27694 20066 27746 20078
rect 16046 20018 16098 20030
rect 13682 19966 13694 20018
rect 13746 19966 13758 20018
rect 16046 19954 16098 19966
rect 21870 20018 21922 20030
rect 26014 20018 26066 20030
rect 22978 19966 22990 20018
rect 23042 19966 23054 20018
rect 23986 19966 23998 20018
rect 24050 19966 24062 20018
rect 21870 19954 21922 19966
rect 26014 19954 26066 19966
rect 26574 20018 26626 20030
rect 26574 19954 26626 19966
rect 26910 20018 26962 20030
rect 26910 19954 26962 19966
rect 27246 20018 27298 20030
rect 27246 19954 27298 19966
rect 27582 20018 27634 20030
rect 27582 19954 27634 19966
rect 27918 20018 27970 20030
rect 27918 19954 27970 19966
rect 28030 20018 28082 20030
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 28030 19954 28082 19966
rect 22206 19906 22258 19918
rect 10882 19854 10894 19906
rect 10946 19854 10958 19906
rect 13010 19854 13022 19906
rect 13074 19854 13086 19906
rect 20514 19854 20526 19906
rect 20578 19854 20590 19906
rect 21522 19854 21534 19906
rect 21586 19854 21598 19906
rect 22206 19842 22258 19854
rect 26798 19906 26850 19918
rect 26798 19842 26850 19854
rect 20190 19794 20242 19806
rect 20190 19730 20242 19742
rect 22318 19794 22370 19806
rect 22318 19730 22370 19742
rect 40014 19794 40066 19806
rect 40014 19730 40066 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 22094 19458 22146 19470
rect 22094 19394 22146 19406
rect 23662 19458 23714 19470
rect 23662 19394 23714 19406
rect 1934 19346 1986 19358
rect 1934 19282 1986 19294
rect 13806 19346 13858 19358
rect 40014 19346 40066 19358
rect 20290 19294 20302 19346
rect 20354 19294 20366 19346
rect 26450 19294 26462 19346
rect 26514 19294 26526 19346
rect 28578 19294 28590 19346
rect 28642 19294 28654 19346
rect 13806 19282 13858 19294
rect 40014 19282 40066 19294
rect 13918 19234 13970 19246
rect 4274 19182 4286 19234
rect 4338 19182 4350 19234
rect 13918 19170 13970 19182
rect 14254 19234 14306 19246
rect 14254 19170 14306 19182
rect 16494 19234 16546 19246
rect 16494 19170 16546 19182
rect 20638 19234 20690 19246
rect 23326 19234 23378 19246
rect 21522 19182 21534 19234
rect 21586 19182 21598 19234
rect 22194 19182 22206 19234
rect 22258 19182 22270 19234
rect 22530 19182 22542 19234
rect 22594 19182 22606 19234
rect 23090 19182 23102 19234
rect 23154 19182 23166 19234
rect 20638 19170 20690 19182
rect 23326 19170 23378 19182
rect 23550 19234 23602 19246
rect 25666 19182 25678 19234
rect 25730 19182 25742 19234
rect 29250 19182 29262 19234
rect 29314 19182 29326 19234
rect 37650 19182 37662 19234
rect 37714 19182 37726 19234
rect 23550 19170 23602 19182
rect 13694 19122 13746 19134
rect 15362 19070 15374 19122
rect 15426 19070 15438 19122
rect 16146 19070 16158 19122
rect 16210 19070 16222 19122
rect 21410 19070 21422 19122
rect 21474 19070 21486 19122
rect 13694 19058 13746 19070
rect 14702 19010 14754 19022
rect 14702 18946 14754 18958
rect 15710 19010 15762 19022
rect 15710 18946 15762 18958
rect 20078 19010 20130 19022
rect 20078 18946 20130 18958
rect 20302 19010 20354 19022
rect 20302 18946 20354 18958
rect 25342 19010 25394 19022
rect 29474 18958 29486 19010
rect 29538 18958 29550 19010
rect 25342 18946 25394 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 14702 18674 14754 18686
rect 14702 18610 14754 18622
rect 14814 18674 14866 18686
rect 14814 18610 14866 18622
rect 18622 18674 18674 18686
rect 25902 18674 25954 18686
rect 21746 18622 21758 18674
rect 21810 18622 21822 18674
rect 18622 18610 18674 18622
rect 25902 18610 25954 18622
rect 14926 18562 14978 18574
rect 13570 18510 13582 18562
rect 13634 18510 13646 18562
rect 14926 18498 14978 18510
rect 15822 18562 15874 18574
rect 15822 18498 15874 18510
rect 18510 18562 18562 18574
rect 21422 18562 21474 18574
rect 22766 18562 22818 18574
rect 19618 18510 19630 18562
rect 19682 18510 19694 18562
rect 22418 18510 22430 18562
rect 22482 18510 22494 18562
rect 18510 18498 18562 18510
rect 21422 18498 21474 18510
rect 22766 18498 22818 18510
rect 23550 18562 23602 18574
rect 23550 18498 23602 18510
rect 15374 18450 15426 18462
rect 4274 18398 4286 18450
rect 4338 18398 4350 18450
rect 14354 18398 14366 18450
rect 14418 18398 14430 18450
rect 15374 18386 15426 18398
rect 16046 18450 16098 18462
rect 16046 18386 16098 18398
rect 16158 18450 16210 18462
rect 16158 18386 16210 18398
rect 16270 18450 16322 18462
rect 20302 18450 20354 18462
rect 19954 18398 19966 18450
rect 20018 18398 20030 18450
rect 16270 18386 16322 18398
rect 20302 18386 20354 18398
rect 20750 18450 20802 18462
rect 20750 18386 20802 18398
rect 21198 18450 21250 18462
rect 21198 18386 21250 18398
rect 22094 18450 22146 18462
rect 23438 18450 23490 18462
rect 23090 18398 23102 18450
rect 23154 18398 23166 18450
rect 22094 18386 22146 18398
rect 23438 18386 23490 18398
rect 23774 18450 23826 18462
rect 25678 18450 25730 18462
rect 25442 18398 25454 18450
rect 25506 18398 25518 18450
rect 23774 18386 23826 18398
rect 25678 18386 25730 18398
rect 25790 18450 25842 18462
rect 26114 18398 26126 18450
rect 26178 18398 26190 18450
rect 26450 18398 26462 18450
rect 26514 18398 26526 18450
rect 27234 18398 27246 18450
rect 27298 18398 27310 18450
rect 37874 18398 37886 18450
rect 37938 18398 37950 18450
rect 25790 18386 25842 18398
rect 20526 18338 20578 18350
rect 11442 18286 11454 18338
rect 11506 18286 11518 18338
rect 19282 18286 19294 18338
rect 19346 18286 19358 18338
rect 20526 18274 20578 18286
rect 24670 18338 24722 18350
rect 29362 18286 29374 18338
rect 29426 18286 29438 18338
rect 24670 18274 24722 18286
rect 1934 18226 1986 18238
rect 1934 18162 1986 18174
rect 18622 18226 18674 18238
rect 18622 18162 18674 18174
rect 23102 18226 23154 18238
rect 23102 18162 23154 18174
rect 40014 18226 40066 18238
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 14590 17890 14642 17902
rect 14018 17838 14030 17890
rect 14082 17838 14094 17890
rect 14590 17826 14642 17838
rect 14926 17890 14978 17902
rect 14926 17826 14978 17838
rect 13582 17778 13634 17790
rect 13582 17714 13634 17726
rect 40014 17778 40066 17790
rect 40014 17714 40066 17726
rect 13806 17666 13858 17678
rect 18510 17666 18562 17678
rect 27022 17666 27074 17678
rect 14018 17614 14030 17666
rect 14082 17614 14094 17666
rect 16706 17614 16718 17666
rect 16770 17614 16782 17666
rect 17154 17614 17166 17666
rect 17218 17614 17230 17666
rect 22754 17614 22766 17666
rect 22818 17614 22830 17666
rect 13806 17602 13858 17614
rect 18510 17602 18562 17614
rect 27022 17602 27074 17614
rect 27358 17666 27410 17678
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 27358 17602 27410 17614
rect 13470 17554 13522 17566
rect 13470 17490 13522 17502
rect 14702 17554 14754 17566
rect 14702 17490 14754 17502
rect 17278 17554 17330 17566
rect 27246 17554 27298 17566
rect 18162 17502 18174 17554
rect 18226 17502 18238 17554
rect 19282 17502 19294 17554
rect 19346 17502 19358 17554
rect 20402 17502 20414 17554
rect 20466 17502 20478 17554
rect 24658 17502 24670 17554
rect 24722 17502 24734 17554
rect 17278 17490 17330 17502
rect 27246 17490 27298 17502
rect 17838 17442 17890 17454
rect 19630 17442 19682 17454
rect 18834 17390 18846 17442
rect 18898 17390 18910 17442
rect 17838 17378 17890 17390
rect 19630 17378 19682 17390
rect 20078 17442 20130 17454
rect 20078 17378 20130 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 18510 17106 18562 17118
rect 18510 17042 18562 17054
rect 20302 17106 20354 17118
rect 20302 17042 20354 17054
rect 21086 17106 21138 17118
rect 21086 17042 21138 17054
rect 21982 17106 22034 17118
rect 21982 17042 22034 17054
rect 22990 17106 23042 17118
rect 22990 17042 23042 17054
rect 23102 17106 23154 17118
rect 23102 17042 23154 17054
rect 24334 17106 24386 17118
rect 24334 17042 24386 17054
rect 26462 17106 26514 17118
rect 26462 17042 26514 17054
rect 20862 16994 20914 17006
rect 14690 16942 14702 16994
rect 14754 16942 14766 16994
rect 20862 16930 20914 16942
rect 22094 16994 22146 17006
rect 22094 16930 22146 16942
rect 24222 16994 24274 17006
rect 24222 16930 24274 16942
rect 25230 16994 25282 17006
rect 25230 16930 25282 16942
rect 25342 16994 25394 17006
rect 25342 16930 25394 16942
rect 18398 16882 18450 16894
rect 14018 16830 14030 16882
rect 14082 16830 14094 16882
rect 17714 16830 17726 16882
rect 17778 16830 17790 16882
rect 18398 16818 18450 16830
rect 20414 16882 20466 16894
rect 20414 16818 20466 16830
rect 21310 16882 21362 16894
rect 21310 16818 21362 16830
rect 22654 16882 22706 16894
rect 22654 16818 22706 16830
rect 22766 16882 22818 16894
rect 22766 16818 22818 16830
rect 23998 16882 24050 16894
rect 23998 16818 24050 16830
rect 24670 16882 24722 16894
rect 24670 16818 24722 16830
rect 25566 16882 25618 16894
rect 25566 16818 25618 16830
rect 17390 16770 17442 16782
rect 16818 16718 16830 16770
rect 16882 16718 16894 16770
rect 17390 16706 17442 16718
rect 17502 16770 17554 16782
rect 17502 16706 17554 16718
rect 21198 16770 21250 16782
rect 21198 16706 21250 16718
rect 22878 16770 22930 16782
rect 22878 16706 22930 16718
rect 20302 16658 20354 16670
rect 20302 16594 20354 16606
rect 21982 16658 22034 16670
rect 21982 16594 22034 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 22542 16322 22594 16334
rect 22542 16258 22594 16270
rect 27134 16210 27186 16222
rect 24098 16158 24110 16210
rect 24162 16158 24174 16210
rect 26226 16158 26238 16210
rect 26290 16158 26302 16210
rect 27134 16146 27186 16158
rect 40014 16210 40066 16222
rect 40014 16146 40066 16158
rect 19854 16098 19906 16110
rect 19854 16034 19906 16046
rect 20078 16098 20130 16110
rect 22430 16098 22482 16110
rect 26910 16098 26962 16110
rect 22082 16046 22094 16098
rect 22146 16046 22158 16098
rect 23426 16046 23438 16098
rect 23490 16046 23502 16098
rect 26674 16046 26686 16098
rect 26738 16046 26750 16098
rect 37650 16046 37662 16098
rect 37714 16046 37726 16098
rect 20078 16034 20130 16046
rect 22430 16034 22482 16046
rect 26910 16034 26962 16046
rect 20302 15986 20354 15998
rect 20302 15922 20354 15934
rect 21534 15986 21586 15998
rect 21534 15922 21586 15934
rect 21646 15986 21698 15998
rect 21646 15922 21698 15934
rect 22542 15986 22594 15998
rect 22542 15922 22594 15934
rect 27246 15986 27298 15998
rect 27246 15922 27298 15934
rect 17054 15874 17106 15886
rect 17054 15810 17106 15822
rect 19966 15874 20018 15886
rect 19966 15810 20018 15822
rect 21310 15874 21362 15886
rect 21310 15810 21362 15822
rect 21422 15874 21474 15886
rect 21422 15810 21474 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 21534 15538 21586 15550
rect 21534 15474 21586 15486
rect 21646 15538 21698 15550
rect 21646 15474 21698 15486
rect 21870 15538 21922 15550
rect 21870 15474 21922 15486
rect 27122 15374 27134 15426
rect 27186 15374 27198 15426
rect 20526 15314 20578 15326
rect 20526 15250 20578 15262
rect 20750 15314 20802 15326
rect 26014 15314 26066 15326
rect 22082 15262 22094 15314
rect 22146 15262 22158 15314
rect 26450 15262 26462 15314
rect 26514 15262 26526 15314
rect 20750 15250 20802 15262
rect 26014 15250 26066 15262
rect 18062 15202 18114 15214
rect 18062 15138 18114 15150
rect 21758 15202 21810 15214
rect 29250 15150 29262 15202
rect 29314 15150 29326 15202
rect 21758 15138 21810 15150
rect 21074 15038 21086 15090
rect 21138 15038 21150 15090
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 22878 14754 22930 14766
rect 22878 14690 22930 14702
rect 26462 14754 26514 14766
rect 26462 14690 26514 14702
rect 18734 14642 18786 14654
rect 17266 14590 17278 14642
rect 17330 14590 17342 14642
rect 18734 14578 18786 14590
rect 26126 14642 26178 14654
rect 26126 14578 26178 14590
rect 27694 14642 27746 14654
rect 27694 14578 27746 14590
rect 40014 14642 40066 14654
rect 40014 14578 40066 14590
rect 16494 14530 16546 14542
rect 17614 14530 17666 14542
rect 17154 14478 17166 14530
rect 17218 14478 17230 14530
rect 16494 14466 16546 14478
rect 17614 14466 17666 14478
rect 17726 14530 17778 14542
rect 17726 14466 17778 14478
rect 18510 14530 18562 14542
rect 18510 14466 18562 14478
rect 21870 14530 21922 14542
rect 21870 14466 21922 14478
rect 22094 14530 22146 14542
rect 22094 14466 22146 14478
rect 22542 14530 22594 14542
rect 22542 14466 22594 14478
rect 22766 14530 22818 14542
rect 22766 14466 22818 14478
rect 26238 14530 26290 14542
rect 26238 14466 26290 14478
rect 27022 14530 27074 14542
rect 27234 14478 27246 14530
rect 27298 14478 27310 14530
rect 27906 14478 27918 14530
rect 27970 14478 27982 14530
rect 37650 14478 37662 14530
rect 37714 14478 37726 14530
rect 27022 14466 27074 14478
rect 26910 14418 26962 14430
rect 26910 14354 26962 14366
rect 27582 14418 27634 14430
rect 27582 14354 27634 14366
rect 16382 14306 16434 14318
rect 16382 14242 16434 14254
rect 17390 14306 17442 14318
rect 21982 14306 22034 14318
rect 18162 14254 18174 14306
rect 18226 14254 18238 14306
rect 17390 14242 17442 14254
rect 21982 14242 22034 14254
rect 22878 14306 22930 14318
rect 22878 14242 22930 14254
rect 23438 14306 23490 14318
rect 23438 14242 23490 14254
rect 26126 14306 26178 14318
rect 26126 14242 26178 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 17502 13970 17554 13982
rect 17502 13906 17554 13918
rect 23662 13970 23714 13982
rect 23662 13906 23714 13918
rect 24334 13970 24386 13982
rect 24334 13906 24386 13918
rect 24670 13970 24722 13982
rect 24670 13906 24722 13918
rect 17838 13858 17890 13870
rect 14690 13806 14702 13858
rect 14754 13806 14766 13858
rect 17838 13794 17890 13806
rect 18174 13858 18226 13870
rect 21074 13806 21086 13858
rect 21138 13806 21150 13858
rect 26114 13806 26126 13858
rect 26178 13806 26190 13858
rect 18174 13794 18226 13806
rect 23438 13746 23490 13758
rect 14018 13694 14030 13746
rect 14082 13694 14094 13746
rect 20290 13694 20302 13746
rect 20354 13694 20366 13746
rect 23438 13682 23490 13694
rect 23774 13746 23826 13758
rect 25330 13694 25342 13746
rect 25394 13694 25406 13746
rect 23774 13682 23826 13694
rect 16818 13582 16830 13634
rect 16882 13582 16894 13634
rect 23202 13582 23214 13634
rect 23266 13582 23278 13634
rect 28242 13582 28254 13634
rect 28306 13582 28318 13634
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 20302 13074 20354 13086
rect 24782 13074 24834 13086
rect 17602 13022 17614 13074
rect 17666 13022 17678 13074
rect 19730 13022 19742 13074
rect 19794 13022 19806 13074
rect 22082 13022 22094 13074
rect 22146 13022 22158 13074
rect 24210 13022 24222 13074
rect 24274 13022 24286 13074
rect 20302 13010 20354 13022
rect 24782 13010 24834 13022
rect 16930 12910 16942 12962
rect 16994 12910 17006 12962
rect 21298 12910 21310 12962
rect 21362 12910 21374 12962
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 19070 4450 19122 4462
rect 19070 4386 19122 4398
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 18622 3666 18674 3678
rect 18622 3602 18674 3614
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 17938 3502 17950 3554
rect 18002 3502 18014 3554
rect 23538 3502 23550 3554
rect 23602 3502 23614 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 22194 3390 22206 3442
rect 22258 3390 22270 3442
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 19182 38222 19234 38274
rect 26126 38222 26178 38274
rect 22206 38110 22258 38162
rect 19742 37998 19794 38050
rect 23774 37998 23826 38050
rect 25566 37998 25618 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 18398 37438 18450 37490
rect 21422 37438 21474 37490
rect 26798 37438 26850 37490
rect 17390 37214 17442 37266
rect 20414 37214 20466 37266
rect 25902 37214 25954 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 25678 28702 25730 28754
rect 22766 28590 22818 28642
rect 23550 28478 23602 28530
rect 22430 28366 22482 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 19518 28030 19570 28082
rect 25342 28030 25394 28082
rect 18958 27918 19010 27970
rect 19070 27806 19122 27858
rect 19294 27806 19346 27858
rect 19630 27806 19682 27858
rect 20078 27806 20130 27858
rect 23326 27806 23378 27858
rect 23550 27806 23602 27858
rect 23998 27806 24050 27858
rect 25118 27806 25170 27858
rect 25454 27806 25506 27858
rect 20750 27694 20802 27746
rect 22878 27694 22930 27746
rect 23438 27694 23490 27746
rect 24334 27694 24386 27746
rect 18958 27582 19010 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 1934 27134 1986 27186
rect 18062 27134 18114 27186
rect 20190 27134 20242 27186
rect 23774 27134 23826 27186
rect 25902 27134 25954 27186
rect 4286 27022 4338 27074
rect 17390 27022 17442 27074
rect 20638 27022 20690 27074
rect 21198 27022 21250 27074
rect 22654 27022 22706 27074
rect 23102 27022 23154 27074
rect 21422 26910 21474 26962
rect 21534 26910 21586 26962
rect 21758 26910 21810 26962
rect 21982 26910 22034 26962
rect 22094 26910 22146 26962
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 20750 26462 20802 26514
rect 22430 26462 22482 26514
rect 23102 26462 23154 26514
rect 25118 26462 25170 26514
rect 25342 26462 25394 26514
rect 22206 26350 22258 26402
rect 4286 26238 4338 26290
rect 13918 26238 13970 26290
rect 17502 26238 17554 26290
rect 22094 26238 22146 26290
rect 23326 26238 23378 26290
rect 23774 26238 23826 26290
rect 25454 26238 25506 26290
rect 14702 26126 14754 26178
rect 16830 26126 16882 26178
rect 18174 26126 18226 26178
rect 20302 26126 20354 26178
rect 23214 26126 23266 26178
rect 1934 26014 1986 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 15822 25678 15874 25730
rect 17502 25678 17554 25730
rect 18062 25678 18114 25730
rect 22430 25678 22482 25730
rect 2046 25566 2098 25618
rect 13694 25566 13746 25618
rect 4286 25454 4338 25506
rect 12798 25454 12850 25506
rect 14590 25454 14642 25506
rect 16606 25454 16658 25506
rect 16942 25454 16994 25506
rect 17166 25454 17218 25506
rect 18286 25454 18338 25506
rect 19518 25454 19570 25506
rect 12574 25342 12626 25394
rect 14030 25342 14082 25394
rect 14366 25342 14418 25394
rect 15934 25342 15986 25394
rect 16830 25342 16882 25394
rect 17726 25342 17778 25394
rect 18622 25342 18674 25394
rect 19182 25342 19234 25394
rect 19406 25342 19458 25394
rect 21646 25342 21698 25394
rect 22318 25342 22370 25394
rect 13806 25230 13858 25282
rect 16718 25230 16770 25282
rect 18062 25230 18114 25282
rect 18510 25230 18562 25282
rect 21982 25230 22034 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 14814 24894 14866 24946
rect 13582 24782 13634 24834
rect 23662 24782 23714 24834
rect 24110 24782 24162 24834
rect 14254 24670 14306 24722
rect 21870 24670 21922 24722
rect 23326 24670 23378 24722
rect 24222 24670 24274 24722
rect 37662 24670 37714 24722
rect 11454 24558 11506 24610
rect 14702 24558 14754 24610
rect 15486 24558 15538 24610
rect 22318 24558 22370 24610
rect 24670 24558 24722 24610
rect 15038 24446 15090 24498
rect 24110 24446 24162 24498
rect 40014 24446 40066 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 24782 23998 24834 24050
rect 28366 23998 28418 24050
rect 40014 23998 40066 24050
rect 20526 23886 20578 23938
rect 21534 23886 21586 23938
rect 21870 23886 21922 23938
rect 25454 23886 25506 23938
rect 37662 23886 37714 23938
rect 22654 23774 22706 23826
rect 26238 23774 26290 23826
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 14366 23326 14418 23378
rect 25790 23326 25842 23378
rect 26686 23326 26738 23378
rect 16606 23214 16658 23266
rect 17950 23214 18002 23266
rect 26574 23214 26626 23266
rect 4286 23102 4338 23154
rect 13918 23102 13970 23154
rect 14814 23102 14866 23154
rect 15150 23102 15202 23154
rect 15374 23102 15426 23154
rect 16494 23102 16546 23154
rect 16830 23102 16882 23154
rect 17838 23102 17890 23154
rect 18174 23102 18226 23154
rect 22990 23102 23042 23154
rect 25678 23102 25730 23154
rect 25902 23102 25954 23154
rect 26350 23102 26402 23154
rect 11006 22990 11058 23042
rect 13134 22990 13186 23042
rect 14926 22990 14978 23042
rect 17502 22990 17554 23042
rect 21758 22990 21810 23042
rect 25342 22990 25394 23042
rect 1934 22878 1986 22930
rect 26686 22878 26738 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 13694 22430 13746 22482
rect 14926 22430 14978 22482
rect 17054 22430 17106 22482
rect 18174 22430 18226 22482
rect 20302 22430 20354 22482
rect 22766 22430 22818 22482
rect 24334 22430 24386 22482
rect 28254 22430 28306 22482
rect 40014 22430 40066 22482
rect 14142 22318 14194 22370
rect 17502 22318 17554 22370
rect 21534 22318 21586 22370
rect 23326 22318 23378 22370
rect 23550 22318 23602 22370
rect 23886 22318 23938 22370
rect 24670 22318 24722 22370
rect 25342 22318 25394 22370
rect 37662 22318 37714 22370
rect 20750 22206 20802 22258
rect 22654 22206 22706 22258
rect 23662 22206 23714 22258
rect 24894 22206 24946 22258
rect 25006 22206 25058 22258
rect 26126 22206 26178 22258
rect 20638 22094 20690 22146
rect 21310 22094 21362 22146
rect 21982 22094 22034 22146
rect 22318 22094 22370 22146
rect 22878 22094 22930 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 14142 21758 14194 21810
rect 14814 21758 14866 21810
rect 15486 21758 15538 21810
rect 16494 21758 16546 21810
rect 26126 21758 26178 21810
rect 14590 21646 14642 21698
rect 15934 21646 15986 21698
rect 17390 21646 17442 21698
rect 18174 21646 18226 21698
rect 22990 21646 23042 21698
rect 26238 21646 26290 21698
rect 4286 21534 4338 21586
rect 13470 21534 13522 21586
rect 13918 21534 13970 21586
rect 14142 21534 14194 21586
rect 14478 21534 14530 21586
rect 14926 21534 14978 21586
rect 15374 21534 15426 21586
rect 15710 21534 15762 21586
rect 16718 21534 16770 21586
rect 17726 21534 17778 21586
rect 19070 21534 19122 21586
rect 19406 21534 19458 21586
rect 25678 21534 25730 21586
rect 26014 21534 26066 21586
rect 10558 21422 10610 21474
rect 12686 21422 12738 21474
rect 18622 21422 18674 21474
rect 1934 21310 1986 21362
rect 18062 21310 18114 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 12350 20974 12402 21026
rect 20750 20974 20802 21026
rect 22206 20974 22258 21026
rect 24222 20974 24274 21026
rect 12238 20862 12290 20914
rect 14142 20862 14194 20914
rect 19182 20862 19234 20914
rect 21870 20862 21922 20914
rect 23886 20862 23938 20914
rect 14478 20750 14530 20802
rect 20078 20750 20130 20802
rect 21422 20750 21474 20802
rect 22318 20750 22370 20802
rect 23214 20750 23266 20802
rect 14030 20638 14082 20690
rect 14142 20638 14194 20690
rect 14254 20638 14306 20690
rect 20414 20638 20466 20690
rect 20638 20638 20690 20690
rect 22990 20638 23042 20690
rect 19742 20526 19794 20578
rect 24110 20526 24162 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 14254 20190 14306 20242
rect 18062 20190 18114 20242
rect 23214 20190 23266 20242
rect 15710 20078 15762 20130
rect 17726 20078 17778 20130
rect 18398 20078 18450 20130
rect 18734 20078 18786 20130
rect 20414 20078 20466 20130
rect 20862 20078 20914 20130
rect 21198 20078 21250 20130
rect 21646 20078 21698 20130
rect 23774 20078 23826 20130
rect 26350 20078 26402 20130
rect 27694 20078 27746 20130
rect 13694 19966 13746 20018
rect 16046 19966 16098 20018
rect 21870 19966 21922 20018
rect 22990 19966 23042 20018
rect 23998 19966 24050 20018
rect 26014 19966 26066 20018
rect 26574 19966 26626 20018
rect 26910 19966 26962 20018
rect 27246 19966 27298 20018
rect 27582 19966 27634 20018
rect 27918 19966 27970 20018
rect 28030 19966 28082 20018
rect 37662 19966 37714 20018
rect 10894 19854 10946 19906
rect 13022 19854 13074 19906
rect 20526 19854 20578 19906
rect 21534 19854 21586 19906
rect 22206 19854 22258 19906
rect 26798 19854 26850 19906
rect 20190 19742 20242 19794
rect 22318 19742 22370 19794
rect 40014 19742 40066 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 22094 19406 22146 19458
rect 23662 19406 23714 19458
rect 1934 19294 1986 19346
rect 13806 19294 13858 19346
rect 20302 19294 20354 19346
rect 26462 19294 26514 19346
rect 28590 19294 28642 19346
rect 40014 19294 40066 19346
rect 4286 19182 4338 19234
rect 13918 19182 13970 19234
rect 14254 19182 14306 19234
rect 16494 19182 16546 19234
rect 20638 19182 20690 19234
rect 21534 19182 21586 19234
rect 22206 19182 22258 19234
rect 22542 19182 22594 19234
rect 23102 19182 23154 19234
rect 23326 19182 23378 19234
rect 23550 19182 23602 19234
rect 25678 19182 25730 19234
rect 29262 19182 29314 19234
rect 37662 19182 37714 19234
rect 13694 19070 13746 19122
rect 15374 19070 15426 19122
rect 16158 19070 16210 19122
rect 21422 19070 21474 19122
rect 14702 18958 14754 19010
rect 15710 18958 15762 19010
rect 20078 18958 20130 19010
rect 20302 18958 20354 19010
rect 25342 18958 25394 19010
rect 29486 18958 29538 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 14702 18622 14754 18674
rect 14814 18622 14866 18674
rect 18622 18622 18674 18674
rect 21758 18622 21810 18674
rect 25902 18622 25954 18674
rect 13582 18510 13634 18562
rect 14926 18510 14978 18562
rect 15822 18510 15874 18562
rect 18510 18510 18562 18562
rect 19630 18510 19682 18562
rect 21422 18510 21474 18562
rect 22430 18510 22482 18562
rect 22766 18510 22818 18562
rect 23550 18510 23602 18562
rect 4286 18398 4338 18450
rect 14366 18398 14418 18450
rect 15374 18398 15426 18450
rect 16046 18398 16098 18450
rect 16158 18398 16210 18450
rect 16270 18398 16322 18450
rect 19966 18398 20018 18450
rect 20302 18398 20354 18450
rect 20750 18398 20802 18450
rect 21198 18398 21250 18450
rect 22094 18398 22146 18450
rect 23102 18398 23154 18450
rect 23438 18398 23490 18450
rect 23774 18398 23826 18450
rect 25454 18398 25506 18450
rect 25678 18398 25730 18450
rect 25790 18398 25842 18450
rect 26126 18398 26178 18450
rect 26462 18398 26514 18450
rect 27246 18398 27298 18450
rect 37886 18398 37938 18450
rect 11454 18286 11506 18338
rect 19294 18286 19346 18338
rect 20526 18286 20578 18338
rect 24670 18286 24722 18338
rect 29374 18286 29426 18338
rect 1934 18174 1986 18226
rect 18622 18174 18674 18226
rect 23102 18174 23154 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 14030 17838 14082 17890
rect 14590 17838 14642 17890
rect 14926 17838 14978 17890
rect 13582 17726 13634 17778
rect 40014 17726 40066 17778
rect 13806 17614 13858 17666
rect 14030 17614 14082 17666
rect 16718 17614 16770 17666
rect 17166 17614 17218 17666
rect 18510 17614 18562 17666
rect 22766 17614 22818 17666
rect 27022 17614 27074 17666
rect 27358 17614 27410 17666
rect 37662 17614 37714 17666
rect 13470 17502 13522 17554
rect 14702 17502 14754 17554
rect 17278 17502 17330 17554
rect 18174 17502 18226 17554
rect 19294 17502 19346 17554
rect 20414 17502 20466 17554
rect 24670 17502 24722 17554
rect 27246 17502 27298 17554
rect 17838 17390 17890 17442
rect 18846 17390 18898 17442
rect 19630 17390 19682 17442
rect 20078 17390 20130 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 18510 17054 18562 17106
rect 20302 17054 20354 17106
rect 21086 17054 21138 17106
rect 21982 17054 22034 17106
rect 22990 17054 23042 17106
rect 23102 17054 23154 17106
rect 24334 17054 24386 17106
rect 26462 17054 26514 17106
rect 14702 16942 14754 16994
rect 20862 16942 20914 16994
rect 22094 16942 22146 16994
rect 24222 16942 24274 16994
rect 25230 16942 25282 16994
rect 25342 16942 25394 16994
rect 14030 16830 14082 16882
rect 17726 16830 17778 16882
rect 18398 16830 18450 16882
rect 20414 16830 20466 16882
rect 21310 16830 21362 16882
rect 22654 16830 22706 16882
rect 22766 16830 22818 16882
rect 23998 16830 24050 16882
rect 24670 16830 24722 16882
rect 25566 16830 25618 16882
rect 16830 16718 16882 16770
rect 17390 16718 17442 16770
rect 17502 16718 17554 16770
rect 21198 16718 21250 16770
rect 22878 16718 22930 16770
rect 20302 16606 20354 16658
rect 21982 16606 22034 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 22542 16270 22594 16322
rect 24110 16158 24162 16210
rect 26238 16158 26290 16210
rect 27134 16158 27186 16210
rect 40014 16158 40066 16210
rect 19854 16046 19906 16098
rect 20078 16046 20130 16098
rect 22094 16046 22146 16098
rect 22430 16046 22482 16098
rect 23438 16046 23490 16098
rect 26686 16046 26738 16098
rect 26910 16046 26962 16098
rect 37662 16046 37714 16098
rect 20302 15934 20354 15986
rect 21534 15934 21586 15986
rect 21646 15934 21698 15986
rect 22542 15934 22594 15986
rect 27246 15934 27298 15986
rect 17054 15822 17106 15874
rect 19966 15822 20018 15874
rect 21310 15822 21362 15874
rect 21422 15822 21474 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 21534 15486 21586 15538
rect 21646 15486 21698 15538
rect 21870 15486 21922 15538
rect 27134 15374 27186 15426
rect 20526 15262 20578 15314
rect 20750 15262 20802 15314
rect 22094 15262 22146 15314
rect 26014 15262 26066 15314
rect 26462 15262 26514 15314
rect 18062 15150 18114 15202
rect 21758 15150 21810 15202
rect 29262 15150 29314 15202
rect 21086 15038 21138 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 22878 14702 22930 14754
rect 26462 14702 26514 14754
rect 17278 14590 17330 14642
rect 18734 14590 18786 14642
rect 26126 14590 26178 14642
rect 27694 14590 27746 14642
rect 40014 14590 40066 14642
rect 16494 14478 16546 14530
rect 17166 14478 17218 14530
rect 17614 14478 17666 14530
rect 17726 14478 17778 14530
rect 18510 14478 18562 14530
rect 21870 14478 21922 14530
rect 22094 14478 22146 14530
rect 22542 14478 22594 14530
rect 22766 14478 22818 14530
rect 26238 14478 26290 14530
rect 27022 14478 27074 14530
rect 27246 14478 27298 14530
rect 27918 14478 27970 14530
rect 37662 14478 37714 14530
rect 26910 14366 26962 14418
rect 27582 14366 27634 14418
rect 16382 14254 16434 14306
rect 17390 14254 17442 14306
rect 18174 14254 18226 14306
rect 21982 14254 22034 14306
rect 22878 14254 22930 14306
rect 23438 14254 23490 14306
rect 26126 14254 26178 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 17502 13918 17554 13970
rect 23662 13918 23714 13970
rect 24334 13918 24386 13970
rect 24670 13918 24722 13970
rect 14702 13806 14754 13858
rect 17838 13806 17890 13858
rect 18174 13806 18226 13858
rect 21086 13806 21138 13858
rect 26126 13806 26178 13858
rect 14030 13694 14082 13746
rect 20302 13694 20354 13746
rect 23438 13694 23490 13746
rect 23774 13694 23826 13746
rect 25342 13694 25394 13746
rect 16830 13582 16882 13634
rect 23214 13582 23266 13634
rect 28254 13582 28306 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 17614 13022 17666 13074
rect 19742 13022 19794 13074
rect 20302 13022 20354 13074
rect 22094 13022 22146 13074
rect 24222 13022 24274 13074
rect 24782 13022 24834 13074
rect 16942 12910 16994 12962
rect 21310 12910 21362 12962
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 19070 4398 19122 4450
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18622 3614 18674 3666
rect 25566 3614 25618 3666
rect 17950 3502 18002 3554
rect 23550 3502 23602 3554
rect 24558 3502 24610 3554
rect 22206 3390 22258 3442
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 16800 41200 16912 42000
rect 19488 41200 19600 42000
rect 20160 41200 20272 42000
rect 22176 41200 22288 42000
rect 24864 41200 24976 42000
rect 25536 41200 25648 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 16828 37492 16884 41200
rect 19180 38276 19236 38286
rect 19516 38276 19572 41200
rect 19180 38274 19572 38276
rect 19180 38222 19182 38274
rect 19234 38222 19572 38274
rect 19180 38220 19572 38222
rect 19180 38210 19236 38220
rect 19740 38052 19796 38062
rect 19404 38050 19796 38052
rect 19404 37998 19742 38050
rect 19794 37998 19796 38050
rect 19404 37996 19796 37998
rect 16828 37426 16884 37436
rect 18396 37492 18452 37502
rect 18396 37398 18452 37436
rect 17388 37266 17444 37278
rect 17388 37214 17390 37266
rect 17442 37214 17444 37266
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 17388 31948 17444 37214
rect 16828 31892 17444 31948
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4172 27636 4228 27646
rect 1932 27186 1988 27198
rect 1932 27134 1934 27186
rect 1986 27134 1988 27186
rect 1932 26292 1988 27134
rect 1932 26226 1988 26236
rect 1932 26066 1988 26078
rect 1932 26014 1934 26066
rect 1986 26014 1988 26066
rect 1932 25620 1988 26014
rect 1932 25554 1988 25564
rect 2044 25618 2100 25630
rect 2044 25566 2046 25618
rect 2098 25566 2100 25618
rect 2044 24948 2100 25566
rect 2044 24882 2100 24892
rect 1932 22932 1988 22942
rect 1932 22838 1988 22876
rect 1932 21362 1988 21374
rect 1932 21310 1934 21362
rect 1986 21310 1988 21362
rect 1932 20916 1988 21310
rect 1932 20850 1988 20860
rect 4172 20580 4228 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4284 27076 4340 27086
rect 4284 26982 4340 27020
rect 14364 27076 14420 27086
rect 4284 26292 4340 26302
rect 4284 26198 4340 26236
rect 12572 26292 12628 26302
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4284 25508 4340 25518
rect 4284 25414 4340 25452
rect 11452 25508 11508 25518
rect 11452 24610 11508 25452
rect 12572 25394 12628 26236
rect 13916 26290 13972 26302
rect 13916 26238 13918 26290
rect 13970 26238 13972 26290
rect 13692 25620 13748 25630
rect 13580 25618 13748 25620
rect 13580 25566 13694 25618
rect 13746 25566 13748 25618
rect 13580 25564 13748 25566
rect 12796 25508 12852 25518
rect 12796 25414 12852 25452
rect 12572 25342 12574 25394
rect 12626 25342 12628 25394
rect 12572 25330 12628 25342
rect 13580 24834 13636 25564
rect 13692 25554 13748 25564
rect 13804 25284 13860 25294
rect 13804 25190 13860 25228
rect 13580 24782 13582 24834
rect 13634 24782 13636 24834
rect 13580 24770 13636 24782
rect 13916 24724 13972 26238
rect 14028 25396 14084 25406
rect 14028 25394 14196 25396
rect 14028 25342 14030 25394
rect 14082 25342 14196 25394
rect 14028 25340 14196 25342
rect 14028 25330 14084 25340
rect 14140 25060 14196 25340
rect 14364 25394 14420 27020
rect 16604 26404 16660 26414
rect 14700 26180 14756 26190
rect 14700 26086 14756 26124
rect 15820 26180 15876 26190
rect 15820 25730 15876 26124
rect 15820 25678 15822 25730
rect 15874 25678 15876 25730
rect 15820 25666 15876 25678
rect 14588 25508 14644 25518
rect 16604 25508 16660 26348
rect 16828 26180 16884 31892
rect 18956 27972 19012 27982
rect 18844 27970 19012 27972
rect 18844 27918 18958 27970
rect 19010 27918 19012 27970
rect 18844 27916 19012 27918
rect 18060 27636 18116 27646
rect 18060 27186 18116 27580
rect 18060 27134 18062 27186
rect 18114 27134 18116 27186
rect 18060 27122 18116 27134
rect 17388 27076 17444 27086
rect 17388 27074 17556 27076
rect 17388 27022 17390 27074
rect 17442 27022 17556 27074
rect 17388 27020 17556 27022
rect 17388 27010 17444 27020
rect 17500 26290 17556 27020
rect 18844 26908 18900 27916
rect 18956 27906 19012 27916
rect 19068 27860 19124 27870
rect 19292 27860 19348 27870
rect 19068 27858 19348 27860
rect 19068 27806 19070 27858
rect 19122 27806 19294 27858
rect 19346 27806 19348 27858
rect 19068 27804 19348 27806
rect 19068 27794 19124 27804
rect 19292 27794 19348 27804
rect 18956 27636 19012 27646
rect 18956 27542 19012 27580
rect 18844 26852 19348 26908
rect 17500 26238 17502 26290
rect 17554 26238 17556 26290
rect 16828 26178 16996 26180
rect 16828 26126 16830 26178
rect 16882 26126 16996 26178
rect 16828 26124 16996 26126
rect 16828 26114 16884 26124
rect 14644 25452 14868 25508
rect 14588 25414 14644 25452
rect 14364 25342 14366 25394
rect 14418 25342 14420 25394
rect 14364 25330 14420 25342
rect 14140 25004 14756 25060
rect 14252 24724 14308 24734
rect 13916 24722 14308 24724
rect 13916 24670 14254 24722
rect 14306 24670 14308 24722
rect 13916 24668 14308 24670
rect 11452 24558 11454 24610
rect 11506 24558 11508 24610
rect 11452 24546 11508 24558
rect 14252 24612 14308 24668
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 14252 23380 14308 24556
rect 14700 24610 14756 25004
rect 14812 24946 14868 25452
rect 16380 25506 16660 25508
rect 16380 25454 16606 25506
rect 16658 25454 16660 25506
rect 16380 25452 16660 25454
rect 15932 25396 15988 25406
rect 15932 25302 15988 25340
rect 14812 24894 14814 24946
rect 14866 24894 14868 24946
rect 14812 24882 14868 24894
rect 14700 24558 14702 24610
rect 14754 24558 14756 24610
rect 14700 24546 14756 24558
rect 15484 24612 15540 24622
rect 15484 24518 15540 24556
rect 15036 24498 15092 24510
rect 15036 24446 15038 24498
rect 15090 24446 15092 24498
rect 14364 23380 14420 23390
rect 13916 23378 14420 23380
rect 13916 23326 14366 23378
rect 14418 23326 14420 23378
rect 13916 23324 14420 23326
rect 4284 23156 4340 23166
rect 4284 23062 4340 23100
rect 11004 23156 11060 23166
rect 13916 23156 13972 23324
rect 11004 23042 11060 23100
rect 13692 23154 13972 23156
rect 13692 23102 13918 23154
rect 13970 23102 13972 23154
rect 13692 23100 13972 23102
rect 11004 22990 11006 23042
rect 11058 22990 11060 23042
rect 11004 22978 11060 22990
rect 13132 23042 13188 23054
rect 13132 22990 13134 23042
rect 13186 22990 13188 23042
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 13132 21812 13188 22990
rect 13692 22484 13748 23100
rect 13916 23090 13972 23100
rect 13132 21746 13188 21756
rect 13468 22482 13748 22484
rect 13468 22430 13694 22482
rect 13746 22430 13748 22482
rect 13468 22428 13748 22430
rect 4284 21588 4340 21598
rect 4284 21494 4340 21532
rect 10556 21588 10612 21598
rect 10556 21474 10612 21532
rect 13468 21588 13524 22428
rect 13692 22418 13748 22428
rect 14028 23044 14084 23054
rect 14028 21812 14084 22988
rect 14140 22370 14196 23324
rect 14364 23314 14420 23324
rect 14476 23156 14532 23166
rect 14812 23156 14868 23166
rect 14532 23100 14756 23156
rect 14476 23090 14532 23100
rect 14364 22372 14420 22382
rect 14140 22318 14142 22370
rect 14194 22318 14196 22370
rect 14140 22306 14196 22318
rect 14252 22316 14364 22372
rect 13916 21756 14084 21812
rect 14140 21812 14196 21822
rect 13468 21586 13748 21588
rect 13468 21534 13470 21586
rect 13522 21534 13748 21586
rect 13468 21532 13748 21534
rect 13468 21522 13524 21532
rect 12684 21476 12740 21486
rect 10556 21422 10558 21474
rect 10610 21422 10612 21474
rect 10556 21410 10612 21422
rect 12348 21474 12740 21476
rect 12348 21422 12686 21474
rect 12738 21422 12740 21474
rect 12348 21420 12740 21422
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 12348 21026 12404 21420
rect 12684 21410 12740 21420
rect 12348 20974 12350 21026
rect 12402 20974 12404 21026
rect 12348 20962 12404 20974
rect 12236 20916 12292 20926
rect 12236 20822 12292 20860
rect 4172 20514 4228 20524
rect 13692 20244 13748 21532
rect 13692 20018 13748 20188
rect 13692 19966 13694 20018
rect 13746 19966 13748 20018
rect 13692 19954 13748 19966
rect 13916 21586 13972 21756
rect 14140 21718 14196 21756
rect 13916 21534 13918 21586
rect 13970 21534 13972 21586
rect 10892 19906 10948 19918
rect 10892 19854 10894 19906
rect 10946 19854 10948 19906
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 1932 19346 1988 19358
rect 1932 19294 1934 19346
rect 1986 19294 1988 19346
rect 1932 18900 1988 19294
rect 4284 19236 4340 19246
rect 4284 19142 4340 19180
rect 1932 18834 1988 18844
rect 4284 18452 4340 18462
rect 4284 18358 4340 18396
rect 10892 18452 10948 19854
rect 13020 19906 13076 19918
rect 13020 19854 13022 19906
rect 13074 19854 13076 19906
rect 10892 18386 10948 18396
rect 11452 19236 11508 19246
rect 11452 18564 11508 19180
rect 11452 18338 11508 18508
rect 11452 18286 11454 18338
rect 11506 18286 11508 18338
rect 11452 18274 11508 18286
rect 1932 18228 1988 18238
rect 1932 18134 1988 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 13020 17780 13076 19854
rect 13804 19348 13860 19358
rect 13468 19346 13860 19348
rect 13468 19294 13806 19346
rect 13858 19294 13860 19346
rect 13468 19292 13860 19294
rect 13468 18564 13524 19292
rect 13804 19282 13860 19292
rect 13916 19236 13972 21534
rect 14140 21588 14196 21598
rect 14252 21588 14308 22316
rect 14364 22306 14420 22316
rect 14700 21812 14756 23100
rect 14812 23062 14868 23100
rect 14924 23042 14980 23054
rect 14924 22990 14926 23042
rect 14978 22990 14980 23042
rect 14924 22482 14980 22990
rect 14924 22430 14926 22482
rect 14978 22430 14980 22482
rect 14924 22418 14980 22430
rect 14812 21812 14868 21822
rect 14700 21810 14868 21812
rect 14700 21758 14814 21810
rect 14866 21758 14868 21810
rect 14700 21756 14868 21758
rect 14812 21746 14868 21756
rect 14588 21698 14644 21710
rect 14588 21646 14590 21698
rect 14642 21646 14644 21698
rect 14140 21586 14308 21588
rect 14140 21534 14142 21586
rect 14194 21534 14308 21586
rect 14140 21532 14308 21534
rect 14364 21588 14420 21598
rect 14140 21522 14196 21532
rect 14028 21476 14084 21486
rect 14028 20690 14084 21420
rect 14140 20916 14196 20926
rect 14140 20822 14196 20860
rect 14028 20638 14030 20690
rect 14082 20638 14084 20690
rect 14028 20626 14084 20638
rect 14140 20690 14196 20702
rect 14140 20638 14142 20690
rect 14194 20638 14196 20690
rect 14140 19460 14196 20638
rect 14252 20692 14308 20702
rect 14364 20692 14420 21532
rect 14476 21588 14532 21598
rect 14588 21588 14644 21646
rect 14476 21586 14644 21588
rect 14476 21534 14478 21586
rect 14530 21534 14644 21586
rect 14476 21532 14644 21534
rect 14924 21586 14980 21598
rect 14924 21534 14926 21586
rect 14978 21534 14980 21586
rect 14476 21522 14532 21532
rect 14924 21476 14980 21534
rect 14924 21410 14980 21420
rect 15036 21588 15092 24446
rect 15148 23154 15204 23166
rect 15148 23102 15150 23154
rect 15202 23102 15204 23154
rect 15148 23044 15204 23102
rect 15148 22978 15204 22988
rect 15372 23154 15428 23166
rect 15932 23156 15988 23166
rect 15372 23102 15374 23154
rect 15426 23102 15428 23154
rect 15372 21812 15428 23102
rect 15820 23100 15932 23156
rect 15484 21812 15540 21822
rect 15372 21810 15540 21812
rect 15372 21758 15486 21810
rect 15538 21758 15540 21810
rect 15372 21756 15540 21758
rect 15484 21746 15540 21756
rect 15372 21588 15428 21598
rect 15036 21586 15652 21588
rect 15036 21534 15374 21586
rect 15426 21534 15652 21586
rect 15036 21532 15652 21534
rect 15036 21252 15092 21532
rect 15372 21522 15428 21532
rect 14476 21196 15092 21252
rect 14476 20802 14532 21196
rect 14476 20750 14478 20802
rect 14530 20750 14532 20802
rect 14476 20738 14532 20750
rect 14252 20690 14420 20692
rect 14252 20638 14254 20690
rect 14306 20638 14420 20690
rect 14252 20636 14420 20638
rect 14252 20626 14308 20636
rect 14252 20244 14308 20254
rect 14252 20150 14308 20188
rect 14140 19394 14196 19404
rect 15596 20132 15652 21532
rect 15708 21586 15764 21598
rect 15708 21534 15710 21586
rect 15762 21534 15764 21586
rect 15708 21476 15764 21534
rect 15708 21410 15764 21420
rect 15820 20580 15876 23100
rect 15932 23090 15988 23100
rect 16380 21812 16436 25452
rect 16604 25442 16660 25452
rect 16940 25506 16996 26124
rect 17500 25730 17556 26238
rect 18172 26180 18228 26190
rect 18172 26178 18340 26180
rect 18172 26126 18174 26178
rect 18226 26126 18340 26178
rect 18172 26124 18340 26126
rect 18172 26114 18228 26124
rect 17500 25678 17502 25730
rect 17554 25678 17556 25730
rect 17500 25666 17556 25678
rect 18060 25730 18116 25742
rect 18060 25678 18062 25730
rect 18114 25678 18116 25730
rect 16940 25454 16942 25506
rect 16994 25454 16996 25506
rect 16940 25442 16996 25454
rect 17164 25506 17220 25518
rect 17164 25454 17166 25506
rect 17218 25454 17220 25506
rect 16828 25396 16884 25406
rect 16828 25302 16884 25340
rect 17164 25396 17220 25454
rect 17164 25330 17220 25340
rect 17724 25396 17780 25406
rect 17724 25302 17780 25340
rect 16716 25284 16772 25294
rect 16716 25190 16772 25228
rect 18060 25282 18116 25678
rect 18284 25506 18340 26124
rect 18284 25454 18286 25506
rect 18338 25454 18340 25506
rect 18284 25442 18340 25454
rect 18620 25396 18676 25406
rect 19180 25396 19236 25406
rect 18620 25394 19236 25396
rect 18620 25342 18622 25394
rect 18674 25342 19182 25394
rect 19234 25342 19236 25394
rect 18620 25340 19236 25342
rect 18620 25330 18676 25340
rect 19180 25330 19236 25340
rect 18060 25230 18062 25282
rect 18114 25230 18116 25282
rect 18060 24612 18116 25230
rect 16604 23266 16660 23278
rect 16604 23214 16606 23266
rect 16658 23214 16660 23266
rect 16492 23156 16548 23166
rect 16492 23062 16548 23100
rect 16492 21812 16548 21822
rect 15932 21810 16548 21812
rect 15932 21758 16494 21810
rect 16546 21758 16548 21810
rect 15932 21756 16548 21758
rect 15932 21698 15988 21756
rect 16492 21746 16548 21756
rect 15932 21646 15934 21698
rect 15986 21646 15988 21698
rect 15932 21634 15988 21646
rect 16604 21476 16660 23214
rect 17948 23268 18004 23278
rect 17948 23174 18004 23212
rect 16828 23156 16884 23166
rect 16828 23062 16884 23100
rect 17836 23156 17892 23166
rect 17836 23062 17892 23100
rect 17500 23042 17556 23054
rect 17500 22990 17502 23042
rect 17554 22990 17556 23042
rect 17052 22482 17108 22494
rect 17052 22430 17054 22482
rect 17106 22430 17108 22482
rect 17052 21924 17108 22430
rect 17500 22484 17556 22990
rect 17500 22370 17556 22428
rect 18060 22484 18116 24556
rect 18508 25282 18564 25294
rect 18508 25230 18510 25282
rect 18562 25230 18564 25282
rect 18060 22418 18116 22428
rect 18172 23154 18228 23166
rect 18172 23102 18174 23154
rect 18226 23102 18228 23154
rect 18172 22482 18228 23102
rect 18172 22430 18174 22482
rect 18226 22430 18228 22482
rect 18172 22418 18228 22430
rect 17500 22318 17502 22370
rect 17554 22318 17556 22370
rect 17500 22306 17556 22318
rect 18508 22372 18564 25230
rect 19292 23268 19348 26852
rect 19404 26180 19460 37996
rect 19740 37986 19796 37996
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20188 37492 20244 41200
rect 22204 38162 22260 41200
rect 24892 38276 24948 41200
rect 25564 39172 25620 41200
rect 25564 39116 25844 39172
rect 24892 38210 24948 38220
rect 22204 38110 22206 38162
rect 22258 38110 22260 38162
rect 22204 38098 22260 38110
rect 23772 38050 23828 38062
rect 23772 37998 23774 38050
rect 23826 37998 23828 38050
rect 20188 37426 20244 37436
rect 21420 37492 21476 37502
rect 21420 37398 21476 37436
rect 20412 37266 20468 37278
rect 20412 37214 20414 37266
rect 20466 37214 20468 37266
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19516 28084 19572 28094
rect 20412 28084 20468 37214
rect 22764 28642 22820 28654
rect 22764 28590 22766 28642
rect 22818 28590 22820 28642
rect 22428 28420 22484 28430
rect 22764 28420 22820 28590
rect 22428 28418 22820 28420
rect 22428 28366 22430 28418
rect 22482 28366 22820 28418
rect 22428 28364 22820 28366
rect 22428 28354 22484 28364
rect 19516 27990 19572 28028
rect 20188 28028 20412 28084
rect 19628 27858 19684 27870
rect 19628 27806 19630 27858
rect 19682 27806 19684 27858
rect 19628 26908 19684 27806
rect 20076 27858 20132 27870
rect 20076 27806 20078 27858
rect 20130 27806 20132 27858
rect 20076 26964 20132 27806
rect 20188 27186 20244 28028
rect 20412 28018 20468 28028
rect 22428 27860 22484 27870
rect 22316 27804 22428 27860
rect 20748 27748 20804 27758
rect 21980 27748 22036 27758
rect 20748 27746 21252 27748
rect 20748 27694 20750 27746
rect 20802 27694 21252 27746
rect 20748 27692 21252 27694
rect 20748 27682 20804 27692
rect 20188 27134 20190 27186
rect 20242 27134 20244 27186
rect 20188 27122 20244 27134
rect 20636 27076 20692 27086
rect 20300 27020 20636 27076
rect 20692 27020 20804 27076
rect 20300 26964 20356 27020
rect 20636 26982 20692 27020
rect 20076 26908 20356 26964
rect 19404 25394 19460 26124
rect 19516 26852 19684 26908
rect 20188 26852 20580 26908
rect 19516 25508 19572 26852
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20300 26180 20356 26190
rect 20300 26086 20356 26124
rect 19516 25414 19572 25452
rect 19404 25342 19406 25394
rect 19458 25342 19460 25394
rect 19404 25330 19460 25342
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20524 23940 20580 26852
rect 20748 26514 20804 27020
rect 21196 27074 21252 27692
rect 21196 27022 21198 27074
rect 21250 27022 21252 27074
rect 21196 27010 21252 27022
rect 20748 26462 20750 26514
rect 20802 26462 20804 26514
rect 20748 26450 20804 26462
rect 21420 26962 21476 26974
rect 21420 26910 21422 26962
rect 21474 26910 21476 26962
rect 21420 26180 21476 26910
rect 21532 26964 21588 26974
rect 21756 26964 21812 26974
rect 21532 26962 21812 26964
rect 21532 26910 21534 26962
rect 21586 26910 21758 26962
rect 21810 26910 21812 26962
rect 21532 26908 21812 26910
rect 21532 26898 21588 26908
rect 21756 26898 21812 26908
rect 21980 26962 22036 27692
rect 21980 26910 21982 26962
rect 22034 26910 22036 26962
rect 21980 26898 22036 26910
rect 22092 26962 22148 26974
rect 22092 26910 22094 26962
rect 22146 26910 22148 26962
rect 22092 26516 22148 26910
rect 21420 26114 21476 26124
rect 21980 26460 22148 26516
rect 21980 26292 22036 26460
rect 22204 26404 22260 26414
rect 22204 26310 22260 26348
rect 21644 25508 21700 25518
rect 21980 25508 22036 26236
rect 21700 25452 22036 25508
rect 22092 26290 22148 26302
rect 22092 26238 22094 26290
rect 22146 26238 22148 26290
rect 22092 26180 22148 26238
rect 21644 25394 21700 25452
rect 21644 25342 21646 25394
rect 21698 25342 21700 25394
rect 21644 25330 21700 25342
rect 21980 25282 22036 25294
rect 21980 25230 21982 25282
rect 22034 25230 22036 25282
rect 21868 24724 21924 24734
rect 21980 24724 22036 25230
rect 21868 24722 22036 24724
rect 21868 24670 21870 24722
rect 21922 24670 22036 24722
rect 21868 24668 22036 24670
rect 21868 24658 21924 24668
rect 20524 23846 20580 23884
rect 21532 23940 21588 23950
rect 21868 23940 21924 23950
rect 21588 23938 21924 23940
rect 21588 23886 21870 23938
rect 21922 23886 21924 23938
rect 21588 23884 21924 23886
rect 21532 23846 21588 23884
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19292 23202 19348 23212
rect 20188 23268 20244 23278
rect 18508 22306 18564 22316
rect 19836 21980 20100 21990
rect 17052 21858 17108 21868
rect 18172 21924 18228 21934
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 17388 21698 17444 21710
rect 17388 21646 17390 21698
rect 17442 21646 17444 21698
rect 16604 21410 16660 21420
rect 16716 21586 16772 21598
rect 16716 21534 16718 21586
rect 16770 21534 16772 21586
rect 15820 20524 16212 20580
rect 15708 20132 15764 20142
rect 15596 20130 15764 20132
rect 15596 20078 15710 20130
rect 15762 20078 15764 20130
rect 15596 20076 15764 20078
rect 13692 19122 13748 19134
rect 13692 19070 13694 19122
rect 13746 19070 13748 19122
rect 13692 19012 13748 19070
rect 13580 18564 13636 18574
rect 13468 18562 13636 18564
rect 13468 18510 13582 18562
rect 13634 18510 13636 18562
rect 13468 18508 13636 18510
rect 13580 18498 13636 18508
rect 13580 17780 13636 17790
rect 13020 17778 13636 17780
rect 13020 17726 13582 17778
rect 13634 17726 13636 17778
rect 13020 17724 13636 17726
rect 13580 17714 13636 17724
rect 13468 17556 13524 17566
rect 13692 17556 13748 18956
rect 13804 17892 13860 17902
rect 13804 17666 13860 17836
rect 13804 17614 13806 17666
rect 13858 17614 13860 17666
rect 13804 17602 13860 17614
rect 13916 17668 13972 19180
rect 14252 19236 14308 19246
rect 14252 19234 14868 19236
rect 14252 19182 14254 19234
rect 14306 19182 14868 19234
rect 14252 19180 14868 19182
rect 14252 19170 14308 19180
rect 14700 19012 14756 19022
rect 14588 19010 14756 19012
rect 14588 18958 14702 19010
rect 14754 18958 14756 19010
rect 14588 18956 14756 18958
rect 14364 18452 14420 18462
rect 14588 18452 14644 18956
rect 14700 18946 14756 18956
rect 14700 18676 14756 18686
rect 14700 18582 14756 18620
rect 14812 18674 14868 19180
rect 15372 19124 15428 19134
rect 15372 19030 15428 19068
rect 14812 18622 14814 18674
rect 14866 18622 14868 18674
rect 14812 18610 14868 18622
rect 15596 18676 15652 20076
rect 15708 20066 15764 20076
rect 16044 20020 16100 20030
rect 16044 19926 16100 19964
rect 16044 19460 16100 19470
rect 15708 19012 15764 19022
rect 15708 19010 15876 19012
rect 15708 18958 15710 19010
rect 15762 18958 15876 19010
rect 15708 18956 15876 18958
rect 15708 18946 15764 18956
rect 15596 18610 15652 18620
rect 14924 18564 14980 18574
rect 14924 18470 14980 18508
rect 15820 18564 15876 18956
rect 16044 18676 16100 19404
rect 16156 19124 16212 20524
rect 16492 19236 16548 19246
rect 16716 19236 16772 21534
rect 17388 21476 17444 21646
rect 18172 21698 18228 21868
rect 18172 21646 18174 21698
rect 18226 21646 18228 21698
rect 18172 21634 18228 21646
rect 17388 21410 17444 21420
rect 17724 21586 17780 21598
rect 17724 21534 17726 21586
rect 17778 21534 17780 21586
rect 17724 21476 17780 21534
rect 19068 21588 19124 21598
rect 19404 21588 19460 21598
rect 19068 21494 19124 21532
rect 19180 21586 19460 21588
rect 19180 21534 19406 21586
rect 19458 21534 19460 21586
rect 19180 21532 19460 21534
rect 17724 21410 17780 21420
rect 18620 21476 18676 21486
rect 18060 21362 18116 21374
rect 18060 21310 18062 21362
rect 18114 21310 18116 21362
rect 16492 19234 16772 19236
rect 16492 19182 16494 19234
rect 16546 19182 16772 19234
rect 16492 19180 16772 19182
rect 16492 19170 16548 19180
rect 16156 19030 16212 19068
rect 16044 18620 16212 18676
rect 15820 18470 15876 18508
rect 14364 18450 14644 18452
rect 14364 18398 14366 18450
rect 14418 18398 14644 18450
rect 14364 18396 14644 18398
rect 14700 18452 14756 18462
rect 14028 18004 14084 18014
rect 14028 17890 14084 17948
rect 14028 17838 14030 17890
rect 14082 17838 14084 17890
rect 14028 17826 14084 17838
rect 14028 17668 14084 17678
rect 13916 17666 14084 17668
rect 13916 17614 14030 17666
rect 14082 17614 14084 17666
rect 13916 17612 14084 17614
rect 14028 17602 14084 17612
rect 13468 17554 13748 17556
rect 13468 17502 13470 17554
rect 13522 17502 13748 17554
rect 13468 17500 13748 17502
rect 13468 17490 13524 17500
rect 14028 16884 14084 16894
rect 14364 16884 14420 18396
rect 14476 18004 14532 18014
rect 14476 17892 14532 17948
rect 14588 17892 14644 17902
rect 14476 17890 14644 17892
rect 14476 17838 14590 17890
rect 14642 17838 14644 17890
rect 14476 17836 14644 17838
rect 14588 17826 14644 17836
rect 14700 17554 14756 18396
rect 15372 18450 15428 18462
rect 15372 18398 15374 18450
rect 15426 18398 15428 18450
rect 14924 17892 14980 17902
rect 14924 17798 14980 17836
rect 15372 17668 15428 18398
rect 15372 17602 15428 17612
rect 16044 18450 16100 18462
rect 16044 18398 16046 18450
rect 16098 18398 16100 18450
rect 14700 17502 14702 17554
rect 14754 17502 14756 17554
rect 14700 17490 14756 17502
rect 14700 17108 14756 17118
rect 14700 16994 14756 17052
rect 16044 17108 16100 18398
rect 16156 18450 16212 18620
rect 16156 18398 16158 18450
rect 16210 18398 16212 18450
rect 16156 18386 16212 18398
rect 16268 18452 16324 18462
rect 16268 18358 16324 18396
rect 16716 18340 16772 19180
rect 17500 20916 17556 20926
rect 16716 18274 16772 18284
rect 17164 18564 17220 18574
rect 16716 17668 16772 17678
rect 16716 17574 16772 17612
rect 17164 17666 17220 18508
rect 17164 17614 17166 17666
rect 17218 17614 17220 17666
rect 17164 17602 17220 17614
rect 17388 18452 17444 18462
rect 16044 17042 16100 17052
rect 17276 17554 17332 17566
rect 17276 17502 17278 17554
rect 17330 17502 17332 17554
rect 14700 16942 14702 16994
rect 14754 16942 14756 16994
rect 14700 16930 14756 16942
rect 14028 16882 14420 16884
rect 14028 16830 14030 16882
rect 14082 16830 14420 16882
rect 14028 16828 14420 16830
rect 17276 16884 17332 17502
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 14028 13972 14084 16828
rect 17276 16818 17332 16828
rect 17388 17556 17444 18396
rect 16828 16772 16884 16782
rect 16828 16678 16884 16716
rect 17388 16770 17444 17500
rect 17388 16718 17390 16770
rect 17442 16718 17444 16770
rect 17388 16706 17444 16718
rect 17500 16770 17556 20860
rect 18060 20244 18116 21310
rect 18060 20150 18116 20188
rect 18620 20692 18676 21420
rect 17724 20132 17780 20142
rect 17724 20038 17780 20076
rect 18396 20130 18452 20142
rect 18396 20078 18398 20130
rect 18450 20078 18452 20130
rect 18396 20020 18452 20078
rect 18396 19954 18452 19964
rect 18508 20132 18564 20142
rect 18508 18564 18564 20076
rect 18620 18674 18676 20636
rect 19180 20914 19236 21532
rect 19404 21522 19460 21532
rect 19180 20862 19182 20914
rect 19234 20862 19236 20914
rect 19180 20580 19236 20862
rect 20076 20804 20132 20814
rect 20076 20710 20132 20748
rect 19740 20580 19796 20590
rect 19180 20514 19236 20524
rect 19516 20578 19796 20580
rect 19516 20526 19742 20578
rect 19794 20526 19796 20578
rect 19516 20524 19796 20526
rect 18732 20132 18788 20142
rect 18732 20038 18788 20076
rect 18620 18622 18622 18674
rect 18674 18622 18676 18674
rect 18620 18610 18676 18622
rect 19516 18676 19572 20524
rect 19740 20514 19796 20524
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 18508 18470 18564 18508
rect 18172 18452 18228 18462
rect 18172 17554 18228 18396
rect 19292 18340 19348 18350
rect 19292 18246 19348 18284
rect 18620 18226 18676 18238
rect 18620 18174 18622 18226
rect 18674 18174 18676 18226
rect 18172 17502 18174 17554
rect 18226 17502 18228 17554
rect 18172 17490 18228 17502
rect 18508 17668 18564 17678
rect 17836 17442 17892 17454
rect 17836 17390 17838 17442
rect 17890 17390 17892 17442
rect 17724 17108 17780 17118
rect 17724 16882 17780 17052
rect 17724 16830 17726 16882
rect 17778 16830 17780 16882
rect 17724 16818 17780 16830
rect 17500 16718 17502 16770
rect 17554 16718 17556 16770
rect 17052 15874 17108 15886
rect 17052 15822 17054 15874
rect 17106 15822 17108 15874
rect 16492 14532 16548 14542
rect 16492 14438 16548 14476
rect 14028 13746 14084 13916
rect 14700 14308 14756 14318
rect 14700 13858 14756 14252
rect 16380 14308 16436 14318
rect 16380 14214 16436 14252
rect 14700 13806 14702 13858
rect 14754 13806 14756 13858
rect 14700 13794 14756 13806
rect 16940 13972 16996 13982
rect 17052 13972 17108 15822
rect 17164 14756 17220 14766
rect 17164 14530 17220 14700
rect 17164 14478 17166 14530
rect 17218 14478 17220 14530
rect 17164 14466 17220 14478
rect 17276 14642 17332 14654
rect 17276 14590 17278 14642
rect 17330 14590 17332 14642
rect 17276 14532 17332 14590
rect 17500 14532 17556 16718
rect 17836 16772 17892 17390
rect 18508 17106 18564 17612
rect 18508 17054 18510 17106
rect 18562 17054 18564 17106
rect 18508 17042 18564 17054
rect 17836 16706 17892 16716
rect 17948 16884 18004 16894
rect 17948 15148 18004 16828
rect 18396 16882 18452 16894
rect 18396 16830 18398 16882
rect 18450 16830 18452 16882
rect 18284 16772 18340 16782
rect 18396 16772 18452 16830
rect 18340 16716 18452 16772
rect 18284 16706 18340 16716
rect 18620 16100 18676 18174
rect 19516 17892 19572 18620
rect 19628 20132 19684 20142
rect 19628 18564 19684 20076
rect 20188 20020 20244 23212
rect 21756 23042 21812 23884
rect 21868 23874 21924 23884
rect 21980 23716 22036 24668
rect 21756 22990 21758 23042
rect 21810 22990 21812 23042
rect 20300 22482 20356 22494
rect 20300 22430 20302 22482
rect 20354 22430 20356 22482
rect 20300 22372 20356 22430
rect 21756 22484 21812 22990
rect 21756 22418 21812 22428
rect 21868 23660 22036 23716
rect 21868 23492 21924 23660
rect 21532 22372 21588 22382
rect 20300 22316 20804 22372
rect 20748 22260 20804 22316
rect 21084 22370 21588 22372
rect 21084 22318 21534 22370
rect 21586 22318 21588 22370
rect 21084 22316 21588 22318
rect 20748 22258 20916 22260
rect 20748 22206 20750 22258
rect 20802 22206 20916 22258
rect 20748 22204 20916 22206
rect 20748 22194 20804 22204
rect 20636 22146 20692 22158
rect 20636 22094 20638 22146
rect 20690 22094 20692 22146
rect 20636 20804 20692 22094
rect 20748 22036 20804 22046
rect 20748 21026 20804 21980
rect 20748 20974 20750 21026
rect 20802 20974 20804 21026
rect 20748 20962 20804 20974
rect 20860 21588 20916 22204
rect 20412 20692 20468 20702
rect 20300 20690 20468 20692
rect 20300 20638 20414 20690
rect 20466 20638 20468 20690
rect 20300 20636 20468 20638
rect 20300 20244 20356 20636
rect 20412 20626 20468 20636
rect 20636 20690 20692 20748
rect 20636 20638 20638 20690
rect 20690 20638 20692 20690
rect 20636 20626 20692 20638
rect 20636 20356 20692 20366
rect 20300 20178 20356 20188
rect 20524 20244 20580 20254
rect 20412 20132 20468 20142
rect 20412 20038 20468 20076
rect 20188 19964 20356 20020
rect 20188 19796 20244 19806
rect 20188 19702 20244 19740
rect 20300 19346 20356 19964
rect 20524 19906 20580 20188
rect 20524 19854 20526 19906
rect 20578 19854 20580 19906
rect 20524 19842 20580 19854
rect 20300 19294 20302 19346
rect 20354 19294 20356 19346
rect 20300 19282 20356 19294
rect 20412 19796 20468 19806
rect 20076 19012 20132 19050
rect 20300 19012 20356 19022
rect 20076 18946 20132 18956
rect 20188 19010 20356 19012
rect 20188 18958 20302 19010
rect 20354 18958 20356 19010
rect 20188 18956 20356 18958
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 18470 19684 18508
rect 19516 17826 19572 17836
rect 19964 18450 20020 18462
rect 19964 18398 19966 18450
rect 20018 18398 20020 18450
rect 19964 18340 20020 18398
rect 19292 17556 19348 17566
rect 19292 17462 19348 17500
rect 18844 17442 18900 17454
rect 18844 17390 18846 17442
rect 18898 17390 18900 17442
rect 18844 17108 18900 17390
rect 18844 17042 18900 17052
rect 19628 17444 19684 17454
rect 19964 17444 20020 18284
rect 20188 17556 20244 18956
rect 20300 18946 20356 18956
rect 20300 18564 20356 18574
rect 20300 18450 20356 18508
rect 20300 18398 20302 18450
rect 20354 18398 20356 18450
rect 20300 18386 20356 18398
rect 20412 17556 20468 19740
rect 20636 19234 20692 20300
rect 20860 20130 20916 21532
rect 20860 20078 20862 20130
rect 20914 20078 20916 20130
rect 20860 20066 20916 20078
rect 20636 19182 20638 19234
rect 20690 19182 20692 19234
rect 20524 18340 20580 18350
rect 20524 18246 20580 18284
rect 20188 17490 20244 17500
rect 20300 17554 20468 17556
rect 20300 17502 20414 17554
rect 20466 17502 20468 17554
rect 20300 17500 20468 17502
rect 20076 17444 20132 17454
rect 19628 17442 20132 17444
rect 19628 17390 19630 17442
rect 19682 17390 20078 17442
rect 20130 17390 20132 17442
rect 19628 17388 20132 17390
rect 18620 16034 18676 16044
rect 18732 15876 18788 15886
rect 17724 15092 18004 15148
rect 18060 15202 18116 15214
rect 18060 15150 18062 15202
rect 18114 15150 18116 15202
rect 17612 14532 17668 14542
rect 17500 14476 17612 14532
rect 17276 14466 17332 14476
rect 17612 14438 17668 14476
rect 17724 14530 17780 15092
rect 18060 14756 18116 15150
rect 18060 14690 18116 14700
rect 18732 14642 18788 15820
rect 18732 14590 18734 14642
rect 18786 14590 18788 14642
rect 18732 14578 18788 14590
rect 17724 14478 17726 14530
rect 17778 14478 17780 14530
rect 17724 14466 17780 14478
rect 18508 14532 18564 14542
rect 18508 14438 18564 14476
rect 16996 13916 17108 13972
rect 17388 14306 17444 14318
rect 17388 14254 17390 14306
rect 17442 14254 17444 14306
rect 14028 13694 14030 13746
rect 14082 13694 14084 13746
rect 14028 13682 14084 13694
rect 16828 13634 16884 13646
rect 16828 13582 16830 13634
rect 16882 13582 16884 13634
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 16828 12740 16884 13582
rect 16940 12962 16996 13916
rect 16940 12910 16942 12962
rect 16994 12910 16996 12962
rect 16940 12898 16996 12910
rect 17388 12740 17444 14254
rect 18172 14306 18228 14318
rect 18172 14254 18174 14306
rect 18226 14254 18228 14306
rect 17500 13972 17556 13982
rect 17500 13878 17556 13916
rect 17836 13860 17892 13870
rect 17612 13858 17892 13860
rect 17612 13806 17838 13858
rect 17890 13806 17892 13858
rect 17612 13804 17892 13806
rect 17612 13074 17668 13804
rect 17836 13794 17892 13804
rect 18172 13858 18228 14254
rect 18172 13806 18174 13858
rect 18226 13806 18228 13858
rect 18172 13794 18228 13806
rect 17612 13022 17614 13074
rect 17666 13022 17668 13074
rect 17612 13010 17668 13022
rect 19628 13076 19684 17388
rect 20076 17378 20132 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20076 17108 20132 17118
rect 19852 16100 19908 16110
rect 19852 16006 19908 16044
rect 20076 16098 20132 17052
rect 20300 17106 20356 17500
rect 20412 17490 20468 17500
rect 20300 17054 20302 17106
rect 20354 17054 20356 17106
rect 20300 17042 20356 17054
rect 20412 16884 20468 16894
rect 20636 16884 20692 19182
rect 20748 18452 20804 18462
rect 21084 18452 21140 22316
rect 21532 22306 21588 22316
rect 21644 22372 21700 22382
rect 21308 22148 21364 22158
rect 21644 22148 21700 22316
rect 21308 22146 21700 22148
rect 21308 22094 21310 22146
rect 21362 22094 21700 22146
rect 21308 22092 21700 22094
rect 21308 22082 21364 22092
rect 21756 22036 21812 22046
rect 21868 22036 21924 23436
rect 21812 21980 21924 22036
rect 21980 22148 22036 22158
rect 21756 21970 21812 21980
rect 21532 21588 21588 21598
rect 21420 20802 21476 20814
rect 21420 20750 21422 20802
rect 21474 20750 21476 20802
rect 21420 20692 21476 20750
rect 21196 20132 21252 20142
rect 21196 20038 21252 20076
rect 21420 19122 21476 20636
rect 21532 20356 21588 21532
rect 21980 21140 22036 22092
rect 21532 19906 21588 20300
rect 21756 21084 22036 21140
rect 21532 19854 21534 19906
rect 21586 19854 21588 19906
rect 21532 19842 21588 19854
rect 21644 20132 21700 20142
rect 21420 19070 21422 19122
rect 21474 19070 21476 19122
rect 21420 19058 21476 19070
rect 21532 19234 21588 19246
rect 21532 19182 21534 19234
rect 21586 19182 21588 19234
rect 21420 18564 21476 18574
rect 21420 18470 21476 18508
rect 21196 18452 21252 18462
rect 21084 18450 21364 18452
rect 21084 18398 21198 18450
rect 21250 18398 21364 18450
rect 21084 18396 21364 18398
rect 20748 18358 20804 18396
rect 21196 18386 21252 18396
rect 21196 18228 21252 18238
rect 21196 17780 21252 18172
rect 21084 17556 21140 17566
rect 21084 17106 21140 17500
rect 21084 17054 21086 17106
rect 21138 17054 21140 17106
rect 21084 17042 21140 17054
rect 20412 16882 20692 16884
rect 20412 16830 20414 16882
rect 20466 16830 20692 16882
rect 20412 16828 20692 16830
rect 20860 16994 20916 17006
rect 20860 16942 20862 16994
rect 20914 16942 20916 16994
rect 20412 16818 20468 16828
rect 20860 16772 20916 16942
rect 21196 16996 21252 17724
rect 21308 17108 21364 18396
rect 21532 17668 21588 19182
rect 21644 18452 21700 20076
rect 21756 20020 21812 21084
rect 21868 20914 21924 20926
rect 21868 20862 21870 20914
rect 21922 20862 21924 20914
rect 21868 20244 21924 20862
rect 21868 20178 21924 20188
rect 21868 20020 21924 20030
rect 21756 20018 21924 20020
rect 21756 19966 21870 20018
rect 21922 19966 21924 20018
rect 21756 19964 21924 19966
rect 21868 19954 21924 19964
rect 22092 19458 22148 26124
rect 22316 25732 22372 27804
rect 22428 27794 22484 27804
rect 22652 27076 22708 27086
rect 22764 27076 22820 28364
rect 22876 28532 22932 28542
rect 23548 28532 23604 28542
rect 22876 27748 22932 28476
rect 23436 28530 23604 28532
rect 23436 28478 23550 28530
rect 23602 28478 23604 28530
rect 23436 28476 23604 28478
rect 23436 27972 23492 28476
rect 23548 28466 23604 28476
rect 23772 28532 23828 37998
rect 25564 38052 25620 38062
rect 25564 38050 25732 38052
rect 25564 37998 25566 38050
rect 25618 37998 25732 38050
rect 25564 37996 25732 37998
rect 25564 37986 25620 37996
rect 25676 28756 25732 37996
rect 25788 37492 25844 39116
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 26124 38276 26180 38286
rect 26124 38182 26180 38220
rect 25788 37426 25844 37436
rect 26796 37492 26852 37502
rect 26796 37398 26852 37436
rect 23772 28466 23828 28476
rect 25340 28754 25732 28756
rect 25340 28702 25678 28754
rect 25730 28702 25732 28754
rect 25340 28700 25732 28702
rect 25340 28082 25396 28700
rect 25676 28690 25732 28700
rect 25900 37266 25956 37278
rect 25900 37214 25902 37266
rect 25954 37214 25956 37266
rect 25340 28030 25342 28082
rect 25394 28030 25396 28082
rect 25340 28018 25396 28030
rect 23436 27906 23492 27916
rect 23324 27858 23380 27870
rect 23324 27806 23326 27858
rect 23378 27806 23380 27858
rect 22876 27654 22932 27692
rect 23100 27748 23156 27758
rect 23100 27076 23156 27692
rect 22708 27074 23156 27076
rect 22708 27022 23102 27074
rect 23154 27022 23156 27074
rect 22708 27020 23156 27022
rect 22652 26982 22708 27020
rect 23100 27010 23156 27020
rect 23324 26740 23380 27806
rect 23548 27860 23604 27870
rect 23548 27766 23604 27804
rect 23996 27858 24052 27870
rect 23996 27806 23998 27858
rect 24050 27806 24052 27858
rect 23436 27746 23492 27758
rect 23436 27694 23438 27746
rect 23490 27694 23492 27746
rect 23436 27636 23492 27694
rect 23436 27580 23828 27636
rect 23772 27186 23828 27580
rect 23772 27134 23774 27186
rect 23826 27134 23828 27186
rect 23772 27122 23828 27134
rect 22988 26684 23380 26740
rect 23772 26964 23828 26974
rect 22428 26516 22484 26526
rect 22988 26516 23044 26684
rect 23100 26516 23156 26526
rect 22428 26514 23156 26516
rect 22428 26462 22430 26514
rect 22482 26462 23102 26514
rect 23154 26462 23156 26514
rect 22428 26460 23156 26462
rect 22428 26450 22484 26460
rect 23100 26450 23156 26460
rect 23436 26404 23492 26414
rect 23492 26348 23604 26404
rect 23436 26338 23492 26348
rect 23324 26292 23380 26302
rect 23324 26198 23380 26236
rect 23212 26180 23268 26190
rect 23212 26086 23268 26124
rect 22428 25732 22484 25742
rect 22316 25730 22484 25732
rect 22316 25678 22430 25730
rect 22482 25678 22484 25730
rect 22316 25676 22484 25678
rect 22428 25666 22484 25676
rect 22316 25396 22372 25406
rect 22204 25394 22372 25396
rect 22204 25342 22318 25394
rect 22370 25342 22372 25394
rect 22204 25340 22372 25342
rect 22204 25284 22260 25340
rect 22316 25330 22372 25340
rect 22428 25396 22484 25406
rect 22204 21026 22260 25228
rect 22316 24612 22372 24622
rect 22428 24612 22484 25340
rect 23324 24724 23380 24734
rect 22372 24556 22484 24612
rect 23212 24722 23380 24724
rect 23212 24670 23326 24722
rect 23378 24670 23380 24722
rect 23212 24668 23380 24670
rect 22316 24518 22372 24556
rect 22652 23826 22708 23838
rect 22652 23774 22654 23826
rect 22706 23774 22708 23826
rect 22652 22484 22708 23774
rect 23212 23492 23268 24668
rect 23324 24658 23380 24668
rect 23212 23426 23268 23436
rect 23324 24500 23380 24510
rect 22988 23154 23044 23166
rect 22988 23102 22990 23154
rect 23042 23102 23044 23154
rect 22764 22484 22820 22494
rect 22652 22482 22820 22484
rect 22652 22430 22766 22482
rect 22818 22430 22820 22482
rect 22652 22428 22820 22430
rect 22764 22418 22820 22428
rect 22428 22372 22484 22382
rect 22484 22316 22708 22372
rect 22428 22306 22484 22316
rect 22652 22258 22708 22316
rect 22652 22206 22654 22258
rect 22706 22206 22708 22258
rect 22652 22194 22708 22206
rect 22316 22146 22372 22158
rect 22876 22148 22932 22158
rect 22316 22094 22318 22146
rect 22370 22094 22372 22146
rect 22316 22036 22372 22094
rect 22764 22146 22932 22148
rect 22764 22094 22878 22146
rect 22930 22094 22932 22146
rect 22764 22092 22932 22094
rect 22764 22036 22820 22092
rect 22876 22082 22932 22092
rect 22316 21980 22820 22036
rect 22204 20974 22206 21026
rect 22258 20974 22260 21026
rect 22204 20962 22260 20974
rect 22316 20802 22372 20814
rect 22316 20750 22318 20802
rect 22370 20750 22372 20802
rect 22316 20692 22372 20750
rect 22540 20692 22596 20702
rect 22316 20636 22540 20692
rect 22092 19406 22094 19458
rect 22146 19406 22148 19458
rect 22092 19394 22148 19406
rect 22204 19906 22260 19918
rect 22204 19854 22206 19906
rect 22258 19854 22260 19906
rect 22204 19796 22260 19854
rect 22204 19234 22260 19740
rect 22204 19182 22206 19234
rect 22258 19182 22260 19234
rect 22204 19170 22260 19182
rect 22316 19794 22372 19806
rect 22316 19742 22318 19794
rect 22370 19742 22372 19794
rect 21868 19012 21924 19022
rect 21756 18676 21812 18686
rect 21868 18676 21924 18956
rect 22204 18788 22260 18798
rect 22316 18788 22372 19742
rect 22260 18732 22372 18788
rect 22428 18788 22484 20636
rect 22540 20626 22596 20636
rect 22652 20580 22708 20590
rect 22764 20580 22820 21980
rect 22988 21700 23044 23102
rect 23324 22370 23380 24444
rect 23548 23492 23604 26348
rect 23772 26290 23828 26908
rect 23996 26516 24052 27806
rect 25116 27858 25172 27870
rect 25116 27806 25118 27858
rect 25170 27806 25172 27858
rect 24332 27748 24388 27758
rect 24332 27654 24388 27692
rect 25116 26964 25172 27806
rect 25452 27858 25508 27870
rect 25452 27806 25454 27858
rect 25506 27806 25508 27858
rect 25452 27300 25508 27806
rect 25116 26898 25172 26908
rect 25228 27244 25508 27300
rect 23996 26450 24052 26460
rect 25116 26516 25172 26526
rect 25116 26422 25172 26460
rect 23772 26238 23774 26290
rect 23826 26238 23828 26290
rect 23772 26226 23828 26238
rect 25228 26292 25284 27244
rect 25900 27188 25956 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 25340 27186 25956 27188
rect 25340 27134 25902 27186
rect 25954 27134 25956 27186
rect 25340 27132 25956 27134
rect 25340 26514 25396 27132
rect 25900 27122 25956 27132
rect 25340 26462 25342 26514
rect 25394 26462 25396 26514
rect 25340 26450 25396 26462
rect 25452 26292 25508 26302
rect 25228 26290 25620 26292
rect 25228 26238 25454 26290
rect 25506 26238 25620 26290
rect 25228 26236 25620 26238
rect 25452 26226 25508 26236
rect 23660 24836 23716 24846
rect 23660 24742 23716 24780
rect 24108 24834 24164 24846
rect 24108 24782 24110 24834
rect 24162 24782 24164 24834
rect 24108 24724 24164 24782
rect 25564 24836 25620 26236
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 24108 24658 24164 24668
rect 24220 24722 24276 24734
rect 24220 24670 24222 24722
rect 24274 24670 24276 24722
rect 24220 24612 24276 24670
rect 24780 24724 24836 24734
rect 24668 24612 24724 24622
rect 24276 24610 24724 24612
rect 24276 24558 24670 24610
rect 24722 24558 24724 24610
rect 24276 24556 24724 24558
rect 24220 24518 24276 24556
rect 24108 24500 24164 24510
rect 24108 24406 24164 24444
rect 23548 23436 23716 23492
rect 23324 22318 23326 22370
rect 23378 22318 23380 22370
rect 23324 22306 23380 22318
rect 23548 22372 23604 22382
rect 23548 22278 23604 22316
rect 23660 22258 23716 23436
rect 24668 23268 24724 24556
rect 24780 24050 24836 24668
rect 24780 23998 24782 24050
rect 24834 23998 24836 24050
rect 24780 23986 24836 23998
rect 25452 23938 25508 23950
rect 25452 23886 25454 23938
rect 25506 23886 25508 23938
rect 24668 23212 24836 23268
rect 23884 23156 23940 23166
rect 23884 22370 23940 23100
rect 24332 22484 24388 22494
rect 24332 22390 24388 22428
rect 24668 22372 24724 22382
rect 23884 22318 23886 22370
rect 23938 22318 23940 22370
rect 23884 22306 23940 22318
rect 24444 22370 24724 22372
rect 24444 22318 24670 22370
rect 24722 22318 24724 22370
rect 24444 22316 24724 22318
rect 23660 22206 23662 22258
rect 23714 22206 23716 22258
rect 23660 22194 23716 22206
rect 22708 20524 22820 20580
rect 22876 21698 23044 21700
rect 22876 21646 22990 21698
rect 23042 21646 23044 21698
rect 22876 21644 23044 21646
rect 22540 20020 22596 20030
rect 22540 19234 22596 19964
rect 22540 19182 22542 19234
rect 22594 19182 22596 19234
rect 22540 19170 22596 19182
rect 22428 18732 22596 18788
rect 21980 18676 22036 18686
rect 21756 18674 21980 18676
rect 21756 18622 21758 18674
rect 21810 18622 21980 18674
rect 21756 18620 21980 18622
rect 21756 18610 21812 18620
rect 21980 18610 22036 18620
rect 21644 18386 21700 18396
rect 22092 18452 22148 18462
rect 22092 18358 22148 18396
rect 21588 17612 22036 17668
rect 21532 17574 21588 17612
rect 21308 17052 21476 17108
rect 21196 16940 21364 16996
rect 21308 16882 21364 16940
rect 21308 16830 21310 16882
rect 21362 16830 21364 16882
rect 21308 16818 21364 16830
rect 20524 16716 20860 16772
rect 20076 16046 20078 16098
rect 20130 16046 20132 16098
rect 20076 16034 20132 16046
rect 20300 16658 20356 16670
rect 20300 16606 20302 16658
rect 20354 16606 20356 16658
rect 20300 15988 20356 16606
rect 20300 15894 20356 15932
rect 19964 15876 20020 15886
rect 19964 15874 20244 15876
rect 19964 15822 19966 15874
rect 20018 15822 20244 15874
rect 19964 15820 20244 15822
rect 19964 15810 20020 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20188 14980 20244 15820
rect 20524 15314 20580 16716
rect 20860 16706 20916 16716
rect 21196 16770 21252 16782
rect 21196 16718 21198 16770
rect 21250 16718 21252 16770
rect 20524 15262 20526 15314
rect 20578 15262 20580 15314
rect 20524 15250 20580 15262
rect 20748 16212 20804 16222
rect 20748 15314 20804 16156
rect 20748 15262 20750 15314
rect 20802 15262 20804 15314
rect 20748 15250 20804 15262
rect 21196 15148 21252 16718
rect 21420 16212 21476 17052
rect 21980 17106 22036 17612
rect 21980 17054 21982 17106
rect 22034 17054 22036 17106
rect 21980 17042 22036 17054
rect 22092 16996 22148 17006
rect 22204 16996 22260 18732
rect 22428 18562 22484 18574
rect 22428 18510 22430 18562
rect 22482 18510 22484 18562
rect 22428 18340 22484 18510
rect 22428 18274 22484 18284
rect 22092 16994 22260 16996
rect 22092 16942 22094 16994
rect 22146 16942 22260 16994
rect 22092 16940 22260 16942
rect 22092 16930 22148 16940
rect 21420 16146 21476 16156
rect 21756 16884 21812 16894
rect 21532 16100 21588 16110
rect 21532 15986 21588 16044
rect 21532 15934 21534 15986
rect 21586 15934 21588 15986
rect 21532 15922 21588 15934
rect 21644 15988 21700 15998
rect 21644 15894 21700 15932
rect 21308 15876 21364 15886
rect 21308 15782 21364 15820
rect 21420 15874 21476 15886
rect 21420 15822 21422 15874
rect 21474 15822 21476 15874
rect 21420 15652 21476 15822
rect 21756 15764 21812 16828
rect 22540 16772 22596 18732
rect 22652 17108 22708 20524
rect 22764 18788 22820 18798
rect 22764 18562 22820 18732
rect 22764 18510 22766 18562
rect 22818 18510 22820 18562
rect 22764 18498 22820 18510
rect 22764 17668 22820 17678
rect 22876 17668 22932 21644
rect 22988 21634 23044 21644
rect 23212 22148 23268 22158
rect 23212 20802 23268 22092
rect 24444 21364 24500 22316
rect 24668 22306 24724 22316
rect 24220 21308 24500 21364
rect 24220 21026 24276 21308
rect 24220 20974 24222 21026
rect 24274 20974 24276 21026
rect 24220 20962 24276 20974
rect 23884 20916 23940 20926
rect 23884 20822 23940 20860
rect 23212 20750 23214 20802
rect 23266 20750 23268 20802
rect 23212 20738 23268 20750
rect 22988 20692 23044 20702
rect 22988 20598 23044 20636
rect 24108 20580 24164 20590
rect 24108 20486 24164 20524
rect 23212 20244 23268 20254
rect 23212 20150 23268 20188
rect 23772 20130 23828 20142
rect 23772 20078 23774 20130
rect 23826 20078 23828 20130
rect 22988 20020 23044 20030
rect 22988 19236 23044 19964
rect 23660 19460 23716 19470
rect 23660 19366 23716 19404
rect 23100 19236 23156 19246
rect 22988 19234 23156 19236
rect 22988 19182 23102 19234
rect 23154 19182 23156 19234
rect 22988 19180 23156 19182
rect 23100 19170 23156 19180
rect 23324 19234 23380 19246
rect 23324 19182 23326 19234
rect 23378 19182 23380 19234
rect 23100 18676 23156 18686
rect 23100 18450 23156 18620
rect 23100 18398 23102 18450
rect 23154 18398 23156 18450
rect 23100 18386 23156 18398
rect 23324 18452 23380 19182
rect 23548 19234 23604 19246
rect 23772 19236 23828 20078
rect 23548 19182 23550 19234
rect 23602 19182 23604 19234
rect 23548 18788 23604 19182
rect 23548 18722 23604 18732
rect 23660 19180 23828 19236
rect 23996 20018 24052 20030
rect 23996 19966 23998 20018
rect 24050 19966 24052 20018
rect 23548 18564 23604 18574
rect 23660 18564 23716 19180
rect 23604 18508 23716 18564
rect 23548 18470 23604 18508
rect 23324 18386 23380 18396
rect 23436 18450 23492 18462
rect 23436 18398 23438 18450
rect 23490 18398 23492 18450
rect 22764 17666 22932 17668
rect 22764 17614 22766 17666
rect 22818 17614 22932 17666
rect 22764 17612 22932 17614
rect 22988 18340 23044 18350
rect 22764 17602 22820 17612
rect 22652 16882 22708 17052
rect 22988 17106 23044 18284
rect 23100 18226 23156 18238
rect 23100 18174 23102 18226
rect 23154 18174 23156 18226
rect 23100 18116 23156 18174
rect 23436 18116 23492 18398
rect 23772 18452 23828 18462
rect 23772 18358 23828 18396
rect 23100 18060 23492 18116
rect 23996 18116 24052 19966
rect 24332 18452 24388 18462
rect 22988 17054 22990 17106
rect 23042 17054 23044 17106
rect 22988 17042 23044 17054
rect 23100 17892 23156 17902
rect 23100 17106 23156 17836
rect 23100 17054 23102 17106
rect 23154 17054 23156 17106
rect 23100 17042 23156 17054
rect 22652 16830 22654 16882
rect 22706 16830 22708 16882
rect 22652 16818 22708 16830
rect 22764 16882 22820 16894
rect 22764 16830 22766 16882
rect 22818 16830 22820 16882
rect 21420 15586 21476 15596
rect 21532 15708 21812 15764
rect 21980 16660 22036 16670
rect 21532 15538 21588 15708
rect 21868 15652 21924 15662
rect 21532 15486 21534 15538
rect 21586 15486 21588 15538
rect 21532 15474 21588 15486
rect 21644 15540 21700 15550
rect 21644 15446 21700 15484
rect 21868 15538 21924 15596
rect 21868 15486 21870 15538
rect 21922 15486 21924 15538
rect 21868 15474 21924 15486
rect 21980 15540 22036 16604
rect 22540 16548 22596 16716
rect 22764 16660 22820 16830
rect 22876 16772 22932 16782
rect 22876 16678 22932 16716
rect 22764 16594 22820 16604
rect 22540 16492 22708 16548
rect 22540 16324 22596 16334
rect 22092 16322 22596 16324
rect 22092 16270 22542 16322
rect 22594 16270 22596 16322
rect 22092 16268 22596 16270
rect 22092 16098 22148 16268
rect 22540 16258 22596 16268
rect 22092 16046 22094 16098
rect 22146 16046 22148 16098
rect 22092 16034 22148 16046
rect 22428 16100 22484 16110
rect 22428 16006 22484 16044
rect 22540 15988 22596 15998
rect 22652 15988 22708 16492
rect 22540 15986 22708 15988
rect 22540 15934 22542 15986
rect 22594 15934 22708 15986
rect 22540 15932 22708 15934
rect 22540 15922 22596 15932
rect 23324 15876 23380 18060
rect 23996 18050 24052 18060
rect 24220 18396 24332 18452
rect 24220 16994 24276 18396
rect 24332 18386 24388 18396
rect 24668 18340 24724 18350
rect 24668 17554 24724 18284
rect 24668 17502 24670 17554
rect 24722 17502 24724 17554
rect 24668 17490 24724 17502
rect 24220 16942 24222 16994
rect 24274 16942 24276 16994
rect 24220 16930 24276 16942
rect 24332 17106 24388 17118
rect 24332 17054 24334 17106
rect 24386 17054 24388 17106
rect 23996 16884 24052 16894
rect 23996 16790 24052 16828
rect 24108 16212 24164 16222
rect 24332 16212 24388 17054
rect 24668 16884 24724 16894
rect 24668 16790 24724 16828
rect 24108 16210 24388 16212
rect 24108 16158 24110 16210
rect 24162 16158 24388 16210
rect 24108 16156 24388 16158
rect 24108 16146 24164 16156
rect 23324 15810 23380 15820
rect 23436 16098 23492 16110
rect 23436 16046 23438 16098
rect 23490 16046 23492 16098
rect 21980 15474 22036 15484
rect 22092 15314 22148 15326
rect 22092 15262 22094 15314
rect 22146 15262 22148 15314
rect 21756 15202 21812 15214
rect 21756 15150 21758 15202
rect 21810 15150 21812 15202
rect 21084 15092 21140 15102
rect 21196 15092 21588 15148
rect 21084 14998 21140 15036
rect 20188 14914 20244 14924
rect 21532 14644 21588 15092
rect 21532 14578 21588 14588
rect 21756 14420 21812 15150
rect 22092 15148 22148 15262
rect 21868 15092 21924 15102
rect 22092 15092 22932 15148
rect 21868 14532 21924 15036
rect 21868 14438 21924 14476
rect 22092 14980 22148 14990
rect 22092 14644 22148 14924
rect 22876 14754 22932 15092
rect 22876 14702 22878 14754
rect 22930 14702 22932 14754
rect 22876 14690 22932 14702
rect 22092 14530 22148 14588
rect 22092 14478 22094 14530
rect 22146 14478 22148 14530
rect 22092 14466 22148 14478
rect 22540 14530 22596 14542
rect 22540 14478 22542 14530
rect 22594 14478 22596 14530
rect 21084 14364 21812 14420
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20300 13972 20356 13982
rect 20300 13746 20356 13916
rect 21084 13858 21140 14364
rect 21980 14306 22036 14318
rect 21980 14254 21982 14306
rect 22034 14254 22036 14306
rect 21084 13806 21086 13858
rect 21138 13806 21140 13858
rect 21084 13794 21140 13806
rect 21308 13972 21364 13982
rect 20300 13694 20302 13746
rect 20354 13694 20356 13746
rect 19740 13076 19796 13086
rect 19628 13074 19796 13076
rect 19628 13022 19742 13074
rect 19794 13022 19796 13074
rect 19628 13020 19796 13022
rect 19740 13010 19796 13020
rect 20300 13074 20356 13694
rect 20300 13022 20302 13074
rect 20354 13022 20356 13074
rect 20300 13010 20356 13022
rect 21308 12962 21364 13916
rect 21980 13076 22036 14254
rect 22540 13748 22596 14478
rect 22764 14532 22820 14542
rect 22764 14438 22820 14476
rect 22540 13682 22596 13692
rect 22876 14306 22932 14318
rect 22876 14254 22878 14306
rect 22930 14254 22932 14306
rect 22876 13636 22932 14254
rect 23436 14306 23492 16046
rect 24780 15148 24836 23212
rect 25340 23044 25396 23054
rect 25452 23044 25508 23886
rect 25564 23604 25620 24780
rect 37660 24724 37716 24734
rect 37660 24630 37716 24668
rect 40012 24498 40068 24510
rect 40012 24446 40014 24498
rect 40066 24446 40068 24498
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 40012 24276 40068 24446
rect 40012 24210 40068 24220
rect 26908 24052 26964 24062
rect 26236 23828 26292 23838
rect 25564 23538 25620 23548
rect 25788 23826 26292 23828
rect 25788 23774 26238 23826
rect 26290 23774 26292 23826
rect 25788 23772 26292 23774
rect 25788 23378 25844 23772
rect 26236 23762 26292 23772
rect 25788 23326 25790 23378
rect 25842 23326 25844 23378
rect 25788 23314 25844 23326
rect 26236 23604 26292 23614
rect 26236 23380 26292 23548
rect 26684 23380 26740 23390
rect 26908 23380 26964 23996
rect 28364 24052 28420 24062
rect 28364 23958 28420 23996
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 37660 23940 37716 23950
rect 37660 23846 37716 23884
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 26236 23324 26628 23380
rect 25676 23156 25732 23166
rect 25676 23062 25732 23100
rect 25900 23154 25956 23166
rect 25900 23102 25902 23154
rect 25954 23102 25956 23154
rect 25340 23042 25508 23044
rect 25340 22990 25342 23042
rect 25394 22990 25508 23042
rect 25340 22988 25508 22990
rect 25340 22484 25396 22988
rect 25340 22370 25396 22428
rect 25340 22318 25342 22370
rect 25394 22318 25396 22370
rect 25340 22306 25396 22318
rect 24892 22260 24948 22270
rect 24892 22166 24948 22204
rect 25004 22258 25060 22270
rect 25004 22206 25006 22258
rect 25058 22206 25060 22258
rect 25004 21812 25060 22206
rect 25004 21746 25060 21756
rect 25676 21588 25732 21598
rect 25676 21494 25732 21532
rect 25900 20244 25956 23102
rect 26124 22260 26180 22270
rect 26124 22166 26180 22204
rect 26124 21812 26180 21822
rect 26124 21718 26180 21756
rect 26012 21700 26068 21710
rect 26012 21586 26068 21644
rect 26236 21698 26292 23324
rect 26572 23266 26628 23324
rect 26684 23378 26964 23380
rect 26684 23326 26686 23378
rect 26738 23326 26964 23378
rect 26684 23324 26964 23326
rect 26684 23314 26740 23324
rect 26572 23214 26574 23266
rect 26626 23214 26628 23266
rect 26572 23202 26628 23214
rect 26348 23154 26404 23166
rect 26348 23102 26350 23154
rect 26402 23102 26404 23154
rect 26348 22932 26404 23102
rect 26684 22932 26740 22942
rect 26348 22930 26740 22932
rect 26348 22878 26686 22930
rect 26738 22878 26740 22930
rect 26348 22876 26740 22878
rect 26684 22866 26740 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 26236 21646 26238 21698
rect 26290 21646 26292 21698
rect 26236 21634 26292 21646
rect 28252 22484 28308 22494
rect 28252 21700 28308 22428
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 37660 22372 37716 22382
rect 37660 22278 37716 22316
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 28252 21634 28308 21644
rect 26012 21534 26014 21586
rect 26066 21534 26068 21586
rect 26012 21522 26068 21534
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 27356 20244 27412 20254
rect 25900 20178 25956 20188
rect 26348 20130 26404 20142
rect 26348 20078 26350 20130
rect 26402 20078 26404 20130
rect 25900 20020 25956 20030
rect 25676 19234 25732 19246
rect 25676 19182 25678 19234
rect 25730 19182 25732 19234
rect 25340 19012 25396 19022
rect 25676 19012 25732 19182
rect 25340 19010 25732 19012
rect 25340 18958 25342 19010
rect 25394 18958 25732 19010
rect 25340 18956 25732 18958
rect 25340 18340 25396 18956
rect 25900 18676 25956 19964
rect 26012 20018 26068 20030
rect 26012 19966 26014 20018
rect 26066 19966 26068 20018
rect 26012 19460 26068 19966
rect 26012 19394 26068 19404
rect 26348 20020 26404 20078
rect 27132 20132 27412 20188
rect 27468 20132 27748 20188
rect 26572 20020 26628 20030
rect 26348 20018 26628 20020
rect 26348 19966 26574 20018
rect 26626 19966 26628 20018
rect 26348 19964 26628 19966
rect 25900 18582 25956 18620
rect 25452 18452 25508 18462
rect 25452 18358 25508 18396
rect 25676 18450 25732 18462
rect 25676 18398 25678 18450
rect 25730 18398 25732 18450
rect 25340 18274 25396 18284
rect 25676 17892 25732 18398
rect 25788 18452 25844 18462
rect 25788 18358 25844 18396
rect 26124 18452 26180 18462
rect 26348 18452 26404 19964
rect 26572 19954 26628 19964
rect 26908 20020 26964 20030
rect 26908 19926 26964 19964
rect 26796 19906 26852 19918
rect 26796 19854 26798 19906
rect 26850 19854 26852 19906
rect 26460 19348 26516 19358
rect 26796 19348 26852 19854
rect 27132 19796 27188 20132
rect 27244 20020 27300 20030
rect 27468 20020 27524 20132
rect 27692 20130 27748 20132
rect 27692 20078 27694 20130
rect 27746 20078 27748 20130
rect 27692 20066 27748 20078
rect 27244 20018 27524 20020
rect 27244 19966 27246 20018
rect 27298 19966 27524 20018
rect 27244 19964 27524 19966
rect 27580 20018 27636 20030
rect 27580 19966 27582 20018
rect 27634 19966 27636 20018
rect 27244 19954 27300 19964
rect 27580 19796 27636 19966
rect 27916 20020 27972 20030
rect 27916 19926 27972 19964
rect 28028 20018 28084 20030
rect 28028 19966 28030 20018
rect 28082 19966 28084 20018
rect 27132 19740 27636 19796
rect 26460 19346 26852 19348
rect 26460 19294 26462 19346
rect 26514 19294 26852 19346
rect 26460 19292 26852 19294
rect 26460 19282 26516 19292
rect 26124 18450 26404 18452
rect 26124 18398 26126 18450
rect 26178 18398 26404 18450
rect 26124 18396 26404 18398
rect 26460 18450 26516 18462
rect 26460 18398 26462 18450
rect 26514 18398 26516 18450
rect 25676 17826 25732 17836
rect 25228 17108 25284 17118
rect 25228 16994 25284 17052
rect 25228 16942 25230 16994
rect 25282 16942 25284 16994
rect 25228 16930 25284 16942
rect 25340 16996 25396 17006
rect 25340 16902 25396 16940
rect 25564 16884 25620 16894
rect 25564 16790 25620 16828
rect 26124 16100 26180 18396
rect 26460 18340 26516 18398
rect 27244 18452 27300 18462
rect 27244 18358 27300 18396
rect 26460 17106 26516 18284
rect 27020 17892 27076 17902
rect 27020 17666 27076 17836
rect 27020 17614 27022 17666
rect 27074 17614 27076 17666
rect 27020 17602 27076 17614
rect 27356 17668 27412 17678
rect 27580 17668 27636 19740
rect 28028 19460 28084 19966
rect 28028 19394 28084 19404
rect 28588 20020 28644 20030
rect 28588 19346 28644 19964
rect 37660 20020 37716 20030
rect 37660 19926 37716 19964
rect 40012 19794 40068 19806
rect 40012 19742 40014 19794
rect 40066 19742 40068 19794
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 40012 19572 40068 19742
rect 40012 19506 40068 19516
rect 28588 19294 28590 19346
rect 28642 19294 28644 19346
rect 28588 19282 28644 19294
rect 40012 19346 40068 19358
rect 40012 19294 40014 19346
rect 40066 19294 40068 19346
rect 29260 19234 29316 19246
rect 29260 19182 29262 19234
rect 29314 19182 29316 19234
rect 29260 18900 29316 19182
rect 37660 19234 37716 19246
rect 37660 19182 37662 19234
rect 37714 19182 37716 19234
rect 29484 19012 29540 19022
rect 29484 18918 29540 18956
rect 37660 18900 37716 19182
rect 29316 18844 29428 18900
rect 29260 18834 29316 18844
rect 27356 17666 27636 17668
rect 27356 17614 27358 17666
rect 27410 17614 27636 17666
rect 27356 17612 27636 17614
rect 29372 18338 29428 18844
rect 37660 18834 37716 18844
rect 37884 19012 37940 19022
rect 37884 18450 37940 18956
rect 40012 18900 40068 19294
rect 40012 18834 40068 18844
rect 37884 18398 37886 18450
rect 37938 18398 37940 18450
rect 37884 18386 37940 18398
rect 29372 18286 29374 18338
rect 29426 18286 29428 18338
rect 27356 17602 27412 17612
rect 27244 17556 27300 17566
rect 27244 17462 27300 17500
rect 29372 17556 29428 18286
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 29372 17490 29428 17500
rect 37660 17666 37716 17678
rect 37660 17614 37662 17666
rect 37714 17614 37716 17666
rect 26460 17054 26462 17106
rect 26514 17054 26516 17106
rect 26236 16996 26292 17006
rect 26236 16210 26292 16940
rect 26236 16158 26238 16210
rect 26290 16158 26292 16210
rect 26236 16146 26292 16158
rect 26124 16034 26180 16044
rect 23436 14254 23438 14306
rect 23490 14254 23492 14306
rect 23436 13972 23492 14254
rect 24556 15092 24836 15148
rect 26012 15316 26068 15326
rect 26460 15316 26516 17054
rect 37660 16996 37716 17614
rect 37660 16930 37716 16940
rect 40012 16884 40068 17726
rect 40012 16818 40068 16828
rect 26684 16772 26740 16782
rect 26684 16098 26740 16716
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 27132 16212 27188 16222
rect 27132 16210 27748 16212
rect 27132 16158 27134 16210
rect 27186 16158 27748 16210
rect 27132 16156 27748 16158
rect 27132 16146 27188 16156
rect 26684 16046 26686 16098
rect 26738 16046 26740 16098
rect 26684 16034 26740 16046
rect 26796 16100 26852 16110
rect 26908 16100 26964 16110
rect 26852 16098 26964 16100
rect 26852 16046 26910 16098
rect 26962 16046 26964 16098
rect 26852 16044 26964 16046
rect 26012 15314 26516 15316
rect 26012 15262 26014 15314
rect 26066 15262 26462 15314
rect 26514 15262 26516 15314
rect 26012 15260 26516 15262
rect 24556 14868 24612 15092
rect 23436 13906 23492 13916
rect 23660 13972 23716 13982
rect 24332 13972 24388 13982
rect 24556 13972 24612 14812
rect 23660 13970 23940 13972
rect 23660 13918 23662 13970
rect 23714 13918 23940 13970
rect 23660 13916 23940 13918
rect 23660 13906 23716 13916
rect 23436 13748 23492 13758
rect 23436 13654 23492 13692
rect 23772 13748 23828 13758
rect 23772 13654 23828 13692
rect 23212 13636 23268 13646
rect 22876 13634 23268 13636
rect 22876 13582 23214 13634
rect 23266 13582 23268 13634
rect 22876 13580 23268 13582
rect 22092 13076 22148 13086
rect 21980 13074 22148 13076
rect 21980 13022 22094 13074
rect 22146 13022 22148 13074
rect 21980 13020 22148 13022
rect 22092 13010 22148 13020
rect 21308 12910 21310 12962
rect 21362 12910 21364 12962
rect 21308 12898 21364 12910
rect 16828 12684 17444 12740
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 16828 8428 16884 12684
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 16828 8372 18004 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 17500 3668 17556 3678
rect 17500 800 17556 3612
rect 17948 3554 18004 8372
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19068 4452 19124 4462
rect 18844 4450 19124 4452
rect 18844 4398 19070 4450
rect 19122 4398 19124 4450
rect 18844 4396 19124 4398
rect 18620 3668 18676 3678
rect 18620 3574 18676 3612
rect 17948 3502 17950 3554
rect 18002 3502 18004 3554
rect 17948 3490 18004 3502
rect 18844 800 18900 4396
rect 19068 4386 19124 4396
rect 23212 3556 23268 13580
rect 23884 13076 23940 13916
rect 24332 13970 24612 13972
rect 24332 13918 24334 13970
rect 24386 13918 24612 13970
rect 24332 13916 24612 13918
rect 24668 13972 24724 13982
rect 26012 13972 26068 15260
rect 26460 15250 26516 15260
rect 26460 14756 26516 14766
rect 26796 14756 26852 16044
rect 26908 16034 26964 16044
rect 27244 15986 27300 15998
rect 27244 15934 27246 15986
rect 27298 15934 27300 15986
rect 27132 15428 27188 15438
rect 27244 15428 27300 15934
rect 27132 15426 27300 15428
rect 27132 15374 27134 15426
rect 27186 15374 27300 15426
rect 27132 15372 27300 15374
rect 27132 15362 27188 15372
rect 26460 14754 26852 14756
rect 26460 14702 26462 14754
rect 26514 14702 26852 14754
rect 26460 14700 26852 14702
rect 26460 14690 26516 14700
rect 26124 14644 26180 14654
rect 26124 14550 26180 14588
rect 27692 14642 27748 16156
rect 40012 16210 40068 16222
rect 40012 16158 40014 16210
rect 40066 16158 40068 16210
rect 37660 16098 37716 16110
rect 37660 16046 37662 16098
rect 37714 16046 37716 16098
rect 27692 14590 27694 14642
rect 27746 14590 27748 14642
rect 27692 14578 27748 14590
rect 27916 15204 27972 15214
rect 26236 14532 26292 14542
rect 26236 14438 26292 14476
rect 27020 14532 27076 14542
rect 27020 14438 27076 14476
rect 27244 14530 27300 14542
rect 27244 14478 27246 14530
rect 27298 14478 27300 14530
rect 26908 14420 26964 14430
rect 26908 14326 26964 14364
rect 24724 13916 24836 13972
rect 24332 13748 24388 13916
rect 24668 13878 24724 13916
rect 24332 13682 24388 13692
rect 24780 13748 24836 13916
rect 26012 13906 26068 13916
rect 26124 14306 26180 14318
rect 26124 14254 26126 14306
rect 26178 14254 26180 14306
rect 26124 13858 26180 14254
rect 27244 14308 27300 14478
rect 27916 14530 27972 15148
rect 29260 15204 29316 15214
rect 29260 15110 29316 15148
rect 37660 15204 37716 16046
rect 40012 15540 40068 16158
rect 40012 15474 40068 15484
rect 37660 15138 37716 15148
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 40012 14642 40068 14654
rect 40012 14590 40014 14642
rect 40066 14590 40068 14642
rect 27916 14478 27918 14530
rect 27970 14478 27972 14530
rect 27916 14466 27972 14478
rect 37660 14532 37716 14542
rect 37660 14438 37716 14476
rect 27580 14420 27636 14430
rect 27580 14326 27636 14364
rect 27244 14242 27300 14252
rect 28252 14308 28308 14318
rect 26124 13806 26126 13858
rect 26178 13806 26180 13858
rect 26124 13794 26180 13806
rect 25340 13748 25396 13758
rect 24780 13746 25396 13748
rect 24780 13694 25342 13746
rect 25394 13694 25396 13746
rect 24780 13692 25396 13694
rect 24220 13076 24276 13086
rect 23884 13074 24276 13076
rect 23884 13022 24222 13074
rect 24274 13022 24276 13074
rect 23884 13020 24276 13022
rect 24220 8428 24276 13020
rect 24780 13074 24836 13692
rect 25340 13682 25396 13692
rect 28252 13634 28308 14252
rect 40012 14196 40068 14590
rect 40012 14130 40068 14140
rect 28252 13582 28254 13634
rect 28306 13582 28308 13634
rect 28252 13570 28308 13582
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 24780 13022 24782 13074
rect 24834 13022 24836 13074
rect 24780 13010 24836 13022
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 24220 8372 24612 8428
rect 23772 3668 23828 3678
rect 23548 3556 23604 3566
rect 23212 3554 23604 3556
rect 23212 3502 23550 3554
rect 23602 3502 23604 3554
rect 23212 3500 23604 3502
rect 23548 3490 23604 3500
rect 22204 3442 22260 3454
rect 22204 3390 22206 3442
rect 22258 3390 22260 3442
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 22204 800 22260 3390
rect 23772 980 23828 3612
rect 24556 3554 24612 8372
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 23548 924 23828 980
rect 23548 800 23604 924
rect 17472 0 17584 800
rect 18816 0 18928 800
rect 22176 0 22288 800
rect 23520 0 23632 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 16828 37436 16884 37492
rect 18396 37490 18452 37492
rect 18396 37438 18398 37490
rect 18398 37438 18450 37490
rect 18450 37438 18452 37490
rect 18396 37436 18452 37438
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4172 27580 4228 27636
rect 1932 26236 1988 26292
rect 1932 25564 1988 25620
rect 2044 24892 2100 24948
rect 1932 22930 1988 22932
rect 1932 22878 1934 22930
rect 1934 22878 1986 22930
rect 1986 22878 1988 22930
rect 1932 22876 1988 22878
rect 1932 20860 1988 20916
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4284 27074 4340 27076
rect 4284 27022 4286 27074
rect 4286 27022 4338 27074
rect 4338 27022 4340 27074
rect 4284 27020 4340 27022
rect 14364 27020 14420 27076
rect 4284 26290 4340 26292
rect 4284 26238 4286 26290
rect 4286 26238 4338 26290
rect 4338 26238 4340 26290
rect 4284 26236 4340 26238
rect 12572 26236 12628 26292
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4284 25506 4340 25508
rect 4284 25454 4286 25506
rect 4286 25454 4338 25506
rect 4338 25454 4340 25506
rect 4284 25452 4340 25454
rect 11452 25452 11508 25508
rect 12796 25506 12852 25508
rect 12796 25454 12798 25506
rect 12798 25454 12850 25506
rect 12850 25454 12852 25506
rect 12796 25452 12852 25454
rect 13804 25282 13860 25284
rect 13804 25230 13806 25282
rect 13806 25230 13858 25282
rect 13858 25230 13860 25282
rect 13804 25228 13860 25230
rect 16604 26348 16660 26404
rect 14700 26178 14756 26180
rect 14700 26126 14702 26178
rect 14702 26126 14754 26178
rect 14754 26126 14756 26178
rect 14700 26124 14756 26126
rect 15820 26124 15876 26180
rect 18060 27580 18116 27636
rect 18956 27634 19012 27636
rect 18956 27582 18958 27634
rect 18958 27582 19010 27634
rect 19010 27582 19012 27634
rect 18956 27580 19012 27582
rect 14588 25506 14644 25508
rect 14588 25454 14590 25506
rect 14590 25454 14642 25506
rect 14642 25454 14644 25506
rect 14588 25452 14644 25454
rect 14252 24556 14308 24612
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 15932 25394 15988 25396
rect 15932 25342 15934 25394
rect 15934 25342 15986 25394
rect 15986 25342 15988 25394
rect 15932 25340 15988 25342
rect 15484 24610 15540 24612
rect 15484 24558 15486 24610
rect 15486 24558 15538 24610
rect 15538 24558 15540 24610
rect 15484 24556 15540 24558
rect 4284 23154 4340 23156
rect 4284 23102 4286 23154
rect 4286 23102 4338 23154
rect 4338 23102 4340 23154
rect 4284 23100 4340 23102
rect 11004 23100 11060 23156
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 13132 21756 13188 21812
rect 4284 21586 4340 21588
rect 4284 21534 4286 21586
rect 4286 21534 4338 21586
rect 4338 21534 4340 21586
rect 4284 21532 4340 21534
rect 10556 21532 10612 21588
rect 14028 22988 14084 23044
rect 14476 23100 14532 23156
rect 14364 22316 14420 22372
rect 14140 21810 14196 21812
rect 14140 21758 14142 21810
rect 14142 21758 14194 21810
rect 14194 21758 14196 21810
rect 14140 21756 14196 21758
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 12236 20914 12292 20916
rect 12236 20862 12238 20914
rect 12238 20862 12290 20914
rect 12290 20862 12292 20914
rect 12236 20860 12292 20862
rect 4172 20524 4228 20580
rect 13692 20188 13748 20244
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4284 19234 4340 19236
rect 4284 19182 4286 19234
rect 4286 19182 4338 19234
rect 4338 19182 4340 19234
rect 4284 19180 4340 19182
rect 1932 18844 1988 18900
rect 4284 18450 4340 18452
rect 4284 18398 4286 18450
rect 4286 18398 4338 18450
rect 4338 18398 4340 18450
rect 4284 18396 4340 18398
rect 10892 18396 10948 18452
rect 11452 19180 11508 19236
rect 11452 18508 11508 18564
rect 1932 18226 1988 18228
rect 1932 18174 1934 18226
rect 1934 18174 1986 18226
rect 1986 18174 1988 18226
rect 1932 18172 1988 18174
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 14812 23154 14868 23156
rect 14812 23102 14814 23154
rect 14814 23102 14866 23154
rect 14866 23102 14868 23154
rect 14812 23100 14868 23102
rect 14364 21532 14420 21588
rect 14028 21420 14084 21476
rect 14140 20914 14196 20916
rect 14140 20862 14142 20914
rect 14142 20862 14194 20914
rect 14194 20862 14196 20914
rect 14140 20860 14196 20862
rect 14924 21420 14980 21476
rect 15148 22988 15204 23044
rect 15932 23100 15988 23156
rect 14252 20242 14308 20244
rect 14252 20190 14254 20242
rect 14254 20190 14306 20242
rect 14306 20190 14308 20242
rect 14252 20188 14308 20190
rect 14140 19404 14196 19460
rect 15708 21420 15764 21476
rect 16828 25394 16884 25396
rect 16828 25342 16830 25394
rect 16830 25342 16882 25394
rect 16882 25342 16884 25394
rect 16828 25340 16884 25342
rect 17164 25340 17220 25396
rect 17724 25394 17780 25396
rect 17724 25342 17726 25394
rect 17726 25342 17778 25394
rect 17778 25342 17780 25394
rect 17724 25340 17780 25342
rect 16716 25282 16772 25284
rect 16716 25230 16718 25282
rect 16718 25230 16770 25282
rect 16770 25230 16772 25282
rect 16716 25228 16772 25230
rect 18060 24556 18116 24612
rect 16492 23154 16548 23156
rect 16492 23102 16494 23154
rect 16494 23102 16546 23154
rect 16546 23102 16548 23154
rect 16492 23100 16548 23102
rect 17948 23266 18004 23268
rect 17948 23214 17950 23266
rect 17950 23214 18002 23266
rect 18002 23214 18004 23266
rect 17948 23212 18004 23214
rect 16828 23154 16884 23156
rect 16828 23102 16830 23154
rect 16830 23102 16882 23154
rect 16882 23102 16884 23154
rect 16828 23100 16884 23102
rect 17836 23154 17892 23156
rect 17836 23102 17838 23154
rect 17838 23102 17890 23154
rect 17890 23102 17892 23154
rect 17836 23100 17892 23102
rect 17500 22428 17556 22484
rect 18060 22428 18116 22484
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 24892 38220 24948 38276
rect 20188 37436 20244 37492
rect 21420 37490 21476 37492
rect 21420 37438 21422 37490
rect 21422 37438 21474 37490
rect 21474 37438 21476 37490
rect 21420 37436 21476 37438
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19516 28082 19572 28084
rect 19516 28030 19518 28082
rect 19518 28030 19570 28082
rect 19570 28030 19572 28082
rect 19516 28028 19572 28030
rect 20412 28028 20468 28084
rect 22428 27804 22484 27860
rect 20636 27074 20692 27076
rect 20636 27022 20638 27074
rect 20638 27022 20690 27074
rect 20690 27022 20692 27074
rect 20636 27020 20692 27022
rect 19404 26124 19460 26180
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20300 26178 20356 26180
rect 20300 26126 20302 26178
rect 20302 26126 20354 26178
rect 20354 26126 20356 26178
rect 20300 26124 20356 26126
rect 19516 25506 19572 25508
rect 19516 25454 19518 25506
rect 19518 25454 19570 25506
rect 19570 25454 19572 25506
rect 19516 25452 19572 25454
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 21980 27692 22036 27748
rect 21420 26124 21476 26180
rect 22204 26402 22260 26404
rect 22204 26350 22206 26402
rect 22206 26350 22258 26402
rect 22258 26350 22260 26402
rect 22204 26348 22260 26350
rect 21980 26236 22036 26292
rect 21644 25452 21700 25508
rect 22092 26124 22148 26180
rect 20524 23938 20580 23940
rect 20524 23886 20526 23938
rect 20526 23886 20578 23938
rect 20578 23886 20580 23938
rect 20524 23884 20580 23886
rect 21532 23938 21588 23940
rect 21532 23886 21534 23938
rect 21534 23886 21586 23938
rect 21586 23886 21588 23938
rect 21532 23884 21588 23886
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19292 23212 19348 23268
rect 20188 23212 20244 23268
rect 18508 22316 18564 22372
rect 19836 21978 19892 21980
rect 17052 21868 17108 21924
rect 18172 21868 18228 21924
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 16604 21420 16660 21476
rect 13916 19234 13972 19236
rect 13916 19182 13918 19234
rect 13918 19182 13970 19234
rect 13970 19182 13972 19234
rect 13916 19180 13972 19182
rect 13692 18956 13748 19012
rect 13804 17836 13860 17892
rect 14700 18674 14756 18676
rect 14700 18622 14702 18674
rect 14702 18622 14754 18674
rect 14754 18622 14756 18674
rect 14700 18620 14756 18622
rect 15372 19122 15428 19124
rect 15372 19070 15374 19122
rect 15374 19070 15426 19122
rect 15426 19070 15428 19122
rect 15372 19068 15428 19070
rect 16044 20018 16100 20020
rect 16044 19966 16046 20018
rect 16046 19966 16098 20018
rect 16098 19966 16100 20018
rect 16044 19964 16100 19966
rect 16044 19404 16100 19460
rect 15596 18620 15652 18676
rect 14924 18562 14980 18564
rect 14924 18510 14926 18562
rect 14926 18510 14978 18562
rect 14978 18510 14980 18562
rect 14924 18508 14980 18510
rect 17388 21420 17444 21476
rect 19068 21586 19124 21588
rect 19068 21534 19070 21586
rect 19070 21534 19122 21586
rect 19122 21534 19124 21586
rect 19068 21532 19124 21534
rect 17724 21420 17780 21476
rect 18620 21474 18676 21476
rect 18620 21422 18622 21474
rect 18622 21422 18674 21474
rect 18674 21422 18676 21474
rect 18620 21420 18676 21422
rect 16156 19122 16212 19124
rect 16156 19070 16158 19122
rect 16158 19070 16210 19122
rect 16210 19070 16212 19122
rect 16156 19068 16212 19070
rect 15820 18562 15876 18564
rect 15820 18510 15822 18562
rect 15822 18510 15874 18562
rect 15874 18510 15876 18562
rect 15820 18508 15876 18510
rect 14700 18396 14756 18452
rect 14028 17948 14084 18004
rect 14476 17948 14532 18004
rect 14924 17890 14980 17892
rect 14924 17838 14926 17890
rect 14926 17838 14978 17890
rect 14978 17838 14980 17890
rect 14924 17836 14980 17838
rect 15372 17612 15428 17668
rect 14700 17052 14756 17108
rect 16268 18450 16324 18452
rect 16268 18398 16270 18450
rect 16270 18398 16322 18450
rect 16322 18398 16324 18450
rect 16268 18396 16324 18398
rect 17500 20860 17556 20916
rect 16716 18284 16772 18340
rect 17164 18508 17220 18564
rect 16716 17666 16772 17668
rect 16716 17614 16718 17666
rect 16718 17614 16770 17666
rect 16770 17614 16772 17666
rect 16716 17612 16772 17614
rect 17388 18396 17444 18452
rect 16044 17052 16100 17108
rect 17276 16828 17332 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 17388 17500 17444 17556
rect 16828 16770 16884 16772
rect 16828 16718 16830 16770
rect 16830 16718 16882 16770
rect 16882 16718 16884 16770
rect 16828 16716 16884 16718
rect 18060 20242 18116 20244
rect 18060 20190 18062 20242
rect 18062 20190 18114 20242
rect 18114 20190 18116 20242
rect 18060 20188 18116 20190
rect 18620 20636 18676 20692
rect 17724 20130 17780 20132
rect 17724 20078 17726 20130
rect 17726 20078 17778 20130
rect 17778 20078 17780 20130
rect 17724 20076 17780 20078
rect 18396 19964 18452 20020
rect 18508 20076 18564 20132
rect 20076 20802 20132 20804
rect 20076 20750 20078 20802
rect 20078 20750 20130 20802
rect 20130 20750 20132 20802
rect 20076 20748 20132 20750
rect 19180 20524 19236 20580
rect 18732 20130 18788 20132
rect 18732 20078 18734 20130
rect 18734 20078 18786 20130
rect 18786 20078 18788 20130
rect 18732 20076 18788 20078
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19516 18620 19572 18676
rect 18508 18562 18564 18564
rect 18508 18510 18510 18562
rect 18510 18510 18562 18562
rect 18562 18510 18564 18562
rect 18508 18508 18564 18510
rect 18172 18396 18228 18452
rect 19292 18338 19348 18340
rect 19292 18286 19294 18338
rect 19294 18286 19346 18338
rect 19346 18286 19348 18338
rect 19292 18284 19348 18286
rect 18508 17666 18564 17668
rect 18508 17614 18510 17666
rect 18510 17614 18562 17666
rect 18562 17614 18564 17666
rect 18508 17612 18564 17614
rect 17724 17052 17780 17108
rect 16492 14530 16548 14532
rect 16492 14478 16494 14530
rect 16494 14478 16546 14530
rect 16546 14478 16548 14530
rect 16492 14476 16548 14478
rect 14028 13916 14084 13972
rect 14700 14252 14756 14308
rect 16380 14306 16436 14308
rect 16380 14254 16382 14306
rect 16382 14254 16434 14306
rect 16434 14254 16436 14306
rect 16380 14252 16436 14254
rect 17164 14700 17220 14756
rect 17276 14476 17332 14532
rect 17836 16716 17892 16772
rect 17948 16828 18004 16884
rect 18284 16716 18340 16772
rect 19628 20076 19684 20132
rect 21756 22428 21812 22484
rect 21868 23436 21924 23492
rect 20748 21980 20804 22036
rect 20860 21532 20916 21588
rect 20636 20748 20692 20804
rect 20636 20300 20692 20356
rect 20300 20188 20356 20244
rect 20524 20188 20580 20244
rect 20412 20130 20468 20132
rect 20412 20078 20414 20130
rect 20414 20078 20466 20130
rect 20466 20078 20468 20130
rect 20412 20076 20468 20078
rect 20188 19794 20244 19796
rect 20188 19742 20190 19794
rect 20190 19742 20242 19794
rect 20242 19742 20244 19794
rect 20188 19740 20244 19742
rect 20412 19740 20468 19796
rect 20076 19010 20132 19012
rect 20076 18958 20078 19010
rect 20078 18958 20130 19010
rect 20130 18958 20132 19010
rect 20076 18956 20132 18958
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19628 18562 19684 18564
rect 19628 18510 19630 18562
rect 19630 18510 19682 18562
rect 19682 18510 19684 18562
rect 19628 18508 19684 18510
rect 19516 17836 19572 17892
rect 19964 18284 20020 18340
rect 19292 17554 19348 17556
rect 19292 17502 19294 17554
rect 19294 17502 19346 17554
rect 19346 17502 19348 17554
rect 19292 17500 19348 17502
rect 18844 17052 18900 17108
rect 20300 18508 20356 18564
rect 20524 18338 20580 18340
rect 20524 18286 20526 18338
rect 20526 18286 20578 18338
rect 20578 18286 20580 18338
rect 20524 18284 20580 18286
rect 20188 17500 20244 17556
rect 18620 16044 18676 16100
rect 18732 15820 18788 15876
rect 17612 14530 17668 14532
rect 17612 14478 17614 14530
rect 17614 14478 17666 14530
rect 17666 14478 17668 14530
rect 17612 14476 17668 14478
rect 18060 14700 18116 14756
rect 18508 14530 18564 14532
rect 18508 14478 18510 14530
rect 18510 14478 18562 14530
rect 18562 14478 18564 14530
rect 18508 14476 18564 14478
rect 16940 13916 16996 13972
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 17500 13970 17556 13972
rect 17500 13918 17502 13970
rect 17502 13918 17554 13970
rect 17554 13918 17556 13970
rect 17500 13916 17556 13918
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20076 17052 20132 17108
rect 19852 16098 19908 16100
rect 19852 16046 19854 16098
rect 19854 16046 19906 16098
rect 19906 16046 19908 16098
rect 19852 16044 19908 16046
rect 20748 18450 20804 18452
rect 20748 18398 20750 18450
rect 20750 18398 20802 18450
rect 20802 18398 20804 18450
rect 20748 18396 20804 18398
rect 21644 22316 21700 22372
rect 21756 21980 21812 22036
rect 21980 22146 22036 22148
rect 21980 22094 21982 22146
rect 21982 22094 22034 22146
rect 22034 22094 22036 22146
rect 21980 22092 22036 22094
rect 21532 21532 21588 21588
rect 21420 20636 21476 20692
rect 21196 20130 21252 20132
rect 21196 20078 21198 20130
rect 21198 20078 21250 20130
rect 21250 20078 21252 20130
rect 21196 20076 21252 20078
rect 21532 20300 21588 20356
rect 21644 20130 21700 20132
rect 21644 20078 21646 20130
rect 21646 20078 21698 20130
rect 21698 20078 21700 20130
rect 21644 20076 21700 20078
rect 21420 18562 21476 18564
rect 21420 18510 21422 18562
rect 21422 18510 21474 18562
rect 21474 18510 21476 18562
rect 21420 18508 21476 18510
rect 21196 18172 21252 18228
rect 21196 17724 21252 17780
rect 21084 17500 21140 17556
rect 21868 20188 21924 20244
rect 22876 28476 22932 28532
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 26124 38274 26180 38276
rect 26124 38222 26126 38274
rect 26126 38222 26178 38274
rect 26178 38222 26180 38274
rect 26124 38220 26180 38222
rect 25788 37436 25844 37492
rect 26796 37490 26852 37492
rect 26796 37438 26798 37490
rect 26798 37438 26850 37490
rect 26850 37438 26852 37490
rect 26796 37436 26852 37438
rect 23772 28476 23828 28532
rect 23436 27916 23492 27972
rect 22876 27746 22932 27748
rect 22876 27694 22878 27746
rect 22878 27694 22930 27746
rect 22930 27694 22932 27746
rect 22876 27692 22932 27694
rect 23100 27692 23156 27748
rect 22652 27074 22708 27076
rect 22652 27022 22654 27074
rect 22654 27022 22706 27074
rect 22706 27022 22708 27074
rect 22652 27020 22708 27022
rect 23548 27858 23604 27860
rect 23548 27806 23550 27858
rect 23550 27806 23602 27858
rect 23602 27806 23604 27858
rect 23548 27804 23604 27806
rect 23772 26908 23828 26964
rect 23436 26348 23492 26404
rect 23324 26290 23380 26292
rect 23324 26238 23326 26290
rect 23326 26238 23378 26290
rect 23378 26238 23380 26290
rect 23324 26236 23380 26238
rect 23212 26178 23268 26180
rect 23212 26126 23214 26178
rect 23214 26126 23266 26178
rect 23266 26126 23268 26178
rect 23212 26124 23268 26126
rect 22428 25340 22484 25396
rect 22204 25228 22260 25284
rect 22316 24610 22372 24612
rect 22316 24558 22318 24610
rect 22318 24558 22370 24610
rect 22370 24558 22372 24610
rect 22316 24556 22372 24558
rect 23212 23436 23268 23492
rect 23324 24444 23380 24500
rect 22428 22316 22484 22372
rect 22540 20636 22596 20692
rect 22204 19740 22260 19796
rect 21868 18956 21924 19012
rect 22204 18732 22260 18788
rect 24332 27746 24388 27748
rect 24332 27694 24334 27746
rect 24334 27694 24386 27746
rect 24386 27694 24388 27746
rect 24332 27692 24388 27694
rect 25116 26908 25172 26964
rect 23996 26460 24052 26516
rect 25116 26514 25172 26516
rect 25116 26462 25118 26514
rect 25118 26462 25170 26514
rect 25170 26462 25172 26514
rect 25116 26460 25172 26462
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 23660 24834 23716 24836
rect 23660 24782 23662 24834
rect 23662 24782 23714 24834
rect 23714 24782 23716 24834
rect 23660 24780 23716 24782
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 25564 24780 25620 24836
rect 24108 24668 24164 24724
rect 24780 24668 24836 24724
rect 24220 24556 24276 24612
rect 24108 24498 24164 24500
rect 24108 24446 24110 24498
rect 24110 24446 24162 24498
rect 24162 24446 24164 24498
rect 24108 24444 24164 24446
rect 23548 22370 23604 22372
rect 23548 22318 23550 22370
rect 23550 22318 23602 22370
rect 23602 22318 23604 22370
rect 23548 22316 23604 22318
rect 23884 23100 23940 23156
rect 24332 22482 24388 22484
rect 24332 22430 24334 22482
rect 24334 22430 24386 22482
rect 24386 22430 24388 22482
rect 24332 22428 24388 22430
rect 22652 20524 22708 20580
rect 22540 19964 22596 20020
rect 21980 18620 22036 18676
rect 21644 18396 21700 18452
rect 22092 18450 22148 18452
rect 22092 18398 22094 18450
rect 22094 18398 22146 18450
rect 22146 18398 22148 18450
rect 22092 18396 22148 18398
rect 21532 17612 21588 17668
rect 20860 16716 20916 16772
rect 20300 15986 20356 15988
rect 20300 15934 20302 15986
rect 20302 15934 20354 15986
rect 20354 15934 20356 15986
rect 20300 15932 20356 15934
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20748 16156 20804 16212
rect 22428 18284 22484 18340
rect 21420 16156 21476 16212
rect 21756 16828 21812 16884
rect 21532 16044 21588 16100
rect 21644 15986 21700 15988
rect 21644 15934 21646 15986
rect 21646 15934 21698 15986
rect 21698 15934 21700 15986
rect 21644 15932 21700 15934
rect 21308 15874 21364 15876
rect 21308 15822 21310 15874
rect 21310 15822 21362 15874
rect 21362 15822 21364 15874
rect 21308 15820 21364 15822
rect 22764 18732 22820 18788
rect 23212 22092 23268 22148
rect 23884 20914 23940 20916
rect 23884 20862 23886 20914
rect 23886 20862 23938 20914
rect 23938 20862 23940 20914
rect 23884 20860 23940 20862
rect 22988 20690 23044 20692
rect 22988 20638 22990 20690
rect 22990 20638 23042 20690
rect 23042 20638 23044 20690
rect 22988 20636 23044 20638
rect 24108 20578 24164 20580
rect 24108 20526 24110 20578
rect 24110 20526 24162 20578
rect 24162 20526 24164 20578
rect 24108 20524 24164 20526
rect 23212 20242 23268 20244
rect 23212 20190 23214 20242
rect 23214 20190 23266 20242
rect 23266 20190 23268 20242
rect 23212 20188 23268 20190
rect 22988 20018 23044 20020
rect 22988 19966 22990 20018
rect 22990 19966 23042 20018
rect 23042 19966 23044 20018
rect 22988 19964 23044 19966
rect 23660 19458 23716 19460
rect 23660 19406 23662 19458
rect 23662 19406 23714 19458
rect 23714 19406 23716 19458
rect 23660 19404 23716 19406
rect 23100 18620 23156 18676
rect 23548 18732 23604 18788
rect 23548 18562 23604 18564
rect 23548 18510 23550 18562
rect 23550 18510 23602 18562
rect 23602 18510 23604 18562
rect 23548 18508 23604 18510
rect 23324 18396 23380 18452
rect 22988 18284 23044 18340
rect 22652 17052 22708 17108
rect 23772 18450 23828 18452
rect 23772 18398 23774 18450
rect 23774 18398 23826 18450
rect 23826 18398 23828 18450
rect 23772 18396 23828 18398
rect 23996 18060 24052 18116
rect 23100 17836 23156 17892
rect 22540 16716 22596 16772
rect 21420 15596 21476 15652
rect 21980 16658 22036 16660
rect 21980 16606 21982 16658
rect 21982 16606 22034 16658
rect 22034 16606 22036 16658
rect 21980 16604 22036 16606
rect 21868 15596 21924 15652
rect 21644 15538 21700 15540
rect 21644 15486 21646 15538
rect 21646 15486 21698 15538
rect 21698 15486 21700 15538
rect 21644 15484 21700 15486
rect 22876 16770 22932 16772
rect 22876 16718 22878 16770
rect 22878 16718 22930 16770
rect 22930 16718 22932 16770
rect 22876 16716 22932 16718
rect 22764 16604 22820 16660
rect 22428 16098 22484 16100
rect 22428 16046 22430 16098
rect 22430 16046 22482 16098
rect 22482 16046 22484 16098
rect 22428 16044 22484 16046
rect 24332 18396 24388 18452
rect 24668 18338 24724 18340
rect 24668 18286 24670 18338
rect 24670 18286 24722 18338
rect 24722 18286 24724 18338
rect 24668 18284 24724 18286
rect 23996 16882 24052 16884
rect 23996 16830 23998 16882
rect 23998 16830 24050 16882
rect 24050 16830 24052 16882
rect 23996 16828 24052 16830
rect 24668 16882 24724 16884
rect 24668 16830 24670 16882
rect 24670 16830 24722 16882
rect 24722 16830 24724 16882
rect 24668 16828 24724 16830
rect 23324 15820 23380 15876
rect 21980 15484 22036 15540
rect 21084 15090 21140 15092
rect 21084 15038 21086 15090
rect 21086 15038 21138 15090
rect 21138 15038 21140 15090
rect 21084 15036 21140 15038
rect 20188 14924 20244 14980
rect 21532 14588 21588 14644
rect 21868 15036 21924 15092
rect 21868 14530 21924 14532
rect 21868 14478 21870 14530
rect 21870 14478 21922 14530
rect 21922 14478 21924 14530
rect 21868 14476 21924 14478
rect 22092 14924 22148 14980
rect 22092 14588 22148 14644
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20300 13916 20356 13972
rect 21308 13916 21364 13972
rect 22764 14530 22820 14532
rect 22764 14478 22766 14530
rect 22766 14478 22818 14530
rect 22818 14478 22820 14530
rect 22764 14476 22820 14478
rect 22540 13692 22596 13748
rect 37660 24722 37716 24724
rect 37660 24670 37662 24722
rect 37662 24670 37714 24722
rect 37714 24670 37716 24722
rect 37660 24668 37716 24670
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 40012 24220 40068 24276
rect 26908 23996 26964 24052
rect 25564 23548 25620 23604
rect 26236 23548 26292 23604
rect 28364 24050 28420 24052
rect 28364 23998 28366 24050
rect 28366 23998 28418 24050
rect 28418 23998 28420 24050
rect 28364 23996 28420 23998
rect 37660 23938 37716 23940
rect 37660 23886 37662 23938
rect 37662 23886 37714 23938
rect 37714 23886 37716 23938
rect 37660 23884 37716 23886
rect 40012 23548 40068 23604
rect 25676 23154 25732 23156
rect 25676 23102 25678 23154
rect 25678 23102 25730 23154
rect 25730 23102 25732 23154
rect 25676 23100 25732 23102
rect 25340 22428 25396 22484
rect 24892 22258 24948 22260
rect 24892 22206 24894 22258
rect 24894 22206 24946 22258
rect 24946 22206 24948 22258
rect 24892 22204 24948 22206
rect 25004 21756 25060 21812
rect 25676 21586 25732 21588
rect 25676 21534 25678 21586
rect 25678 21534 25730 21586
rect 25730 21534 25732 21586
rect 25676 21532 25732 21534
rect 26124 22258 26180 22260
rect 26124 22206 26126 22258
rect 26126 22206 26178 22258
rect 26178 22206 26180 22258
rect 26124 22204 26180 22206
rect 26124 21810 26180 21812
rect 26124 21758 26126 21810
rect 26126 21758 26178 21810
rect 26178 21758 26180 21810
rect 26124 21756 26180 21758
rect 26012 21644 26068 21700
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 28252 22482 28308 22484
rect 28252 22430 28254 22482
rect 28254 22430 28306 22482
rect 28306 22430 28308 22482
rect 28252 22428 28308 22430
rect 37660 22370 37716 22372
rect 37660 22318 37662 22370
rect 37662 22318 37714 22370
rect 37714 22318 37716 22370
rect 37660 22316 37716 22318
rect 40012 22204 40068 22260
rect 28252 21644 28308 21700
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 25900 20188 25956 20244
rect 27356 20188 27412 20244
rect 25900 19964 25956 20020
rect 26012 19404 26068 19460
rect 25900 18674 25956 18676
rect 25900 18622 25902 18674
rect 25902 18622 25954 18674
rect 25954 18622 25956 18674
rect 25900 18620 25956 18622
rect 25452 18450 25508 18452
rect 25452 18398 25454 18450
rect 25454 18398 25506 18450
rect 25506 18398 25508 18450
rect 25452 18396 25508 18398
rect 25340 18284 25396 18340
rect 25788 18450 25844 18452
rect 25788 18398 25790 18450
rect 25790 18398 25842 18450
rect 25842 18398 25844 18450
rect 25788 18396 25844 18398
rect 26908 20018 26964 20020
rect 26908 19966 26910 20018
rect 26910 19966 26962 20018
rect 26962 19966 26964 20018
rect 26908 19964 26964 19966
rect 27916 20018 27972 20020
rect 27916 19966 27918 20018
rect 27918 19966 27970 20018
rect 27970 19966 27972 20018
rect 27916 19964 27972 19966
rect 25676 17836 25732 17892
rect 25228 17052 25284 17108
rect 25340 16994 25396 16996
rect 25340 16942 25342 16994
rect 25342 16942 25394 16994
rect 25394 16942 25396 16994
rect 25340 16940 25396 16942
rect 25564 16882 25620 16884
rect 25564 16830 25566 16882
rect 25566 16830 25618 16882
rect 25618 16830 25620 16882
rect 25564 16828 25620 16830
rect 27244 18450 27300 18452
rect 27244 18398 27246 18450
rect 27246 18398 27298 18450
rect 27298 18398 27300 18450
rect 27244 18396 27300 18398
rect 26460 18284 26516 18340
rect 27020 17836 27076 17892
rect 28028 19404 28084 19460
rect 28588 19964 28644 20020
rect 37660 20018 37716 20020
rect 37660 19966 37662 20018
rect 37662 19966 37714 20018
rect 37714 19966 37716 20018
rect 37660 19964 37716 19966
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 40012 19516 40068 19572
rect 29484 19010 29540 19012
rect 29484 18958 29486 19010
rect 29486 18958 29538 19010
rect 29538 18958 29540 19010
rect 29484 18956 29540 18958
rect 29260 18844 29316 18900
rect 37660 18844 37716 18900
rect 37884 18956 37940 19012
rect 40012 18844 40068 18900
rect 27244 17554 27300 17556
rect 27244 17502 27246 17554
rect 27246 17502 27298 17554
rect 27298 17502 27300 17554
rect 27244 17500 27300 17502
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 29372 17500 29428 17556
rect 26236 16940 26292 16996
rect 26124 16044 26180 16100
rect 37660 16940 37716 16996
rect 40012 16828 40068 16884
rect 26684 16716 26740 16772
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 26796 16044 26852 16100
rect 24556 14812 24612 14868
rect 23436 13916 23492 13972
rect 23436 13746 23492 13748
rect 23436 13694 23438 13746
rect 23438 13694 23490 13746
rect 23490 13694 23492 13746
rect 23436 13692 23492 13694
rect 23772 13746 23828 13748
rect 23772 13694 23774 13746
rect 23774 13694 23826 13746
rect 23826 13694 23828 13746
rect 23772 13692 23828 13694
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 17500 3612 17556 3668
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 18620 3666 18676 3668
rect 18620 3614 18622 3666
rect 18622 3614 18674 3666
rect 18674 3614 18676 3666
rect 18620 3612 18676 3614
rect 26124 14642 26180 14644
rect 26124 14590 26126 14642
rect 26126 14590 26178 14642
rect 26178 14590 26180 14642
rect 26124 14588 26180 14590
rect 27916 15148 27972 15204
rect 26236 14530 26292 14532
rect 26236 14478 26238 14530
rect 26238 14478 26290 14530
rect 26290 14478 26292 14530
rect 26236 14476 26292 14478
rect 27020 14530 27076 14532
rect 27020 14478 27022 14530
rect 27022 14478 27074 14530
rect 27074 14478 27076 14530
rect 27020 14476 27076 14478
rect 26908 14418 26964 14420
rect 26908 14366 26910 14418
rect 26910 14366 26962 14418
rect 26962 14366 26964 14418
rect 26908 14364 26964 14366
rect 24668 13970 24724 13972
rect 24668 13918 24670 13970
rect 24670 13918 24722 13970
rect 24722 13918 24724 13970
rect 24668 13916 24724 13918
rect 24332 13692 24388 13748
rect 26012 13916 26068 13972
rect 29260 15202 29316 15204
rect 29260 15150 29262 15202
rect 29262 15150 29314 15202
rect 29314 15150 29316 15202
rect 29260 15148 29316 15150
rect 40012 15484 40068 15540
rect 37660 15148 37716 15204
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 37660 14530 37716 14532
rect 37660 14478 37662 14530
rect 37662 14478 37714 14530
rect 37714 14478 37716 14530
rect 37660 14476 37716 14478
rect 27580 14418 27636 14420
rect 27580 14366 27582 14418
rect 27582 14366 27634 14418
rect 27634 14366 27636 14418
rect 27580 14364 27636 14366
rect 27244 14252 27300 14308
rect 28252 14252 28308 14308
rect 40012 14140 40068 14196
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 23772 3612 23828 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 24882 38220 24892 38276
rect 24948 38220 26124 38276
rect 26180 38220 26190 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 16818 37436 16828 37492
rect 16884 37436 18396 37492
rect 18452 37436 18462 37492
rect 20178 37436 20188 37492
rect 20244 37436 21420 37492
rect 21476 37436 21486 37492
rect 25778 37436 25788 37492
rect 25844 37436 26796 37492
rect 26852 37436 26862 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 22866 28476 22876 28532
rect 22932 28476 23772 28532
rect 23828 28476 23838 28532
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 19506 28028 19516 28084
rect 19572 28028 20412 28084
rect 20468 28028 20478 28084
rect 23398 27916 23436 27972
rect 23492 27916 23502 27972
rect 22418 27804 22428 27860
rect 22484 27804 23548 27860
rect 23604 27804 23614 27860
rect 21970 27692 21980 27748
rect 22036 27692 22876 27748
rect 22932 27692 22942 27748
rect 23090 27692 23100 27748
rect 23156 27692 24332 27748
rect 24388 27692 24398 27748
rect 0 27636 800 27664
rect 0 27580 4172 27636
rect 4228 27580 4238 27636
rect 18050 27580 18060 27636
rect 18116 27580 18956 27636
rect 19012 27580 19022 27636
rect 0 27552 800 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 4274 27020 4284 27076
rect 4340 27020 14364 27076
rect 14420 27020 14430 27076
rect 20626 27020 20636 27076
rect 20692 27020 22652 27076
rect 22708 27020 22718 27076
rect 23762 26908 23772 26964
rect 23828 26908 25116 26964
rect 25172 26908 25182 26964
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 23986 26460 23996 26516
rect 24052 26460 25116 26516
rect 25172 26460 25182 26516
rect 16594 26348 16604 26404
rect 16660 26348 22204 26404
rect 22260 26348 23436 26404
rect 23492 26348 23502 26404
rect 0 26292 800 26320
rect 0 26236 1932 26292
rect 1988 26236 1998 26292
rect 4274 26236 4284 26292
rect 4340 26236 12572 26292
rect 12628 26236 12638 26292
rect 21970 26236 21980 26292
rect 22036 26236 23324 26292
rect 23380 26236 23390 26292
rect 0 26208 800 26236
rect 14690 26124 14700 26180
rect 14756 26124 15820 26180
rect 15876 26124 15886 26180
rect 19394 26124 19404 26180
rect 19460 26124 20300 26180
rect 20356 26124 20366 26180
rect 21410 26124 21420 26180
rect 21476 26124 22092 26180
rect 22148 26124 22158 26180
rect 23202 26124 23212 26180
rect 23268 26124 23436 26180
rect 23492 26124 23502 26180
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 0 25620 800 25648
rect 0 25564 1932 25620
rect 1988 25564 1998 25620
rect 0 25536 800 25564
rect 4274 25452 4284 25508
rect 4340 25452 11452 25508
rect 11508 25452 12796 25508
rect 12852 25452 14588 25508
rect 14644 25452 14654 25508
rect 19506 25452 19516 25508
rect 19572 25452 21644 25508
rect 21700 25452 21710 25508
rect 15922 25340 15932 25396
rect 15988 25340 16828 25396
rect 16884 25340 16894 25396
rect 17154 25340 17164 25396
rect 17220 25340 17724 25396
rect 17780 25340 22428 25396
rect 22484 25340 22494 25396
rect 13794 25228 13804 25284
rect 13860 25228 16716 25284
rect 16772 25228 22204 25284
rect 22260 25228 22270 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 0 24948 800 24976
rect 0 24892 2044 24948
rect 2100 24892 2110 24948
rect 0 24864 800 24892
rect 23650 24780 23660 24836
rect 23716 24780 25564 24836
rect 25620 24780 25630 24836
rect 24098 24668 24108 24724
rect 24164 24668 24780 24724
rect 24836 24668 37660 24724
rect 37716 24668 37726 24724
rect 14242 24556 14252 24612
rect 14308 24556 15484 24612
rect 15540 24556 18060 24612
rect 18116 24556 18126 24612
rect 22306 24556 22316 24612
rect 22372 24556 24220 24612
rect 24276 24556 24286 24612
rect 23314 24444 23324 24500
rect 23380 24444 24108 24500
rect 24164 24444 24174 24500
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 41200 24276 42000 24304
rect 40002 24220 40012 24276
rect 40068 24220 42000 24276
rect 41200 24192 42000 24220
rect 26898 23996 26908 24052
rect 26964 23996 28364 24052
rect 28420 23996 31948 24052
rect 31892 23940 31948 23996
rect 20514 23884 20524 23940
rect 20580 23884 21532 23940
rect 21588 23884 21598 23940
rect 31892 23884 37660 23940
rect 37716 23884 37726 23940
rect 41200 23604 42000 23632
rect 25554 23548 25564 23604
rect 25620 23548 26236 23604
rect 26292 23548 26302 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 41200 23520 42000 23548
rect 21858 23436 21868 23492
rect 21924 23436 23212 23492
rect 23268 23436 23278 23492
rect 17938 23212 17948 23268
rect 18004 23212 19292 23268
rect 19348 23212 20188 23268
rect 20244 23212 20254 23268
rect 4274 23100 4284 23156
rect 4340 23100 11004 23156
rect 11060 23100 14476 23156
rect 14532 23100 14542 23156
rect 14802 23100 14812 23156
rect 14868 23100 15932 23156
rect 15988 23100 16492 23156
rect 16548 23100 16558 23156
rect 16818 23100 16828 23156
rect 16884 23100 17836 23156
rect 17892 23100 17902 23156
rect 23874 23100 23884 23156
rect 23940 23100 25676 23156
rect 25732 23100 25742 23156
rect 14018 22988 14028 23044
rect 14084 22988 15148 23044
rect 15204 22988 15214 23044
rect 0 22932 800 22960
rect 0 22876 1932 22932
rect 1988 22876 1998 22932
rect 0 22848 800 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 17490 22428 17500 22484
rect 17556 22428 18060 22484
rect 18116 22428 21756 22484
rect 21812 22428 24332 22484
rect 24388 22428 25340 22484
rect 25396 22428 25406 22484
rect 28242 22428 28252 22484
rect 28308 22428 31948 22484
rect 31892 22372 31948 22428
rect 14354 22316 14364 22372
rect 14420 22316 18508 22372
rect 18564 22316 21644 22372
rect 21700 22316 22428 22372
rect 22484 22316 23548 22372
rect 23604 22316 23614 22372
rect 31892 22316 37660 22372
rect 37716 22316 37726 22372
rect 41200 22260 42000 22288
rect 24882 22204 24892 22260
rect 24948 22204 26124 22260
rect 26180 22204 26190 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 41200 22176 42000 22204
rect 18172 22092 21980 22148
rect 22036 22092 23212 22148
rect 23268 22092 23278 22148
rect 18172 21924 18228 22092
rect 20738 21980 20748 22036
rect 20804 21980 21756 22036
rect 21812 21980 21822 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 17042 21868 17052 21924
rect 17108 21868 18172 21924
rect 18228 21868 18238 21924
rect 13122 21756 13132 21812
rect 13188 21756 14140 21812
rect 14196 21756 14206 21812
rect 24994 21756 25004 21812
rect 25060 21756 26124 21812
rect 26180 21756 26190 21812
rect 26002 21644 26012 21700
rect 26068 21644 28252 21700
rect 28308 21644 28318 21700
rect 4274 21532 4284 21588
rect 4340 21532 10556 21588
rect 10612 21532 14364 21588
rect 14420 21532 14430 21588
rect 19058 21532 19068 21588
rect 19124 21532 20860 21588
rect 20916 21532 20926 21588
rect 21522 21532 21532 21588
rect 21588 21532 25676 21588
rect 25732 21532 25742 21588
rect 14018 21420 14028 21476
rect 14084 21420 14924 21476
rect 14980 21420 15708 21476
rect 15764 21420 16604 21476
rect 16660 21420 17388 21476
rect 17444 21420 17454 21476
rect 17714 21420 17724 21476
rect 17780 21420 18620 21476
rect 18676 21420 18686 21476
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 0 20916 800 20944
rect 0 20860 1932 20916
rect 1988 20860 1998 20916
rect 12226 20860 12236 20916
rect 12292 20860 14140 20916
rect 14196 20860 14206 20916
rect 17490 20860 17500 20916
rect 17556 20860 23884 20916
rect 23940 20860 23950 20916
rect 0 20832 800 20860
rect 20066 20748 20076 20804
rect 20132 20748 20636 20804
rect 20692 20748 20702 20804
rect 18610 20636 18620 20692
rect 18676 20636 21420 20692
rect 21476 20636 21486 20692
rect 22530 20636 22540 20692
rect 22596 20636 22988 20692
rect 23044 20636 23054 20692
rect 4162 20524 4172 20580
rect 4228 20524 19180 20580
rect 19236 20524 19246 20580
rect 22642 20524 22652 20580
rect 22708 20524 24108 20580
rect 24164 20524 24174 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 20626 20300 20636 20356
rect 20692 20300 21532 20356
rect 21588 20300 21598 20356
rect 13682 20188 13692 20244
rect 13748 20188 14252 20244
rect 14308 20188 14318 20244
rect 18050 20188 18060 20244
rect 18116 20188 20300 20244
rect 20356 20188 20366 20244
rect 20514 20188 20524 20244
rect 20580 20188 21868 20244
rect 21924 20188 21934 20244
rect 23202 20188 23212 20244
rect 23268 20188 25900 20244
rect 25956 20188 27356 20244
rect 27412 20188 27422 20244
rect 18732 20132 18788 20188
rect 17714 20076 17724 20132
rect 17780 20076 18508 20132
rect 18564 20076 18574 20132
rect 18722 20076 18732 20132
rect 18788 20076 18798 20132
rect 19618 20076 19628 20132
rect 19684 20076 20412 20132
rect 20468 20076 20478 20132
rect 21186 20076 21196 20132
rect 21252 20076 21644 20132
rect 21700 20076 21710 20132
rect 16034 19964 16044 20020
rect 16100 19964 18396 20020
rect 18452 19964 22540 20020
rect 22596 19964 22988 20020
rect 23044 19964 23054 20020
rect 25890 19964 25900 20020
rect 25956 19964 26908 20020
rect 26964 19964 26974 20020
rect 27906 19964 27916 20020
rect 27972 19964 28588 20020
rect 28644 19964 37660 20020
rect 37716 19964 37726 20020
rect 20178 19740 20188 19796
rect 20244 19740 20412 19796
rect 20468 19740 22204 19796
rect 22260 19740 22270 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 41200 19488 42000 19516
rect 14130 19404 14140 19460
rect 14196 19404 16044 19460
rect 16100 19404 16110 19460
rect 23650 19404 23660 19460
rect 23716 19404 26012 19460
rect 26068 19404 28028 19460
rect 28084 19404 28094 19460
rect 4274 19180 4284 19236
rect 4340 19180 11452 19236
rect 11508 19180 11518 19236
rect 13906 19180 13916 19236
rect 13972 19180 15148 19236
rect 15092 19124 15148 19180
rect 15092 19068 15372 19124
rect 15428 19068 15438 19124
rect 16146 19068 16156 19124
rect 16212 19068 16222 19124
rect 16156 19012 16212 19068
rect 13682 18956 13692 19012
rect 13748 18956 16212 19012
rect 20066 18956 20076 19012
rect 20132 18956 21868 19012
rect 21924 18956 21934 19012
rect 29474 18956 29484 19012
rect 29540 18956 37884 19012
rect 37940 18956 37950 19012
rect 0 18900 800 18928
rect 41200 18900 42000 18928
rect 0 18844 1932 18900
rect 1988 18844 1998 18900
rect 29250 18844 29260 18900
rect 29316 18844 37660 18900
rect 37716 18844 37726 18900
rect 40002 18844 40012 18900
rect 40068 18844 42000 18900
rect 0 18816 800 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 41200 18816 42000 18844
rect 22194 18732 22204 18788
rect 22260 18732 22764 18788
rect 22820 18732 23548 18788
rect 23604 18732 23614 18788
rect 14690 18620 14700 18676
rect 14756 18620 15596 18676
rect 15652 18620 15662 18676
rect 19506 18620 19516 18676
rect 19572 18620 21700 18676
rect 21970 18620 21980 18676
rect 22036 18620 23100 18676
rect 23156 18620 25900 18676
rect 25956 18620 25966 18676
rect 21644 18564 21700 18620
rect 11442 18508 11452 18564
rect 11508 18508 14924 18564
rect 14980 18508 14990 18564
rect 15810 18508 15820 18564
rect 15876 18508 17164 18564
rect 17220 18508 18508 18564
rect 18564 18508 18574 18564
rect 19516 18508 19628 18564
rect 19684 18508 20300 18564
rect 20356 18508 21420 18564
rect 21476 18508 21486 18564
rect 21644 18508 23548 18564
rect 23604 18508 23614 18564
rect 19516 18452 19572 18508
rect 4274 18396 4284 18452
rect 4340 18396 10892 18452
rect 10948 18396 14700 18452
rect 14756 18396 14766 18452
rect 16258 18396 16268 18452
rect 16324 18396 17388 18452
rect 17444 18396 17454 18452
rect 18162 18396 18172 18452
rect 18228 18396 19572 18452
rect 20738 18396 20748 18452
rect 20804 18396 21644 18452
rect 21700 18396 22092 18452
rect 22148 18396 23324 18452
rect 23380 18396 23390 18452
rect 23762 18396 23772 18452
rect 23828 18396 24332 18452
rect 24388 18396 25452 18452
rect 25508 18396 25518 18452
rect 25778 18396 25788 18452
rect 25844 18396 27244 18452
rect 27300 18396 27310 18452
rect 16706 18284 16716 18340
rect 16772 18284 19292 18340
rect 19348 18284 19358 18340
rect 19954 18284 19964 18340
rect 20020 18284 20524 18340
rect 20580 18284 20590 18340
rect 21196 18284 22428 18340
rect 22484 18284 22988 18340
rect 23044 18284 23054 18340
rect 24658 18284 24668 18340
rect 24724 18284 25340 18340
rect 25396 18284 26460 18340
rect 26516 18284 26526 18340
rect 0 18228 800 18256
rect 0 18172 1932 18228
rect 1988 18172 1998 18228
rect 0 18144 800 18172
rect 19292 18116 19348 18284
rect 21196 18228 21252 18284
rect 41200 18228 42000 18256
rect 21186 18172 21196 18228
rect 21252 18172 21262 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 41200 18144 42000 18172
rect 19292 18060 23996 18116
rect 24052 18060 24062 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 14018 17948 14028 18004
rect 14084 17948 14476 18004
rect 14532 17948 14542 18004
rect 23100 17892 23156 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 13794 17836 13804 17892
rect 13860 17836 14924 17892
rect 14980 17836 19516 17892
rect 19572 17836 19582 17892
rect 23090 17836 23100 17892
rect 23156 17836 23166 17892
rect 25666 17836 25676 17892
rect 25732 17836 27020 17892
rect 27076 17836 27086 17892
rect 16716 17724 21196 17780
rect 21252 17724 21262 17780
rect 16716 17668 16772 17724
rect 15362 17612 15372 17668
rect 15428 17612 16716 17668
rect 16772 17612 16782 17668
rect 18498 17612 18508 17668
rect 18564 17612 21532 17668
rect 21588 17612 21598 17668
rect 17378 17500 17388 17556
rect 17444 17500 19292 17556
rect 19348 17500 20188 17556
rect 20244 17500 21084 17556
rect 21140 17500 21150 17556
rect 27234 17500 27244 17556
rect 27300 17500 29372 17556
rect 29428 17500 29438 17556
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 14690 17052 14700 17108
rect 14756 17052 16044 17108
rect 16100 17052 17724 17108
rect 17780 17052 18844 17108
rect 18900 17052 20076 17108
rect 20132 17052 20142 17108
rect 22642 17052 22652 17108
rect 22708 17052 25228 17108
rect 25284 17052 25294 17108
rect 25330 16940 25340 16996
rect 25396 16940 26236 16996
rect 26292 16940 37660 16996
rect 37716 16940 37726 16996
rect 41200 16884 42000 16912
rect 17266 16828 17276 16884
rect 17332 16828 17948 16884
rect 18004 16828 21756 16884
rect 21812 16828 23996 16884
rect 24052 16828 24062 16884
rect 24658 16828 24668 16884
rect 24724 16828 25564 16884
rect 25620 16828 25630 16884
rect 40002 16828 40012 16884
rect 40068 16828 42000 16884
rect 41200 16800 42000 16828
rect 16818 16716 16828 16772
rect 16884 16716 17836 16772
rect 17892 16716 18284 16772
rect 18340 16716 18350 16772
rect 20850 16716 20860 16772
rect 20916 16716 22540 16772
rect 22596 16716 22606 16772
rect 22866 16716 22876 16772
rect 22932 16716 26684 16772
rect 26740 16716 26750 16772
rect 21970 16604 21980 16660
rect 22036 16604 22764 16660
rect 22820 16604 22830 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 20738 16156 20748 16212
rect 20804 16156 21420 16212
rect 21476 16156 22484 16212
rect 22428 16100 22484 16156
rect 18610 16044 18620 16100
rect 18676 16044 19852 16100
rect 19908 16044 21532 16100
rect 21588 16044 21598 16100
rect 22418 16044 22428 16100
rect 22484 16044 22494 16100
rect 26114 16044 26124 16100
rect 26180 16044 26796 16100
rect 26852 16044 26862 16100
rect 20290 15932 20300 15988
rect 20356 15932 21644 15988
rect 21700 15932 21710 15988
rect 18722 15820 18732 15876
rect 18788 15820 21308 15876
rect 21364 15820 23324 15876
rect 23380 15820 23390 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 21410 15596 21420 15652
rect 21476 15596 21868 15652
rect 21924 15596 21934 15652
rect 41200 15540 42000 15568
rect 21634 15484 21644 15540
rect 21700 15484 21980 15540
rect 22036 15484 22046 15540
rect 40002 15484 40012 15540
rect 40068 15484 42000 15540
rect 41200 15456 42000 15484
rect 27906 15148 27916 15204
rect 27972 15148 29260 15204
rect 29316 15148 37660 15204
rect 37716 15148 37726 15204
rect 21074 15036 21084 15092
rect 21140 15036 21868 15092
rect 21924 15036 21934 15092
rect 20178 14924 20188 14980
rect 20244 14924 22092 14980
rect 22148 14924 22158 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 24546 14812 24556 14868
rect 24612 14812 24622 14868
rect 24556 14756 24612 14812
rect 17154 14700 17164 14756
rect 17220 14700 18060 14756
rect 18116 14700 24612 14756
rect 21522 14588 21532 14644
rect 21588 14588 21598 14644
rect 22082 14588 22092 14644
rect 22148 14588 26124 14644
rect 26180 14588 26190 14644
rect 16482 14476 16492 14532
rect 16548 14476 17276 14532
rect 17332 14476 17342 14532
rect 17602 14476 17612 14532
rect 17668 14476 18508 14532
rect 18564 14476 18574 14532
rect 21532 14420 21588 14588
rect 21858 14476 21868 14532
rect 21924 14476 22764 14532
rect 22820 14476 22830 14532
rect 26226 14476 26236 14532
rect 26292 14476 27020 14532
rect 27076 14476 27086 14532
rect 31892 14476 37660 14532
rect 37716 14476 37726 14532
rect 21532 14364 26908 14420
rect 26964 14364 27580 14420
rect 27636 14364 27646 14420
rect 31892 14308 31948 14476
rect 14690 14252 14700 14308
rect 14756 14252 16380 14308
rect 16436 14252 16446 14308
rect 27234 14252 27244 14308
rect 27300 14252 28252 14308
rect 28308 14252 31948 14308
rect 41200 14196 42000 14224
rect 40002 14140 40012 14196
rect 40068 14140 42000 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 41200 14112 42000 14140
rect 14018 13916 14028 13972
rect 14084 13916 16940 13972
rect 16996 13916 17500 13972
rect 17556 13916 20300 13972
rect 20356 13916 21308 13972
rect 21364 13916 23436 13972
rect 23492 13916 24668 13972
rect 24724 13916 26012 13972
rect 26068 13916 26078 13972
rect 22530 13692 22540 13748
rect 22596 13692 23436 13748
rect 23492 13692 23502 13748
rect 23762 13692 23772 13748
rect 23828 13692 24332 13748
rect 24388 13692 24398 13748
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 17490 3612 17500 3668
rect 17556 3612 18620 3668
rect 18676 3612 18686 3668
rect 23762 3612 23772 3668
rect 23828 3612 25564 3668
rect 25620 3612 25630 3668
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 23436 27916 23492 27972
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 23436 26124 23492 26180
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 23436 27972 23492 27982
rect 23436 26180 23492 27916
rect 23436 26114 23492 26124
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18368 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18256 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _107_
timestamp 1698175906
transform -1 0 15904 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_
timestamp 1698175906
transform 1 0 17696 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20160 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1698175906
transform -1 0 16688 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _111_
timestamp 1698175906
transform -1 0 18928 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1698175906
transform -1 0 16240 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20720 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1698175906
transform 1 0 21952 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14560 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13552 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698175906
transform -1 0 21840 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _119_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19264 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698175906
transform -1 0 17920 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15120 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _122_
timestamp 1698175906
transform -1 0 14560 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _123_
timestamp 1698175906
transform 1 0 18256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1698175906
transform 1 0 19936 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _126_
timestamp 1698175906
transform -1 0 20944 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20272 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698175906
transform -1 0 22176 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _129_
timestamp 1698175906
transform -1 0 22288 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _130_
timestamp 1698175906
transform -1 0 21728 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform 1 0 18368 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform -1 0 19824 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _133_
timestamp 1698175906
transform -1 0 16464 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _134_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14672 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _135_
timestamp 1698175906
transform 1 0 12096 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _136_
timestamp 1698175906
transform 1 0 21280 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _137_
timestamp 1698175906
transform 1 0 22064 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _138_
timestamp 1698175906
transform 1 0 22624 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _139_
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _140_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18928 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _141_
timestamp 1698175906
transform -1 0 18368 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _142_
timestamp 1698175906
transform -1 0 22064 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _143_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20720 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _144_
timestamp 1698175906
transform 1 0 16352 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform 1 0 17696 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _146_
timestamp 1698175906
transform -1 0 17024 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _147_
timestamp 1698175906
transform 1 0 15232 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _148_
timestamp 1698175906
transform 1 0 14672 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _149_
timestamp 1698175906
transform -1 0 23520 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _150_
timestamp 1698175906
transform 1 0 20048 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _151_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _152_
timestamp 1698175906
transform -1 0 15232 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _153_
timestamp 1698175906
transform -1 0 14224 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _154_
timestamp 1698175906
transform 1 0 21616 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _155_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16352 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _156_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18032 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _157_
timestamp 1698175906
transform -1 0 16688 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698175906
transform -1 0 19824 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _159_
timestamp 1698175906
transform -1 0 19264 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _160_
timestamp 1698175906
transform -1 0 20272 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _161_
timestamp 1698175906
transform 1 0 23296 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _162_
timestamp 1698175906
transform 1 0 21840 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _163_
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _164_
timestamp 1698175906
transform -1 0 24752 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _165_
timestamp 1698175906
transform 1 0 23744 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _166_
timestamp 1698175906
transform 1 0 23184 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _167_
timestamp 1698175906
transform -1 0 26432 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _168_
timestamp 1698175906
transform -1 0 25200 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _169_
timestamp 1698175906
transform -1 0 24416 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _170_
timestamp 1698175906
transform 1 0 22512 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _171_
timestamp 1698175906
transform -1 0 21504 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _172_
timestamp 1698175906
transform 1 0 27440 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _173_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22960 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _174_
timestamp 1698175906
transform 1 0 25872 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _175_
timestamp 1698175906
transform -1 0 22288 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _176_
timestamp 1698175906
transform 1 0 22400 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _177_
timestamp 1698175906
transform 1 0 26544 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _178_
timestamp 1698175906
transform 1 0 26768 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _179_
timestamp 1698175906
transform 1 0 18368 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _180_
timestamp 1698175906
transform -1 0 20608 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _181_
timestamp 1698175906
transform 1 0 19712 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _182_
timestamp 1698175906
transform 1 0 25872 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _183_
timestamp 1698175906
transform -1 0 19712 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _184_
timestamp 1698175906
transform -1 0 18816 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _185_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20384 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _186_
timestamp 1698175906
transform -1 0 23968 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _187_
timestamp 1698175906
transform 1 0 21728 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _188_
timestamp 1698175906
transform 1 0 22288 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _189_
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _190_
timestamp 1698175906
transform 1 0 22624 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _191_
timestamp 1698175906
transform -1 0 22288 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _192_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22848 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _193_
timestamp 1698175906
transform 1 0 27440 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _194_
timestamp 1698175906
transform 1 0 26544 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _195_
timestamp 1698175906
transform -1 0 15120 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _196_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _197_
timestamp 1698175906
transform -1 0 27552 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _198_
timestamp 1698175906
transform 1 0 25312 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _199_
timestamp 1698175906
transform 1 0 16352 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _200_
timestamp 1698175906
transform -1 0 16128 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _201_
timestamp 1698175906
transform 1 0 22176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _202_
timestamp 1698175906
transform 1 0 21952 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _203_
timestamp 1698175906
transform -1 0 25648 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _204_
timestamp 1698175906
transform 1 0 23184 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _205_
timestamp 1698175906
transform 1 0 23408 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _206_
timestamp 1698175906
transform 1 0 26432 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _207_
timestamp 1698175906
transform 1 0 25536 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _208_
timestamp 1698175906
transform -1 0 25648 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _209_
timestamp 1698175906
transform 1 0 22960 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14560 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform -1 0 14112 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 19824 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform -1 0 13664 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 13776 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 16688 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 17248 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 14000 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform -1 0 14560 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 13776 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 17136 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 23184 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 25200 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 21728 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 26208 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 25200 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 25536 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform -1 0 14000 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 26320 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 13776 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform 1 0 22848 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 25312 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform 1 0 22624 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _237_
timestamp 1698175906
transform -1 0 14896 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _238_
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _239_
timestamp 1698175906
transform -1 0 13104 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__156__A2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18032 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__A2
timestamp 1698175906
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__A2
timestamp 1698175906
transform -1 0 24416 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__A2
timestamp 1698175906
transform -1 0 17808 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 14672 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 14336 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 24304 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 13664 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 17024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform -1 0 20384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 20496 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 15456 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 20608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 26432 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 24304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 21504 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 25984 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 20720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform -1 0 24864 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 23408 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 25312 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 14224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 18032 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 22624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 22400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 19264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform -1 0 24416 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698175906
transform 1 0 18144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_154
timestamp 1698175906
transform 1 0 18592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_156
timestamp 1698175906
transform 1 0 18816 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_161
timestamp 1698175906
transform 1 0 19376 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_193 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22960 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_123
timestamp 1698175906
transform 1 0 15120 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_131
timestamp 1698175906
transform 1 0 16016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_135
timestamp 1698175906
transform 1 0 16464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_166
timestamp 1698175906
transform 1 0 19936 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_170
timestamp 1698175906
transform 1 0 20384 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_206
timestamp 1698175906
transform 1 0 24416 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_210
timestamp 1698175906
transform 1 0 24864 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_242
timestamp 1698175906
transform 1 0 28448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698175906
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_104
timestamp 1698175906
transform 1 0 12992 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_108
timestamp 1698175906
transform 1 0 13440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_110
timestamp 1698175906
transform 1 0 13664 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_152
timestamp 1698175906
transform 1 0 18368 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_202
timestamp 1698175906
transform 1 0 23968 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_206
timestamp 1698175906
transform 1 0 24416 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_242
timestamp 1698175906
transform 1 0 28448 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_274
timestamp 1698175906
transform 1 0 32032 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_278
timestamp 1698175906
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_131
timestamp 1698175906
transform 1 0 16016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_137
timestamp 1698175906
transform 1 0 16688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_139
timestamp 1698175906
transform 1 0 16912 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_157
timestamp 1698175906
transform 1 0 18928 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698175906
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_181
timestamp 1698175906
transform 1 0 21616 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_195
timestamp 1698175906
transform 1 0 23184 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_199
timestamp 1698175906
transform 1 0 23632 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_215
timestamp 1698175906
transform 1 0 25424 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_239
timestamp 1698175906
transform 1 0 28112 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698175906
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_321
timestamp 1698175906
transform 1 0 37296 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_146
timestamp 1698175906
transform 1 0 17696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_148
timestamp 1698175906
transform 1 0 17920 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_151
timestamp 1698175906
transform 1 0 18256 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_167
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_169
timestamp 1698175906
transform 1 0 20272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_187
timestamp 1698175906
transform 1 0 22288 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_203
timestamp 1698175906
transform 1 0 24080 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698175906
transform 1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_251
timestamp 1698175906
transform 1 0 29456 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_267
timestamp 1698175906
transform 1 0 31248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_275
timestamp 1698175906
transform 1 0 32144 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_139
timestamp 1698175906
transform 1 0 16912 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_142
timestamp 1698175906
transform 1 0 17248 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_158
timestamp 1698175906
transform 1 0 19040 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_162
timestamp 1698175906
transform 1 0 19488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698175906
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_192
timestamp 1698175906
transform 1 0 22848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_194
timestamp 1698175906
transform 1 0 23072 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_224
timestamp 1698175906
transform 1 0 26432 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_233
timestamp 1698175906
transform 1 0 27440 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698175906
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 37296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_104
timestamp 1698175906
transform 1 0 12992 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_108
timestamp 1698175906
transform 1 0 13440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_110
timestamp 1698175906
transform 1 0 13664 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_148
timestamp 1698175906
transform 1 0 17920 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_150
timestamp 1698175906
transform 1 0 18144 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_155
timestamp 1698175906
transform 1 0 18704 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_163
timestamp 1698175906
transform 1 0 19600 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_180
timestamp 1698175906
transform 1 0 21504 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_187
timestamp 1698175906
transform 1 0 22288 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_197
timestamp 1698175906
transform 1 0 23408 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_217
timestamp 1698175906
transform 1 0 25648 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_221
timestamp 1698175906
transform 1 0 26096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_223
timestamp 1698175906
transform 1 0 26320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_226
timestamp 1698175906
transform 1 0 26656 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_258
timestamp 1698175906
transform 1 0 30240 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_274
timestamp 1698175906
transform 1 0 32032 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698175906
transform 1 0 32480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_123
timestamp 1698175906
transform 1 0 15120 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_131
timestamp 1698175906
transform 1 0 16016 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_133
timestamp 1698175906
transform 1 0 16240 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_144
timestamp 1698175906
transform 1 0 17472 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_158
timestamp 1698175906
transform 1 0 19040 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_165
timestamp 1698175906
transform 1 0 19824 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698175906
transform 1 0 20608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_227
timestamp 1698175906
transform 1 0 26768 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_234
timestamp 1698175906
transform 1 0 27552 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_242
timestamp 1698175906
transform 1 0 28448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 4480 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 8064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_88
timestamp 1698175906
transform 1 0 11200 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_126
timestamp 1698175906
transform 1 0 15456 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_135
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_150
timestamp 1698175906
transform 1 0 18144 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_157
timestamp 1698175906
transform 1 0 18928 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_201
timestamp 1698175906
transform 1 0 23856 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_205
timestamp 1698175906
transform 1 0 24304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_207
timestamp 1698175906
transform 1 0 24528 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_252
timestamp 1698175906
transform 1 0 29568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_268
timestamp 1698175906
transform 1 0 31360 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698175906
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698175906
transform 1 0 4928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_117
timestamp 1698175906
transform 1 0 14448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_121
timestamp 1698175906
transform 1 0 14896 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_123
timestamp 1698175906
transform 1 0 15120 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_130
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_137
timestamp 1698175906
transform 1 0 16688 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_153
timestamp 1698175906
transform 1 0 18480 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_161
timestamp 1698175906
transform 1 0 19376 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_165
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698175906
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_201
timestamp 1698175906
transform 1 0 23856 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_209
timestamp 1698175906
transform 1 0 24752 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_213
timestamp 1698175906
transform 1 0 25200 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_253
timestamp 1698175906
transform 1 0 29680 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_285
timestamp 1698175906
transform 1 0 33264 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_301
timestamp 1698175906
transform 1 0 35056 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_309
timestamp 1698175906
transform 1 0 35952 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_313
timestamp 1698175906
transform 1 0 36400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_80
timestamp 1698175906
transform 1 0 10304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_113
timestamp 1698175906
transform 1 0 14000 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_117
timestamp 1698175906
transform 1 0 14448 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_125
timestamp 1698175906
transform 1 0 15344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_133
timestamp 1698175906
transform 1 0 16240 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_137
timestamp 1698175906
transform 1 0 16688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_144
timestamp 1698175906
transform 1 0 17472 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_157
timestamp 1698175906
transform 1 0 18928 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_165
timestamp 1698175906
transform 1 0 19824 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_189
timestamp 1698175906
transform 1 0 22512 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_191
timestamp 1698175906
transform 1 0 22736 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_205
timestamp 1698175906
transform 1 0 24304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_216
timestamp 1698175906
transform 1 0 25536 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_218
timestamp 1698175906
transform 1 0 25760 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_241
timestamp 1698175906
transform 1 0 28336 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_273
timestamp 1698175906
transform 1 0 31920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698175906
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_69
timestamp 1698175906
transform 1 0 9072 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_85
timestamp 1698175906
transform 1 0 10864 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_93
timestamp 1698175906
transform 1 0 11760 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_95
timestamp 1698175906
transform 1 0 11984 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_100
timestamp 1698175906
transform 1 0 12544 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698175906
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_119
timestamp 1698175906
transform 1 0 14672 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_151
timestamp 1698175906
transform 1 0 18256 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_155
timestamp 1698175906
transform 1 0 18704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_157
timestamp 1698175906
transform 1 0 18928 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_160
timestamp 1698175906
transform 1 0 19264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_162
timestamp 1698175906
transform 1 0 19488 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_198
timestamp 1698175906
transform 1 0 23520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_206
timestamp 1698175906
transform 1 0 24416 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_238
timestamp 1698175906
transform 1 0 28000 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1698175906
transform 1 0 28448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 4480 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 8064 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_80
timestamp 1698175906
transform 1 0 10304 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_123
timestamp 1698175906
transform 1 0 15120 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_132
timestamp 1698175906
transform 1 0 16128 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_224
timestamp 1698175906
transform 1 0 26432 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_256
timestamp 1698175906
transform 1 0 30016 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_272
timestamp 1698175906
transform 1 0 31808 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 40096 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 40320 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_109
timestamp 1698175906
transform 1 0 13552 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_112
timestamp 1698175906
transform 1 0 13888 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_202
timestamp 1698175906
transform 1 0 23968 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_204
timestamp 1698175906
transform 1 0 24192 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_242
timestamp 1698175906
transform 1 0 28448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 4480 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_80
timestamp 1698175906
transform 1 0 10304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_84
timestamp 1698175906
transform 1 0 10752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_114
timestamp 1698175906
transform 1 0 14112 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_118
timestamp 1698175906
transform 1 0 14560 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_127
timestamp 1698175906
transform 1 0 15568 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_131
timestamp 1698175906
transform 1 0 16016 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_133
timestamp 1698175906
transform 1 0 16240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_151
timestamp 1698175906
transform 1 0 18256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_155
timestamp 1698175906
transform 1 0 18704 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_206
timestamp 1698175906
transform 1 0 24416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_229
timestamp 1698175906
transform 1 0 26992 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_261
timestamp 1698175906
transform 1 0 30576 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 40320 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_173
timestamp 1698175906
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_179
timestamp 1698175906
transform 1 0 21392 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_211
timestamp 1698175906
transform 1 0 24976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_213
timestamp 1698175906
transform 1 0 25200 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_88
timestamp 1698175906
transform 1 0 11200 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_124
timestamp 1698175906
transform 1 0 15232 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_128
timestamp 1698175906
transform 1 0 15680 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698175906
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_174
timestamp 1698175906
transform 1 0 20832 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_178
timestamp 1698175906
transform 1 0 21280 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_180
timestamp 1698175906
transform 1 0 21504 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_189
timestamp 1698175906
transform 1 0 22512 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_193
timestamp 1698175906
transform 1 0 22960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_206
timestamp 1698175906
transform 1 0 24416 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 36512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 37408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_69
timestamp 1698175906
transform 1 0 9072 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_85
timestamp 1698175906
transform 1 0 10864 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_93
timestamp 1698175906
transform 1 0 11760 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_97
timestamp 1698175906
transform 1 0 12208 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_121
timestamp 1698175906
transform 1 0 14896 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_125
timestamp 1698175906
transform 1 0 15344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_127
timestamp 1698175906
transform 1 0 15568 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_132
timestamp 1698175906
transform 1 0 16128 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_143
timestamp 1698175906
transform 1 0 17360 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_147
timestamp 1698175906
transform 1 0 17808 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_156
timestamp 1698175906
transform 1 0 18816 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_158
timestamp 1698175906
transform 1 0 19040 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_164
timestamp 1698175906
transform 1 0 19712 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698175906
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_179
timestamp 1698175906
transform 1 0 21392 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_190
timestamp 1698175906
transform 1 0 22624 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_222
timestamp 1698175906
transform 1 0 26208 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_238
timestamp 1698175906
transform 1 0 28000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698175906
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 4480 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_104
timestamp 1698175906
transform 1 0 12992 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_108
timestamp 1698175906
transform 1 0 13440 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_110
timestamp 1698175906
transform 1 0 13664 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_171
timestamp 1698175906
transform 1 0 20496 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_175
timestamp 1698175906
transform 1 0 20944 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_183
timestamp 1698175906
transform 1 0 21840 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_189
timestamp 1698175906
transform 1 0 22512 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_201
timestamp 1698175906
transform 1 0 23856 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_217
timestamp 1698175906
transform 1 0 25648 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_249
timestamp 1698175906
transform 1 0 29232 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_265
timestamp 1698175906
transform 1 0 31024 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_273
timestamp 1698175906
transform 1 0 31920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 32368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_139
timestamp 1698175906
transform 1 0 16912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_170
timestamp 1698175906
transform 1 0 20384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698175906
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_187
timestamp 1698175906
transform 1 0 22288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_189
timestamp 1698175906
transform 1 0 22512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_221
timestamp 1698175906
transform 1 0 26096 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_237
timestamp 1698175906
transform 1 0 27888 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_150
timestamp 1698175906
transform 1 0 18144 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_154
timestamp 1698175906
transform 1 0 18592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_194
timestamp 1698175906
transform 1 0 23072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_203
timestamp 1698175906
transform 1 0 24080 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698175906
transform 1 0 24528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_217
timestamp 1698175906
transform 1 0 25648 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_249
timestamp 1698175906
transform 1 0 29232 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_265
timestamp 1698175906
transform 1 0 31024 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_273
timestamp 1698175906
transform 1 0 31920 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_277
timestamp 1698175906
transform 1 0 32368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_279
timestamp 1698175906
transform 1 0 32592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_185
timestamp 1698175906
transform 1 0 22064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_187
timestamp 1698175906
transform 1 0 22288 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_219
timestamp 1698175906
transform 1 0 25872 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_235
timestamp 1698175906
transform 1 0 27664 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_243
timestamp 1698175906
transform 1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_168
timestamp 1698175906
transform 1 0 20160 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_195
timestamp 1698175906
transform 1 0 23184 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698175906
transform 1 0 24080 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 25536 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_243
timestamp 1698175906
transform 1 0 28560 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698175906
transform 1 0 32144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_206
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_210
timestamp 1698175906
transform 1 0 24864 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_237
timestamp 1698175906
transform 1 0 27888 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita63_26 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37520 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 24976 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 37520 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 20384 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 37520 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform -1 0 24192 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 25648 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 37520 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 4480 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 20272 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform -1 0 4480 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 4480 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 24192 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 4480 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform -1 0 4480 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 17472 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 41200 15456 42000 15568 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 24864 41200 24976 42000 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 41200 14112 42000 14224 0 FreeSans 448 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 19488 41200 19600 42000 0 FreeSans 448 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 41200 18816 42000 18928 0 FreeSans 448 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 16800 41200 16912 42000 0 FreeSans 448 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 25536 41200 25648 42000 0 FreeSans 448 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 41200 24192 42000 24304 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 41200 16800 42000 16912 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 20160 41200 20272 42000 0 FreeSans 448 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 13552 18536 13552 18536 0 _000_
rlabel metal3 13664 21784 13664 21784 0 _001_
rlabel metal2 21224 27384 21224 27384 0 _002_
rlabel metal2 12376 21224 12376 21224 0 _003_
rlabel metal2 18872 17248 18872 17248 0 _004_
rlabel metal2 17640 13440 17640 13440 0 _005_
rlabel metal2 18200 22792 18200 22792 0 _006_
rlabel metal2 14952 22736 14952 22736 0 _007_
rlabel metal2 13608 25200 13608 25200 0 _008_
rlabel metal2 14728 14056 14728 14056 0 _009_
rlabel metal2 18088 27384 18088 27384 0 _010_
rlabel metal2 24248 16184 24248 16184 0 _011_
rlabel metal3 25536 22232 25536 22232 0 _012_
rlabel metal2 22736 22456 22736 22456 0 _013_
rlabel metal2 27216 15400 27216 15400 0 _014_
rlabel metal2 26152 14056 26152 14056 0 _015_
rlabel metal2 18312 25816 18312 25816 0 _016_
rlabel metal2 22064 13048 22064 13048 0 _017_
rlabel metal2 21112 14112 21112 14112 0 _018_
rlabel metal2 26656 19320 26656 19320 0 _019_
rlabel metal2 13048 18816 13048 18816 0 _020_
rlabel metal3 26544 18424 26544 18424 0 _021_
rlabel metal2 15848 25928 15848 25928 0 _022_
rlabel metal2 23800 27384 23800 27384 0 _023_
rlabel metal2 25816 23576 25816 23576 0 _024_
rlabel metal3 23352 26152 23352 26152 0 _025_
rlabel metal2 14728 24808 14728 24808 0 _026_
rlabel metal2 24472 13944 24472 13944 0 _027_
rlabel metal2 17752 14812 17752 14812 0 _028_
rlabel metal2 17304 14560 17304 14560 0 _029_
rlabel metal2 19208 27832 19208 27832 0 _030_
rlabel metal2 19656 20552 19656 20552 0 _031_
rlabel metal3 24640 18424 24640 18424 0 _032_
rlabel metal2 22680 16968 22680 16968 0 _033_
rlabel metal3 25144 16856 25144 16856 0 _034_
rlabel metal2 24248 21168 24248 21168 0 _035_
rlabel metal2 25480 27552 25480 27552 0 _036_
rlabel metal3 25592 21784 25592 21784 0 _037_
rlabel metal2 23352 23408 23352 23408 0 _038_
rlabel metal3 24248 14392 24248 14392 0 _039_
rlabel metal2 27720 15400 27720 15400 0 _040_
rlabel metal2 28056 19712 28056 19712 0 _041_
rlabel metal2 26656 14728 26656 14728 0 _042_
rlabel metal3 22400 16632 22400 16632 0 _043_
rlabel metal2 26712 16408 26712 16408 0 _044_
rlabel metal3 26656 14504 26656 14504 0 _045_
rlabel metal3 19264 16072 19264 16072 0 _046_
rlabel metal2 20328 16296 20328 16296 0 _047_
rlabel metal2 22120 14728 22120 14728 0 _048_
rlabel metal2 18928 25368 18928 25368 0 _049_
rlabel metal2 21896 14784 21896 14784 0 _050_
rlabel metal3 23016 13720 23016 13720 0 _051_
rlabel metal2 22120 16184 22120 16184 0 _052_
rlabel metal2 21896 15568 21896 15568 0 _053_
rlabel metal2 22904 14924 22904 14924 0 _054_
rlabel metal2 27384 20188 27384 20188 0 _055_
rlabel metal2 27720 20132 27720 20132 0 _056_
rlabel metal2 14560 17864 14560 17864 0 _057_
rlabel metal2 27048 17752 27048 17752 0 _058_
rlabel metal3 16408 25368 16408 25368 0 _059_
rlabel metal2 22400 27832 22400 27832 0 _060_
rlabel metal2 23072 26488 23072 26488 0 _061_
rlabel metal3 24584 26488 24584 26488 0 _062_
rlabel metal2 23912 22736 23912 22736 0 _063_
rlabel metal2 26544 22904 26544 22904 0 _064_
rlabel metal3 24472 26936 24472 26936 0 _065_
rlabel metal3 18760 20160 18760 20160 0 _066_
rlabel metal2 18536 19320 18536 19320 0 _067_
rlabel metal2 15176 23072 15176 23072 0 _068_
rlabel metal3 19600 18536 19600 18536 0 _069_
rlabel metal2 16632 19208 16632 19208 0 _070_
rlabel metal2 16184 19824 16184 19824 0 _071_
rlabel metal2 18424 20048 18424 20048 0 _072_
rlabel metal2 15680 20104 15680 20104 0 _073_
rlabel metal3 21448 18424 21448 18424 0 _074_
rlabel metal3 16072 17640 16072 17640 0 _075_
rlabel metal2 14840 18928 14840 18928 0 _076_
rlabel metal2 21168 18424 21168 18424 0 _077_
rlabel metal2 18536 23800 18536 23800 0 _078_
rlabel metal2 21448 19936 21448 19936 0 _079_
rlabel metal2 15736 21504 15736 21504 0 _080_
rlabel metal2 14616 21616 14616 21616 0 _081_
rlabel metal2 22008 17360 22008 17360 0 _082_
rlabel metal2 22232 19544 22232 19544 0 _083_
rlabel metal2 22120 22848 22120 22848 0 _084_
rlabel metal2 20664 21392 20664 21392 0 _085_
rlabel metal2 21952 24696 21952 24696 0 _086_
rlabel metal2 19656 27356 19656 27356 0 _087_
rlabel metal2 21672 26936 21672 26936 0 _088_
rlabel metal2 17416 17584 17416 17584 0 _089_
rlabel metal2 16184 18536 16184 18536 0 _090_
rlabel metal3 13216 20888 13216 20888 0 _091_
rlabel metal2 25928 19320 25928 19320 0 _092_
rlabel metal2 22792 18648 22792 18648 0 _093_
rlabel metal3 20048 15848 20048 15848 0 _094_
rlabel metal2 17584 14504 17584 14504 0 _095_
rlabel metal2 18200 14056 18200 14056 0 _096_
rlabel metal2 21560 20720 21560 20720 0 _097_
rlabel metal2 18928 27944 18928 27944 0 _098_
rlabel metal3 17360 23128 17360 23128 0 _099_
rlabel metal2 23688 22848 23688 22848 0 _100_
rlabel metal2 15456 21784 15456 21784 0 _101_
rlabel metal2 22344 20720 22344 20720 0 _102_
rlabel metal2 20552 20048 20552 20048 0 _103_
rlabel metal2 22288 25368 22288 25368 0 _104_
rlabel metal3 2478 27608 2478 27608 0 clk
rlabel metal2 23016 22400 23016 22400 0 clknet_0_clk
rlabel metal2 20328 13384 20328 13384 0 clknet_1_0__leaf_clk
rlabel metal2 23128 27384 23128 27384 0 clknet_1_1__leaf_clk
rlabel metal2 18424 16800 18424 16800 0 dut63.count\[0\]
rlabel metal2 19712 13048 19712 13048 0 dut63.count\[1\]
rlabel metal2 20832 22232 20832 22232 0 dut63.count\[2\]
rlabel metal2 18200 21784 18200 21784 0 dut63.count\[3\]
rlabel metal2 27944 14840 27944 14840 0 net1
rlabel metal2 24584 5964 24584 5964 0 net10
rlabel metal2 23408 3528 23408 3528 0 net11
rlabel metal2 17136 31920 17136 31920 0 net12
rlabel metal2 25648 27160 25648 27160 0 net13
rlabel metal2 24808 24360 24808 24360 0 net14
rlabel metal2 28616 19656 28616 19656 0 net15
rlabel metal2 10920 19152 10920 19152 0 net16
rlabel metal2 28280 22064 28280 22064 0 net17
rlabel metal2 37688 17304 37688 17304 0 net18
rlabel metal2 20216 27608 20216 27608 0 net19
rlabel metal2 26936 23688 26936 23688 0 net2
rlabel metal2 12600 25816 12600 25816 0 net20
rlabel metal2 10584 21504 10584 21504 0 net21
rlabel metal2 22904 28112 22904 28112 0 net22
rlabel metal2 11480 18760 11480 18760 0 net23
rlabel metal2 11032 23072 11032 23072 0 net24
rlabel metal2 17976 5964 17976 5964 0 net25
rlabel metal2 18872 2590 18872 2590 0 net26
rlabel metal2 25368 28392 25368 28392 0 net3
rlabel metal2 28280 13944 28280 13944 0 net4
rlabel metal3 9352 27048 9352 27048 0 net5
rlabel metal2 19600 38024 19600 38024 0 net6
rlabel metal2 37912 18704 37912 18704 0 net7
rlabel metal2 11480 25032 11480 25032 0 net8
rlabel metal2 29288 19040 29288 19040 0 net9
rlabel metal2 40040 15848 40040 15848 0 segm[10]
rlabel metal2 40040 23800 40040 23800 0 segm[11]
rlabel metal2 24920 39746 24920 39746 0 segm[12]
rlabel metal2 40040 14392 40040 14392 0 segm[13]
rlabel metal3 1358 26264 1358 26264 0 segm[1]
rlabel metal2 19544 39746 19544 39746 0 segm[2]
rlabel metal3 40642 18200 40642 18200 0 segm[3]
rlabel metal3 1414 24920 1414 24920 0 segm[4]
rlabel metal2 40040 19096 40040 19096 0 segm[5]
rlabel metal2 23576 854 23576 854 0 segm[6]
rlabel metal2 22232 2086 22232 2086 0 segm[7]
rlabel metal2 16856 39354 16856 39354 0 segm[8]
rlabel metal2 25592 40194 25592 40194 0 segm[9]
rlabel metal2 40040 24360 40040 24360 0 sel[0]
rlabel metal2 40040 19656 40040 19656 0 sel[10]
rlabel metal3 1358 18200 1358 18200 0 sel[11]
rlabel metal2 40040 22344 40040 22344 0 sel[1]
rlabel metal2 40040 17304 40040 17304 0 sel[2]
rlabel metal2 20216 39354 20216 39354 0 sel[3]
rlabel metal3 1358 25592 1358 25592 0 sel[4]
rlabel metal3 1358 20888 1358 20888 0 sel[5]
rlabel metal2 22232 39690 22232 39690 0 sel[6]
rlabel metal3 1358 18872 1358 18872 0 sel[7]
rlabel metal3 1358 22904 1358 22904 0 sel[8]
rlabel metal2 17528 2198 17528 2198 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
