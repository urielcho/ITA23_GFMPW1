// This is the unpowered netlist.
module ita30 (clk,
    segm,
    sel);
 input clk;
 output [13:0] segm;
 output [11:0] sel;

 wire net24;
 wire net25;
 wire net26;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire \dut30.count[0] ;
 wire \dut30.count[1] ;
 wire \dut30.count[2] ;
 wire \dut30.count[3] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__217__A1 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__226__A2 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__228__A2 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__235__B2 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__236__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__237__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__239__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__240__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__241__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__242__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__243__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__244__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__245__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__246__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__248__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__249__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__250__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__251__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__252__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__253__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__255__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__256__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__257__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__259__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_139 ();
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _118_ (.I(\dut30.count[1] ),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _119_ (.I(_076_),
    .Z(_077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _120_ (.I(\dut30.count[3] ),
    .Z(_078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _121_ (.I(\dut30.count[2] ),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _122_ (.I(_079_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _123_ (.A1(_078_),
    .A2(_080_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _124_ (.A1(_077_),
    .A2(_081_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _125_ (.I(_082_),
    .Z(_083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _126_ (.A1(\dut30.count[0] ),
    .A2(_076_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _127_ (.I(_084_),
    .Z(_085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _128_ (.A1(_081_),
    .A2(_085_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _129_ (.I(net23),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _130_ (.I(\dut30.count[1] ),
    .Z(_088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _131_ (.I(\dut30.count[2] ),
    .Z(_089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _132_ (.I(_089_),
    .Z(_090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _133_ (.I(\dut30.count[3] ),
    .Z(_091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _134_ (.A1(_088_),
    .A2(_090_),
    .B(_091_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _135_ (.A1(_087_),
    .A2(_092_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _136_ (.A1(_086_),
    .A2(_093_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _137_ (.A1(_083_),
    .A2(_094_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _138_ (.I(\dut30.count[0] ),
    .Z(_095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _139_ (.I(_095_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _140_ (.I(\dut30.count[1] ),
    .Z(_096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _141_ (.A1(_000_),
    .A2(_096_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _142_ (.A1(_084_),
    .A2(_097_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _143_ (.I(\dut30.count[3] ),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _144_ (.A1(_098_),
    .A2(_090_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _145_ (.I(_079_),
    .Z(_100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _146_ (.A1(_095_),
    .A2(_096_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _147_ (.A1(_100_),
    .A2(_101_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _148_ (.I(_095_),
    .Z(_103_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _149_ (.A1(_103_),
    .A2(_096_),
    .A3(_089_),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _150_ (.A1(_102_),
    .A2(_104_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _151_ (.A1(_099_),
    .A2(_105_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _152_ (.A1(_091_),
    .A2(_104_),
    .Z(_106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _153_ (.I(_091_),
    .Z(_107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _154_ (.A1(_107_),
    .A2(_101_),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _155_ (.A1(_106_),
    .A2(_108_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _156_ (.I(_098_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _157_ (.A1(_109_),
    .A2(_080_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _158_ (.I(_110_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _159_ (.A1(net21),
    .A2(_111_),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _160_ (.A1(_106_),
    .A2(_112_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _161_ (.A1(_098_),
    .A2(_089_),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _162_ (.I(_110_),
    .Z(_114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _163_ (.A1(net19),
    .A2(_114_),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _164_ (.A1(_085_),
    .A2(_113_),
    .B(_115_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _165_ (.A1(_103_),
    .A2(_096_),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _166_ (.A1(_078_),
    .A2(_080_),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _167_ (.A1(_116_),
    .A2(_117_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _168_ (.A1(net18),
    .A2(_111_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _169_ (.A1(_025_),
    .A2(_026_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _170_ (.A1(_078_),
    .A2(_089_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _171_ (.A1(_103_),
    .A2(_088_),
    .A3(_027_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _172_ (.A1(net17),
    .A2(_111_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _173_ (.A1(_028_),
    .A2(_029_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _174_ (.I(_027_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _175_ (.A1(_095_),
    .A2(_077_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _176_ (.I(_031_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _177_ (.A1(net16),
    .A2(_114_),
    .B1(_030_),
    .B2(_032_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _178_ (.I(_033_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _179_ (.A1(_077_),
    .A2(_030_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _180_ (.A1(net15),
    .A2(_081_),
    .A3(_113_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _181_ (.I(_090_),
    .Z(_036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _182_ (.A1(_000_),
    .A2(_077_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _183_ (.I(_027_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _184_ (.I0(_113_),
    .I1(_038_),
    .S(_088_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _185_ (.A1(_036_),
    .A2(_037_),
    .B(_039_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _186_ (.A1(_034_),
    .A2(_035_),
    .B(_040_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _187_ (.A1(net12),
    .A2(_114_),
    .B1(_030_),
    .B2(_116_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _188_ (.I(_041_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _189_ (.A1(_001_),
    .A2(_117_),
    .B1(_027_),
    .B2(_031_),
    .C(_086_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _190_ (.A1(net9),
    .A2(_092_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _191_ (.I(_082_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _192_ (.A1(_092_),
    .A2(_042_),
    .B(_043_),
    .C(_044_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _193_ (.A1(_099_),
    .A2(_116_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _194_ (.A1(_090_),
    .A2(_085_),
    .B(_091_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _195_ (.A1(net10),
    .A2(_046_),
    .B1(_001_),
    .B2(_107_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _196_ (.A1(_045_),
    .A2(_047_),
    .B(_083_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _197_ (.A1(_088_),
    .A2(_036_),
    .B(_107_),
    .C(net11),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _198_ (.A1(_092_),
    .A2(_106_),
    .A3(_025_),
    .A4(_028_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _199_ (.A1(_048_),
    .A2(_049_),
    .B(_083_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _200_ (.A1(_031_),
    .A2(_117_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _201_ (.A1(net6),
    .A2(_111_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _202_ (.A1(_050_),
    .A2(_051_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _203_ (.I(net22),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _204_ (.A1(_052_),
    .A2(_045_),
    .B(_046_),
    .C(_044_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _205_ (.I(_103_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _206_ (.A1(_080_),
    .A2(_101_),
    .B(_109_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _207_ (.A1(net13),
    .A2(_054_),
    .B(_082_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _208_ (.A1(_053_),
    .A2(_083_),
    .B(_055_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _209_ (.A1(net14),
    .A2(_100_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _210_ (.A1(_100_),
    .A2(_101_),
    .B(_056_),
    .C(_109_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _211_ (.A1(_099_),
    .A2(_032_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _212_ (.A1(net7),
    .A2(_110_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _213_ (.A1(_025_),
    .A2(_028_),
    .A3(_057_),
    .A4(_058_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _214_ (.I(_054_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _215_ (.A1(_086_),
    .A2(_032_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _216_ (.A1(net8),
    .A2(_114_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _217_ (.A1(_059_),
    .A2(_060_),
    .B(_061_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _218_ (.A1(_085_),
    .A2(_117_),
    .B1(_030_),
    .B2(_032_),
    .C(_086_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _219_ (.I(net1),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _220_ (.A1(_053_),
    .A2(_082_),
    .B1(_054_),
    .B2(_063_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _221_ (.A1(_062_),
    .A2(_064_),
    .Z(_065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _222_ (.I(_065_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _223_ (.A1(_078_),
    .A2(_104_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _224_ (.A1(_099_),
    .A2(_116_),
    .B(_066_),
    .C(_054_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _225_ (.A1(_039_),
    .A2(_050_),
    .A3(_067_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _226_ (.A1(net2),
    .A2(_059_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _227_ (.A1(_053_),
    .A2(_044_),
    .B1(_068_),
    .B2(_069_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _228_ (.A1(net3),
    .A2(_059_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _229_ (.A1(_100_),
    .A2(_097_),
    .B(_109_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _230_ (.A1(_105_),
    .A2(_071_),
    .B(_067_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _231_ (.A1(_053_),
    .A2(_044_),
    .B1(_070_),
    .B2(_072_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _232_ (.A1(_039_),
    .A2(_050_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _233_ (.A1(_036_),
    .A2(_037_),
    .B(_107_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _234_ (.A1(net4),
    .A2(_036_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _235_ (.A1(_073_),
    .A2(_074_),
    .B1(_075_),
    .B2(_059_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _236_ (.D(_024_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _237_ (.D(_000_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\dut30.count[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _238_ (.D(_001_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\dut30.count[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _239_ (.D(_002_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\dut30.count[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _240_ (.D(_003_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\dut30.count[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _241_ (.D(_004_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _242_ (.D(_005_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _243_ (.D(_006_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _244_ (.D(_007_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net17));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _245_ (.D(_008_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net16));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _246_ (.D(_009_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net15));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _247_ (.D(_010_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net12));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _248_ (.D(_011_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net9));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _249_ (.D(_012_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net10));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _250_ (.D(_013_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net11));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _251_ (.D(_014_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net6));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _252_ (.D(_015_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _253_ (.D(_016_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net13));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _254_ (.D(_017_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net14));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _255_ (.D(_018_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net7));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _256_ (.D(_019_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net8));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _257_ (.D(_020_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _258_ (.D(_021_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net2));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _259_ (.D(_022_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net3));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _260_ (.D(_023_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _264_ (.I(net7),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _265_ (.I(net6),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita30_24 (.ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita30_25 (.ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__tiel ita30_26 (.ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output1 (.I(net1),
    .Z(segm[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output10 (.I(net10),
    .Z(segm[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output11 (.I(net11),
    .Z(segm[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output12 (.I(net12),
    .Z(sel[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output13 (.I(net13),
    .Z(sel[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output14 (.I(net14),
    .Z(sel[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output15 (.I(net15),
    .Z(sel[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output16 (.I(net16),
    .Z(sel[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output17 (.I(net17),
    .Z(sel[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output18 (.I(net18),
    .Z(sel[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output19 (.I(net19),
    .Z(sel[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output2 (.I(net2),
    .Z(segm[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output20 (.I(net20),
    .Z(sel[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output21 (.I(net21),
    .Z(sel[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output22 (.I(net22),
    .Z(sel[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output23 (.I(net23),
    .Z(sel[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output3 (.I(net3),
    .Z(segm[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output4 (.I(net4),
    .Z(segm[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output5 (.I(net5),
    .Z(segm[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output6 (.I(net6),
    .Z(segm[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output7 (.I(net7),
    .Z(segm[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output8 (.I(net8),
    .Z(segm[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output9 (.I(net9),
    .Z(segm[7]));
 assign segm[0] = net24;
 assign segm[3] = net25;
 assign segm[5] = net26;
endmodule

