magic
tech gf180mcuD
magscale 1 5
timestamp 1699642008
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 9417 19055 9423 19081
rect 9449 19055 9455 19081
rect 11097 19055 11103 19081
rect 11129 19055 11135 19081
rect 8969 18999 8975 19025
rect 9001 18999 9007 19025
rect 11881 18999 11887 19025
rect 11913 18999 11919 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 10375 18745 10401 18751
rect 10375 18713 10401 18719
rect 13119 18745 13145 18751
rect 13119 18713 13145 18719
rect 9865 18607 9871 18633
rect 9897 18607 9903 18633
rect 12609 18607 12615 18633
rect 12641 18607 12647 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 8695 18353 8721 18359
rect 8695 18321 8721 18327
rect 8185 18215 8191 18241
rect 8217 18215 8223 18241
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 9479 14041 9505 14047
rect 9305 14015 9311 14041
rect 9337 14015 9343 14041
rect 9479 14009 9505 14015
rect 11495 14041 11521 14047
rect 11495 14009 11521 14015
rect 11215 13985 11241 13991
rect 11215 13953 11241 13959
rect 11271 13929 11297 13935
rect 11271 13897 11297 13903
rect 11551 13929 11577 13935
rect 11551 13897 11577 13903
rect 11215 13817 11241 13823
rect 11215 13785 11241 13791
rect 11495 13817 11521 13823
rect 11495 13785 11521 13791
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 20007 13593 20033 13599
rect 9697 13567 9703 13593
rect 9729 13567 9735 13593
rect 11209 13567 11215 13593
rect 11241 13567 11247 13593
rect 12273 13567 12279 13593
rect 12305 13567 12311 13593
rect 20007 13561 20033 13567
rect 12503 13537 12529 13543
rect 8297 13511 8303 13537
rect 8329 13511 8335 13537
rect 10873 13511 10879 13537
rect 10905 13511 10911 13537
rect 18937 13511 18943 13537
rect 18969 13511 18975 13537
rect 12503 13505 12529 13511
rect 7967 13481 7993 13487
rect 7967 13449 7993 13455
rect 8023 13481 8049 13487
rect 8633 13455 8639 13481
rect 8665 13455 8671 13481
rect 8023 13449 8049 13455
rect 8135 13425 8161 13431
rect 8135 13393 8161 13399
rect 9927 13425 9953 13431
rect 9927 13393 9953 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 9423 13257 9449 13263
rect 9423 13225 9449 13231
rect 11663 13257 11689 13263
rect 11663 13225 11689 13231
rect 11775 13257 11801 13263
rect 11775 13225 11801 13231
rect 9087 13201 9113 13207
rect 9087 13169 9113 13175
rect 9143 13201 9169 13207
rect 9143 13169 9169 13175
rect 9479 13201 9505 13207
rect 9479 13169 9505 13175
rect 9255 13145 9281 13151
rect 11831 13145 11857 13151
rect 2137 13119 2143 13145
rect 2169 13119 2175 13145
rect 6841 13119 6847 13145
rect 6873 13119 6879 13145
rect 8857 13119 8863 13145
rect 8889 13119 8895 13145
rect 9977 13119 9983 13145
rect 10009 13119 10015 13145
rect 13057 13119 13063 13145
rect 13089 13119 13095 13145
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 9255 13113 9281 13119
rect 11831 13113 11857 13119
rect 9815 13089 9841 13095
rect 14687 13089 14713 13095
rect 7177 13063 7183 13089
rect 7209 13063 7215 13089
rect 8241 13063 8247 13089
rect 8273 13063 8279 13089
rect 9081 13063 9087 13089
rect 9113 13063 9119 13089
rect 10369 13063 10375 13089
rect 10401 13063 10407 13089
rect 11433 13063 11439 13089
rect 11465 13063 11471 13089
rect 13393 13063 13399 13089
rect 13425 13063 13431 13089
rect 14457 13063 14463 13089
rect 14489 13063 14495 13089
rect 9815 13057 9841 13063
rect 14687 13057 14713 13063
rect 967 13033 993 13039
rect 967 13001 993 13007
rect 20007 13033 20033 13039
rect 20007 13001 20033 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 10319 12865 10345 12871
rect 10319 12833 10345 12839
rect 9311 12809 9337 12815
rect 9311 12777 9337 12783
rect 7351 12753 7377 12759
rect 7351 12721 7377 12727
rect 7575 12753 7601 12759
rect 7575 12721 7601 12727
rect 8079 12753 8105 12759
rect 8079 12721 8105 12727
rect 8247 12753 8273 12759
rect 8247 12721 8273 12727
rect 10375 12753 10401 12759
rect 10375 12721 10401 12727
rect 13455 12753 13481 12759
rect 13455 12721 13481 12727
rect 13623 12753 13649 12759
rect 13623 12721 13649 12727
rect 14071 12753 14097 12759
rect 14071 12721 14097 12727
rect 14239 12753 14265 12759
rect 14239 12721 14265 12727
rect 14575 12753 14601 12759
rect 14575 12721 14601 12727
rect 7183 12697 7209 12703
rect 7183 12665 7209 12671
rect 7239 12697 7265 12703
rect 7239 12665 7265 12671
rect 7463 12697 7489 12703
rect 7463 12665 7489 12671
rect 7743 12697 7769 12703
rect 7743 12665 7769 12671
rect 7911 12697 7937 12703
rect 7911 12665 7937 12671
rect 9255 12697 9281 12703
rect 9255 12665 9281 12671
rect 9479 12697 9505 12703
rect 9479 12665 9505 12671
rect 10319 12697 10345 12703
rect 10319 12665 10345 12671
rect 13959 12697 13985 12703
rect 13959 12665 13985 12671
rect 14183 12697 14209 12703
rect 14183 12665 14209 12671
rect 14631 12697 14657 12703
rect 14631 12665 14657 12671
rect 14743 12697 14769 12703
rect 14743 12665 14769 12671
rect 7519 12641 7545 12647
rect 7519 12609 7545 12615
rect 8079 12641 8105 12647
rect 8079 12609 8105 12615
rect 8415 12641 8441 12647
rect 8415 12609 8441 12615
rect 9367 12641 9393 12647
rect 9367 12609 9393 12615
rect 11215 12641 11241 12647
rect 11215 12609 11241 12615
rect 13567 12641 13593 12647
rect 13567 12609 13593 12615
rect 13791 12641 13817 12647
rect 13791 12609 13817 12615
rect 13903 12641 13929 12647
rect 13903 12609 13929 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 11271 12473 11297 12479
rect 11657 12447 11663 12473
rect 11689 12447 11695 12473
rect 11271 12441 11297 12447
rect 12055 12417 12081 12423
rect 7121 12391 7127 12417
rect 7153 12391 7159 12417
rect 13729 12391 13735 12417
rect 13761 12391 13767 12417
rect 12055 12385 12081 12391
rect 11551 12361 11577 12367
rect 11999 12361 12025 12367
rect 7513 12335 7519 12361
rect 7545 12335 7551 12361
rect 9641 12335 9647 12361
rect 9673 12335 9679 12361
rect 11377 12335 11383 12361
rect 11409 12335 11415 12361
rect 11769 12335 11775 12361
rect 11801 12335 11807 12361
rect 11551 12329 11577 12335
rect 11999 12329 12025 12335
rect 12167 12361 12193 12367
rect 15023 12361 15049 12367
rect 13337 12335 13343 12361
rect 13369 12335 13375 12361
rect 12167 12329 12193 12335
rect 15023 12329 15049 12335
rect 7743 12305 7769 12311
rect 6057 12279 6063 12305
rect 6089 12279 6095 12305
rect 10033 12279 10039 12305
rect 10065 12279 10071 12305
rect 11097 12279 11103 12305
rect 11129 12279 11135 12305
rect 14793 12279 14799 12305
rect 14825 12279 14831 12305
rect 7743 12273 7769 12279
rect 11215 12249 11241 12255
rect 11215 12217 11241 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 9591 12081 9617 12087
rect 9591 12049 9617 12055
rect 967 12025 993 12031
rect 7071 12025 7097 12031
rect 20007 12025 20033 12031
rect 4993 11999 4999 12025
rect 5025 11999 5031 12025
rect 13001 11999 13007 12025
rect 13033 11999 13039 12025
rect 967 11993 993 11999
rect 7071 11993 7097 11999
rect 20007 11993 20033 11999
rect 9647 11969 9673 11975
rect 13231 11969 13257 11975
rect 2137 11943 2143 11969
rect 2169 11943 2175 11969
rect 6449 11943 6455 11969
rect 6481 11943 6487 11969
rect 9921 11943 9927 11969
rect 9953 11943 9959 11969
rect 10313 11943 10319 11969
rect 10345 11943 10351 11969
rect 10761 11943 10767 11969
rect 10793 11943 10799 11969
rect 10985 11943 10991 11969
rect 11017 11943 11023 11969
rect 11601 11943 11607 11969
rect 11633 11943 11639 11969
rect 18825 11943 18831 11969
rect 18857 11943 18863 11969
rect 9647 11937 9673 11943
rect 13231 11937 13257 11943
rect 6791 11913 6817 11919
rect 6057 11887 6063 11913
rect 6089 11887 6095 11913
rect 6791 11881 6817 11887
rect 6847 11913 6873 11919
rect 6847 11881 6873 11887
rect 7967 11913 7993 11919
rect 7967 11881 7993 11887
rect 8807 11913 8833 11919
rect 10369 11887 10375 11913
rect 10401 11887 10407 11913
rect 11937 11887 11943 11913
rect 11969 11887 11975 11913
rect 8807 11881 8833 11887
rect 6679 11857 6705 11863
rect 6679 11825 6705 11831
rect 8023 11857 8049 11863
rect 8023 11825 8049 11831
rect 8135 11857 8161 11863
rect 8135 11825 8161 11831
rect 8415 11857 8441 11863
rect 8415 11825 8441 11831
rect 8639 11857 8665 11863
rect 8639 11825 8665 11831
rect 8751 11857 8777 11863
rect 8751 11825 8777 11831
rect 11047 11857 11073 11863
rect 11047 11825 11073 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 6455 11689 6481 11695
rect 6455 11657 6481 11663
rect 12055 11689 12081 11695
rect 12055 11657 12081 11663
rect 8695 11633 8721 11639
rect 8695 11601 8721 11607
rect 9087 11633 9113 11639
rect 9087 11601 9113 11607
rect 9591 11633 9617 11639
rect 11999 11633 12025 11639
rect 10201 11607 10207 11633
rect 10233 11607 10239 11633
rect 10649 11607 10655 11633
rect 10681 11607 10687 11633
rect 9591 11601 9617 11607
rect 11999 11601 12025 11607
rect 12167 11633 12193 11639
rect 12167 11601 12193 11607
rect 14183 11633 14209 11639
rect 14737 11607 14743 11633
rect 14769 11607 14775 11633
rect 14183 11601 14209 11607
rect 6399 11577 6425 11583
rect 2137 11551 2143 11577
rect 2169 11551 2175 11577
rect 6399 11545 6425 11551
rect 6511 11577 6537 11583
rect 8863 11577 8889 11583
rect 6673 11551 6679 11577
rect 6705 11551 6711 11577
rect 8297 11551 8303 11577
rect 8329 11551 8335 11577
rect 6511 11545 6537 11551
rect 8863 11545 8889 11551
rect 9143 11577 9169 11583
rect 9143 11545 9169 11551
rect 9311 11577 9337 11583
rect 11887 11577 11913 11583
rect 9473 11551 9479 11577
rect 9505 11551 9511 11577
rect 10425 11551 10431 11577
rect 10457 11551 10463 11577
rect 10537 11551 10543 11577
rect 10569 11551 10575 11577
rect 14065 11551 14071 11577
rect 14097 11551 14103 11577
rect 14345 11551 14351 11577
rect 14377 11551 14383 11577
rect 18825 11551 18831 11577
rect 18857 11551 18863 11577
rect 9311 11545 9337 11551
rect 11887 11545 11913 11551
rect 16031 11521 16057 11527
rect 6841 11495 6847 11521
rect 6873 11495 6879 11521
rect 7905 11495 7911 11521
rect 7937 11495 7943 11521
rect 10313 11495 10319 11521
rect 10345 11495 10351 11521
rect 15801 11495 15807 11521
rect 15833 11495 15839 11521
rect 16031 11489 16057 11495
rect 967 11465 993 11471
rect 967 11433 993 11439
rect 9199 11465 9225 11471
rect 9199 11433 9225 11439
rect 9647 11465 9673 11471
rect 9647 11433 9673 11439
rect 20007 11465 20033 11471
rect 20007 11433 20033 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 8415 11297 8441 11303
rect 14961 11271 14967 11297
rect 14993 11271 14999 11297
rect 8415 11265 8441 11271
rect 967 11241 993 11247
rect 14015 11241 14041 11247
rect 12217 11215 12223 11241
rect 12249 11215 12255 11241
rect 12497 11215 12503 11241
rect 12529 11215 12535 11241
rect 967 11209 993 11215
rect 14015 11209 14041 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 7911 11185 7937 11191
rect 2137 11159 2143 11185
rect 2169 11159 2175 11185
rect 7911 11153 7937 11159
rect 8079 11185 8105 11191
rect 8079 11153 8105 11159
rect 8247 11185 8273 11191
rect 8247 11153 8273 11159
rect 8471 11185 8497 11191
rect 8471 11153 8497 11159
rect 9591 11185 9617 11191
rect 9591 11153 9617 11159
rect 9927 11185 9953 11191
rect 9927 11153 9953 11159
rect 10039 11185 10065 11191
rect 10039 11153 10065 11159
rect 10263 11185 10289 11191
rect 10263 11153 10289 11159
rect 10711 11185 10737 11191
rect 14127 11185 14153 11191
rect 12273 11159 12279 11185
rect 12305 11159 12311 11185
rect 10711 11153 10737 11159
rect 14127 11153 14153 11159
rect 14687 11185 14713 11191
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 14687 11153 14713 11159
rect 8695 11129 8721 11135
rect 8695 11097 8721 11103
rect 8807 11129 8833 11135
rect 12895 11129 12921 11135
rect 11377 11103 11383 11129
rect 11409 11103 11415 11129
rect 11825 11103 11831 11129
rect 11857 11103 11863 11129
rect 8807 11097 8833 11103
rect 12895 11097 12921 11103
rect 12951 11129 12977 11135
rect 12951 11097 12977 11103
rect 14631 11129 14657 11135
rect 14631 11097 14657 11103
rect 14743 11129 14769 11135
rect 14743 11097 14769 11103
rect 8079 11073 8105 11079
rect 8079 11041 8105 11047
rect 8415 11073 8441 11079
rect 8415 11041 8441 11047
rect 8751 11073 8777 11079
rect 9143 11073 9169 11079
rect 8969 11047 8975 11073
rect 9001 11047 9007 11073
rect 8751 11041 8777 11047
rect 9143 11041 9169 11047
rect 9311 11073 9337 11079
rect 9311 11041 9337 11047
rect 10095 11073 10121 11079
rect 10095 11041 10121 11047
rect 12727 11073 12753 11079
rect 12727 11041 12753 11047
rect 13063 11073 13089 11079
rect 14289 11047 14295 11073
rect 14321 11047 14327 11073
rect 13063 11041 13089 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 7127 10905 7153 10911
rect 7127 10873 7153 10879
rect 7743 10905 7769 10911
rect 7743 10873 7769 10879
rect 11495 10905 11521 10911
rect 11495 10873 11521 10879
rect 14407 10905 14433 10911
rect 14407 10873 14433 10879
rect 11607 10849 11633 10855
rect 7569 10823 7575 10849
rect 7601 10823 7607 10849
rect 11607 10817 11633 10823
rect 6679 10793 6705 10799
rect 6393 10767 6399 10793
rect 6425 10767 6431 10793
rect 6561 10767 6567 10793
rect 6593 10767 6599 10793
rect 6679 10761 6705 10767
rect 6791 10793 6817 10799
rect 11663 10793 11689 10799
rect 6897 10767 6903 10793
rect 6929 10767 6935 10793
rect 11321 10767 11327 10793
rect 11353 10767 11359 10793
rect 14177 10767 14183 10793
rect 14209 10767 14215 10793
rect 6791 10761 6817 10767
rect 11663 10761 11689 10767
rect 6735 10737 6761 10743
rect 4937 10711 4943 10737
rect 4969 10711 4975 10737
rect 6001 10711 6007 10737
rect 6033 10711 6039 10737
rect 8801 10711 8807 10737
rect 8833 10711 8839 10737
rect 12721 10711 12727 10737
rect 12753 10711 12759 10737
rect 13785 10711 13791 10737
rect 13817 10711 13823 10737
rect 6735 10705 6761 10711
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 5895 10513 5921 10519
rect 5895 10481 5921 10487
rect 10039 10513 10065 10519
rect 10039 10481 10065 10487
rect 13567 10513 13593 10519
rect 13567 10481 13593 10487
rect 13791 10513 13817 10519
rect 13791 10481 13817 10487
rect 967 10457 993 10463
rect 967 10425 993 10431
rect 5839 10457 5865 10463
rect 14519 10457 14545 10463
rect 7961 10431 7967 10457
rect 7993 10431 7999 10457
rect 9025 10431 9031 10457
rect 9057 10431 9063 10457
rect 5839 10425 5865 10431
rect 14519 10425 14545 10431
rect 20007 10457 20033 10463
rect 20007 10425 20033 10431
rect 10095 10401 10121 10407
rect 2081 10375 2087 10401
rect 2113 10375 2119 10401
rect 7569 10375 7575 10401
rect 7601 10375 7607 10401
rect 9361 10375 9367 10401
rect 9393 10375 9399 10401
rect 10095 10369 10121 10375
rect 10207 10401 10233 10407
rect 13679 10401 13705 10407
rect 14799 10401 14825 10407
rect 10313 10375 10319 10401
rect 10345 10375 10351 10401
rect 10649 10375 10655 10401
rect 10681 10375 10687 10401
rect 13449 10375 13455 10401
rect 13481 10375 13487 10401
rect 14121 10375 14127 10401
rect 14153 10375 14159 10401
rect 10207 10369 10233 10375
rect 13679 10369 13705 10375
rect 14799 10369 14825 10375
rect 14855 10401 14881 10407
rect 18825 10375 18831 10401
rect 18857 10375 18863 10401
rect 14855 10369 14881 10375
rect 13847 10345 13873 10351
rect 9417 10319 9423 10345
rect 9449 10319 9455 10345
rect 9753 10319 9759 10345
rect 9785 10319 9791 10345
rect 12553 10319 12559 10345
rect 12585 10319 12591 10345
rect 13847 10313 13873 10319
rect 14575 10345 14601 10351
rect 14575 10313 14601 10319
rect 14015 10289 14041 10295
rect 9585 10263 9591 10289
rect 9617 10263 9623 10289
rect 14015 10257 14041 10263
rect 14687 10289 14713 10295
rect 14687 10257 14713 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 8857 10095 8863 10121
rect 8889 10095 8895 10121
rect 6169 10039 6175 10065
rect 6201 10039 6207 10065
rect 9361 10039 9367 10065
rect 9393 10039 9399 10065
rect 11265 10039 11271 10065
rect 11297 10039 11303 10065
rect 6623 10009 6649 10015
rect 2137 9983 2143 10009
rect 2169 9983 2175 10009
rect 6281 9983 6287 10009
rect 6313 9983 6319 10009
rect 6505 9983 6511 10009
rect 6537 9983 6543 10009
rect 6623 9977 6649 9983
rect 6735 10009 6761 10015
rect 10263 10009 10289 10015
rect 6841 9983 6847 10009
rect 6873 9983 6879 10009
rect 8745 9983 8751 10009
rect 8777 9983 8783 10009
rect 9809 9983 9815 10009
rect 9841 9983 9847 10009
rect 10649 9983 10655 10009
rect 10681 9983 10687 10009
rect 11041 9983 11047 10009
rect 11073 9983 11079 10009
rect 11321 9983 11327 10009
rect 11353 9983 11359 10009
rect 11601 9983 11607 10009
rect 11633 9983 11639 10009
rect 11825 9983 11831 10009
rect 11857 9983 11863 10009
rect 12609 9983 12615 10009
rect 12641 9983 12647 10009
rect 6735 9977 6761 9983
rect 10263 9977 10289 9983
rect 5727 9953 5753 9959
rect 5727 9921 5753 9927
rect 6679 9953 6705 9959
rect 6679 9921 6705 9927
rect 8415 9953 8441 9959
rect 11439 9953 11465 9959
rect 15471 9953 15497 9959
rect 9865 9927 9871 9953
rect 9897 9927 9903 9953
rect 14569 9927 14575 9953
rect 14601 9927 14607 9953
rect 8415 9921 8441 9927
rect 11439 9921 11465 9927
rect 15471 9921 15497 9927
rect 967 9897 993 9903
rect 967 9865 993 9871
rect 5783 9897 5809 9903
rect 15415 9897 15441 9903
rect 11601 9871 11607 9897
rect 11633 9871 11639 9897
rect 5783 9865 5809 9871
rect 15415 9865 15441 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 6959 9729 6985 9735
rect 6959 9697 6985 9703
rect 13511 9729 13537 9735
rect 13511 9697 13537 9703
rect 967 9673 993 9679
rect 8639 9673 8665 9679
rect 4825 9647 4831 9673
rect 4857 9647 4863 9673
rect 5889 9647 5895 9673
rect 5921 9647 5927 9673
rect 967 9641 993 9647
rect 8639 9641 8665 9647
rect 9423 9673 9449 9679
rect 9423 9641 9449 9647
rect 10431 9673 10457 9679
rect 10431 9641 10457 9647
rect 12503 9673 12529 9679
rect 12503 9641 12529 9647
rect 13399 9673 13425 9679
rect 16025 9647 16031 9673
rect 16057 9647 16063 9673
rect 13399 9641 13425 9647
rect 6679 9617 6705 9623
rect 2137 9591 2143 9617
rect 2169 9591 2175 9617
rect 6281 9591 6287 9617
rect 6313 9591 6319 9617
rect 6679 9585 6705 9591
rect 6903 9617 6929 9623
rect 6903 9585 6929 9591
rect 7071 9617 7097 9623
rect 7071 9585 7097 9591
rect 7183 9617 7209 9623
rect 9087 9617 9113 9623
rect 11159 9617 11185 9623
rect 8969 9591 8975 9617
rect 9001 9591 9007 9617
rect 9641 9591 9647 9617
rect 9673 9591 9679 9617
rect 9809 9591 9815 9617
rect 9841 9591 9847 9617
rect 7183 9585 7209 9591
rect 9087 9585 9113 9591
rect 11159 9585 11185 9591
rect 11495 9617 11521 9623
rect 11495 9585 11521 9591
rect 11663 9617 11689 9623
rect 12279 9617 12305 9623
rect 12049 9591 12055 9617
rect 12081 9591 12087 9617
rect 11663 9585 11689 9591
rect 12279 9585 12305 9591
rect 12391 9617 12417 9623
rect 12391 9585 12417 9591
rect 12559 9617 12585 9623
rect 12559 9585 12585 9591
rect 12727 9617 12753 9623
rect 12727 9585 12753 9591
rect 12895 9617 12921 9623
rect 13791 9617 13817 9623
rect 13673 9591 13679 9617
rect 13705 9591 13711 9617
rect 12895 9585 12921 9591
rect 13791 9585 13817 9591
rect 14071 9617 14097 9623
rect 14071 9585 14097 9591
rect 14183 9617 14209 9623
rect 14183 9585 14209 9591
rect 14295 9617 14321 9623
rect 14569 9591 14575 9617
rect 14601 9591 14607 9617
rect 14295 9585 14321 9591
rect 11271 9561 11297 9567
rect 9305 9535 9311 9561
rect 9337 9535 9343 9561
rect 10761 9535 10767 9561
rect 10793 9535 10799 9561
rect 10929 9535 10935 9561
rect 10961 9535 10967 9561
rect 11271 9529 11297 9535
rect 11775 9561 11801 9567
rect 13057 9535 13063 9561
rect 13089 9535 13095 9561
rect 13953 9535 13959 9561
rect 13985 9535 13991 9561
rect 14961 9535 14967 9561
rect 14993 9535 14999 9561
rect 11775 9529 11801 9535
rect 11663 9505 11689 9511
rect 6897 9479 6903 9505
rect 6929 9479 6935 9505
rect 11663 9473 11689 9479
rect 14351 9505 14377 9511
rect 14351 9473 14377 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 9255 9337 9281 9343
rect 7737 9311 7743 9337
rect 7769 9311 7775 9337
rect 9255 9305 9281 9311
rect 11831 9337 11857 9343
rect 11831 9305 11857 9311
rect 12279 9337 12305 9343
rect 12279 9305 12305 9311
rect 12223 9281 12249 9287
rect 12223 9249 12249 9255
rect 13399 9281 13425 9287
rect 13399 9249 13425 9255
rect 13679 9281 13705 9287
rect 13679 9249 13705 9255
rect 6567 9225 6593 9231
rect 5945 9199 5951 9225
rect 5977 9199 5983 9225
rect 6337 9199 6343 9225
rect 6369 9199 6375 9225
rect 6567 9193 6593 9199
rect 7911 9225 7937 9231
rect 7911 9193 7937 9199
rect 9535 9225 9561 9231
rect 9535 9193 9561 9199
rect 9759 9225 9785 9231
rect 9759 9193 9785 9199
rect 10039 9225 10065 9231
rect 10655 9225 10681 9231
rect 11439 9225 11465 9231
rect 10425 9199 10431 9225
rect 10457 9199 10463 9225
rect 10873 9199 10879 9225
rect 10905 9199 10911 9225
rect 10039 9193 10065 9199
rect 10655 9193 10681 9199
rect 11439 9193 11465 9199
rect 11775 9225 11801 9231
rect 11775 9193 11801 9199
rect 12391 9225 12417 9231
rect 12391 9193 12417 9199
rect 12951 9225 12977 9231
rect 12951 9193 12977 9199
rect 13623 9225 13649 9231
rect 13623 9193 13649 9199
rect 13791 9225 13817 9231
rect 14121 9199 14127 9225
rect 14153 9199 14159 9225
rect 18937 9199 18943 9225
rect 18969 9199 18975 9225
rect 13791 9193 13817 9199
rect 6511 9169 6537 9175
rect 4881 9143 4887 9169
rect 4913 9143 4919 9169
rect 6511 9137 6537 9143
rect 6791 9169 6817 9175
rect 11103 9169 11129 9175
rect 12839 9169 12865 9175
rect 15751 9169 15777 9175
rect 10257 9143 10263 9169
rect 10289 9143 10295 9169
rect 11265 9143 11271 9169
rect 11297 9143 11303 9169
rect 11601 9143 11607 9169
rect 11633 9143 11639 9169
rect 13113 9143 13119 9169
rect 13145 9143 13151 9169
rect 13449 9143 13455 9169
rect 13481 9143 13487 9169
rect 14457 9143 14463 9169
rect 14489 9143 14495 9169
rect 15521 9143 15527 9169
rect 15553 9143 15559 9169
rect 6791 9137 6817 9143
rect 11103 9137 11129 9143
rect 12839 9137 12865 9143
rect 15751 9137 15777 9143
rect 13287 9113 13313 9119
rect 13287 9081 13313 9087
rect 20007 9113 20033 9119
rect 20007 9081 20033 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 7743 8945 7769 8951
rect 7743 8913 7769 8919
rect 9311 8945 9337 8951
rect 9311 8913 9337 8919
rect 9535 8945 9561 8951
rect 9535 8913 9561 8919
rect 9703 8945 9729 8951
rect 9703 8913 9729 8919
rect 15079 8945 15105 8951
rect 15079 8913 15105 8919
rect 967 8889 993 8895
rect 967 8857 993 8863
rect 7407 8889 7433 8895
rect 7407 8857 7433 8863
rect 7687 8889 7713 8895
rect 7687 8857 7713 8863
rect 20007 8889 20033 8895
rect 20007 8857 20033 8863
rect 8079 8833 8105 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 7233 8807 7239 8833
rect 7265 8807 7271 8833
rect 7905 8807 7911 8833
rect 7937 8807 7943 8833
rect 8079 8801 8105 8807
rect 8303 8833 8329 8839
rect 8303 8801 8329 8807
rect 9367 8833 9393 8839
rect 9367 8801 9393 8807
rect 9871 8833 9897 8839
rect 9871 8801 9897 8807
rect 9927 8833 9953 8839
rect 10767 8833 10793 8839
rect 10089 8807 10095 8833
rect 10121 8807 10127 8833
rect 9927 8801 9953 8807
rect 10767 8801 10793 8807
rect 10935 8833 10961 8839
rect 10935 8801 10961 8807
rect 12671 8833 12697 8839
rect 12671 8801 12697 8807
rect 12839 8833 12865 8839
rect 12839 8801 12865 8807
rect 13007 8833 13033 8839
rect 13007 8801 13033 8807
rect 14575 8833 14601 8839
rect 14575 8801 14601 8807
rect 14687 8833 14713 8839
rect 14687 8801 14713 8807
rect 14911 8833 14937 8839
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 14911 8801 14937 8807
rect 8863 8777 8889 8783
rect 8185 8751 8191 8777
rect 8217 8751 8223 8777
rect 8863 8745 8889 8751
rect 9031 8777 9057 8783
rect 9031 8745 9057 8751
rect 10655 8777 10681 8783
rect 10655 8745 10681 8751
rect 15023 8777 15049 8783
rect 15023 8745 15049 8751
rect 6455 8721 6481 8727
rect 6455 8689 6481 8695
rect 7351 8721 7377 8727
rect 7351 8689 7377 8695
rect 7911 8721 7937 8727
rect 7911 8689 7937 8695
rect 8975 8721 9001 8727
rect 8975 8689 9001 8695
rect 9311 8721 9337 8727
rect 9311 8689 9337 8695
rect 9647 8721 9673 8727
rect 9647 8689 9673 8695
rect 10767 8721 10793 8727
rect 10767 8689 10793 8695
rect 12895 8721 12921 8727
rect 12895 8689 12921 8695
rect 14295 8721 14321 8727
rect 14295 8689 14321 8695
rect 14743 8721 14769 8727
rect 14743 8689 14769 8695
rect 15079 8721 15105 8727
rect 15079 8689 15105 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 9703 8553 9729 8559
rect 11775 8553 11801 8559
rect 11041 8527 11047 8553
rect 11073 8527 11079 8553
rect 9703 8521 9729 8527
rect 11775 8521 11801 8527
rect 12839 8553 12865 8559
rect 12839 8521 12865 8527
rect 7575 8497 7601 8503
rect 12951 8497 12977 8503
rect 9305 8471 9311 8497
rect 9337 8471 9343 8497
rect 10537 8471 10543 8497
rect 10569 8471 10575 8497
rect 11377 8471 11383 8497
rect 11409 8471 11415 8497
rect 7575 8465 7601 8471
rect 12951 8465 12977 8471
rect 7743 8441 7769 8447
rect 9759 8441 9785 8447
rect 10879 8441 10905 8447
rect 2137 8415 2143 8441
rect 2169 8415 2175 8441
rect 7401 8415 7407 8441
rect 7433 8415 7439 8441
rect 9417 8415 9423 8441
rect 9449 8415 9455 8441
rect 10425 8415 10431 8441
rect 10457 8415 10463 8441
rect 7743 8409 7769 8415
rect 9759 8409 9785 8415
rect 10879 8409 10905 8415
rect 11215 8441 11241 8447
rect 11215 8409 11241 8415
rect 13007 8441 13033 8447
rect 15527 8441 15553 8447
rect 13841 8415 13847 8441
rect 13873 8415 13879 8441
rect 18825 8415 18831 8441
rect 18857 8415 18863 8441
rect 13007 8409 13033 8415
rect 15527 8409 15553 8415
rect 7631 8385 7657 8391
rect 5945 8359 5951 8385
rect 5977 8359 5983 8385
rect 7009 8359 7015 8385
rect 7041 8359 7047 8385
rect 7631 8353 7657 8359
rect 8079 8385 8105 8391
rect 8079 8353 8105 8359
rect 9871 8385 9897 8391
rect 9871 8353 9897 8359
rect 11663 8385 11689 8391
rect 14233 8359 14239 8385
rect 14265 8359 14271 8385
rect 15297 8359 15303 8385
rect 15329 8359 15335 8385
rect 19945 8359 19951 8385
rect 19977 8359 19983 8385
rect 11663 8353 11689 8359
rect 967 8329 993 8335
rect 967 8297 993 8303
rect 7799 8329 7825 8335
rect 7799 8297 7825 8303
rect 9703 8329 9729 8335
rect 9703 8297 9729 8303
rect 11831 8329 11857 8335
rect 11831 8297 11857 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 7127 8161 7153 8167
rect 7127 8129 7153 8135
rect 7183 8161 7209 8167
rect 7183 8129 7209 8135
rect 7295 8161 7321 8167
rect 7295 8129 7321 8135
rect 7351 8161 7377 8167
rect 7351 8129 7377 8135
rect 9927 8161 9953 8167
rect 9927 8129 9953 8135
rect 14183 8161 14209 8167
rect 14183 8129 14209 8135
rect 7743 8105 7769 8111
rect 13007 8105 13033 8111
rect 11321 8079 11327 8105
rect 11353 8079 11359 8105
rect 12385 8079 12391 8105
rect 12417 8079 12423 8105
rect 7743 8073 7769 8079
rect 13007 8073 13033 8079
rect 20007 8105 20033 8111
rect 20007 8073 20033 8079
rect 9703 8049 9729 8055
rect 9249 8023 9255 8049
rect 9281 8023 9287 8049
rect 9703 8017 9729 8023
rect 9871 8049 9897 8055
rect 12777 8023 12783 8049
rect 12809 8023 12815 8049
rect 15017 8023 15023 8049
rect 15049 8023 15055 8049
rect 18825 8023 18831 8049
rect 18857 8023 18863 8049
rect 9871 8017 9897 8023
rect 7631 7993 7657 7999
rect 7631 7961 7657 7967
rect 7687 7993 7713 7999
rect 14183 7993 14209 7999
rect 9361 7967 9367 7993
rect 9393 7967 9399 7993
rect 9529 7967 9535 7993
rect 9561 7967 9567 7993
rect 7687 7961 7713 7967
rect 14183 7961 14209 7967
rect 14239 7993 14265 7999
rect 14239 7961 14265 7967
rect 14519 7993 14545 7999
rect 14519 7961 14545 7967
rect 14631 7993 14657 7999
rect 14631 7961 14657 7967
rect 14687 7993 14713 7999
rect 14687 7961 14713 7967
rect 15135 7937 15161 7943
rect 15135 7905 15161 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 11495 7769 11521 7775
rect 9977 7743 9983 7769
rect 10009 7743 10015 7769
rect 11495 7737 11521 7743
rect 12111 7769 12137 7775
rect 12111 7737 12137 7743
rect 14295 7769 14321 7775
rect 14295 7737 14321 7743
rect 7911 7713 7937 7719
rect 7009 7687 7015 7713
rect 7041 7687 7047 7713
rect 7911 7681 7937 7687
rect 9703 7713 9729 7719
rect 9703 7681 9729 7687
rect 10655 7713 10681 7719
rect 11769 7687 11775 7713
rect 11801 7687 11807 7713
rect 13001 7687 13007 7713
rect 13033 7687 13039 7713
rect 10655 7681 10681 7687
rect 10151 7657 10177 7663
rect 7345 7631 7351 7657
rect 7377 7631 7383 7657
rect 9417 7631 9423 7657
rect 9449 7631 9455 7657
rect 10151 7625 10177 7631
rect 10375 7657 10401 7663
rect 11887 7657 11913 7663
rect 11601 7631 11607 7657
rect 11633 7631 11639 7657
rect 12665 7631 12671 7657
rect 12697 7631 12703 7657
rect 10375 7625 10401 7631
rect 11887 7625 11913 7631
rect 7631 7601 7657 7607
rect 12167 7601 12193 7607
rect 5945 7575 5951 7601
rect 5977 7575 5983 7601
rect 9305 7575 9311 7601
rect 9337 7575 9343 7601
rect 14065 7575 14071 7601
rect 14097 7575 14103 7601
rect 7631 7569 7657 7575
rect 12167 7569 12193 7575
rect 7855 7545 7881 7551
rect 11601 7519 11607 7545
rect 11633 7519 11639 7545
rect 7855 7513 7881 7519
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 8689 7295 8695 7321
rect 8721 7295 8727 7321
rect 9249 7295 9255 7321
rect 9281 7295 9287 7321
rect 10313 7295 10319 7321
rect 10345 7295 10351 7321
rect 11489 7295 11495 7321
rect 11521 7295 11527 7321
rect 12553 7295 12559 7321
rect 12585 7295 12591 7321
rect 10711 7265 10737 7271
rect 12839 7265 12865 7271
rect 7233 7239 7239 7265
rect 7265 7239 7271 7265
rect 8913 7239 8919 7265
rect 8945 7239 8951 7265
rect 11153 7239 11159 7265
rect 11185 7239 11191 7265
rect 10711 7233 10737 7239
rect 12839 7233 12865 7239
rect 7625 7183 7631 7209
rect 7657 7183 7663 7209
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 8863 6985 8889 6991
rect 8863 6953 8889 6959
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 12783 19111 12809 19137
rect 9423 19055 9449 19081
rect 11103 19055 11129 19081
rect 8975 18999 9001 19025
rect 11887 18999 11913 19025
rect 12279 18999 12305 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 10375 18719 10401 18745
rect 13119 18719 13145 18745
rect 9871 18607 9897 18633
rect 12615 18607 12641 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 8695 18327 8721 18353
rect 8191 18215 8217 18241
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 9311 14015 9337 14041
rect 9479 14015 9505 14041
rect 11495 14015 11521 14041
rect 11215 13959 11241 13985
rect 11271 13903 11297 13929
rect 11551 13903 11577 13929
rect 11215 13791 11241 13817
rect 11495 13791 11521 13817
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 9703 13567 9729 13593
rect 11215 13567 11241 13593
rect 12279 13567 12305 13593
rect 20007 13567 20033 13593
rect 8303 13511 8329 13537
rect 10879 13511 10905 13537
rect 12503 13511 12529 13537
rect 18943 13511 18969 13537
rect 7967 13455 7993 13481
rect 8023 13455 8049 13481
rect 8639 13455 8665 13481
rect 8135 13399 8161 13425
rect 9927 13399 9953 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 9423 13231 9449 13257
rect 11663 13231 11689 13257
rect 11775 13231 11801 13257
rect 9087 13175 9113 13201
rect 9143 13175 9169 13201
rect 9479 13175 9505 13201
rect 2143 13119 2169 13145
rect 6847 13119 6873 13145
rect 8863 13119 8889 13145
rect 9255 13119 9281 13145
rect 9983 13119 10009 13145
rect 11831 13119 11857 13145
rect 13063 13119 13089 13145
rect 18831 13119 18857 13145
rect 7183 13063 7209 13089
rect 8247 13063 8273 13089
rect 9087 13063 9113 13089
rect 9815 13063 9841 13089
rect 10375 13063 10401 13089
rect 11439 13063 11465 13089
rect 13399 13063 13425 13089
rect 14463 13063 14489 13089
rect 14687 13063 14713 13089
rect 967 13007 993 13033
rect 20007 13007 20033 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 10319 12839 10345 12865
rect 9311 12783 9337 12809
rect 7351 12727 7377 12753
rect 7575 12727 7601 12753
rect 8079 12727 8105 12753
rect 8247 12727 8273 12753
rect 10375 12727 10401 12753
rect 13455 12727 13481 12753
rect 13623 12727 13649 12753
rect 14071 12727 14097 12753
rect 14239 12727 14265 12753
rect 14575 12727 14601 12753
rect 7183 12671 7209 12697
rect 7239 12671 7265 12697
rect 7463 12671 7489 12697
rect 7743 12671 7769 12697
rect 7911 12671 7937 12697
rect 9255 12671 9281 12697
rect 9479 12671 9505 12697
rect 10319 12671 10345 12697
rect 13959 12671 13985 12697
rect 14183 12671 14209 12697
rect 14631 12671 14657 12697
rect 14743 12671 14769 12697
rect 7519 12615 7545 12641
rect 8079 12615 8105 12641
rect 8415 12615 8441 12641
rect 9367 12615 9393 12641
rect 11215 12615 11241 12641
rect 13567 12615 13593 12641
rect 13791 12615 13817 12641
rect 13903 12615 13929 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 11271 12447 11297 12473
rect 11663 12447 11689 12473
rect 7127 12391 7153 12417
rect 12055 12391 12081 12417
rect 13735 12391 13761 12417
rect 7519 12335 7545 12361
rect 9647 12335 9673 12361
rect 11383 12335 11409 12361
rect 11551 12335 11577 12361
rect 11775 12335 11801 12361
rect 11999 12335 12025 12361
rect 12167 12335 12193 12361
rect 13343 12335 13369 12361
rect 15023 12335 15049 12361
rect 6063 12279 6089 12305
rect 7743 12279 7769 12305
rect 10039 12279 10065 12305
rect 11103 12279 11129 12305
rect 14799 12279 14825 12305
rect 11215 12223 11241 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 9591 12055 9617 12081
rect 967 11999 993 12025
rect 4999 11999 5025 12025
rect 7071 11999 7097 12025
rect 13007 11999 13033 12025
rect 20007 11999 20033 12025
rect 2143 11943 2169 11969
rect 6455 11943 6481 11969
rect 9647 11943 9673 11969
rect 9927 11943 9953 11969
rect 10319 11943 10345 11969
rect 10767 11943 10793 11969
rect 10991 11943 11017 11969
rect 11607 11943 11633 11969
rect 13231 11943 13257 11969
rect 18831 11943 18857 11969
rect 6063 11887 6089 11913
rect 6791 11887 6817 11913
rect 6847 11887 6873 11913
rect 7967 11887 7993 11913
rect 8807 11887 8833 11913
rect 10375 11887 10401 11913
rect 11943 11887 11969 11913
rect 6679 11831 6705 11857
rect 8023 11831 8049 11857
rect 8135 11831 8161 11857
rect 8415 11831 8441 11857
rect 8639 11831 8665 11857
rect 8751 11831 8777 11857
rect 11047 11831 11073 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 6455 11663 6481 11689
rect 12055 11663 12081 11689
rect 8695 11607 8721 11633
rect 9087 11607 9113 11633
rect 9591 11607 9617 11633
rect 10207 11607 10233 11633
rect 10655 11607 10681 11633
rect 11999 11607 12025 11633
rect 12167 11607 12193 11633
rect 14183 11607 14209 11633
rect 14743 11607 14769 11633
rect 2143 11551 2169 11577
rect 6399 11551 6425 11577
rect 6511 11551 6537 11577
rect 6679 11551 6705 11577
rect 8303 11551 8329 11577
rect 8863 11551 8889 11577
rect 9143 11551 9169 11577
rect 9311 11551 9337 11577
rect 9479 11551 9505 11577
rect 10431 11551 10457 11577
rect 10543 11551 10569 11577
rect 11887 11551 11913 11577
rect 14071 11551 14097 11577
rect 14351 11551 14377 11577
rect 18831 11551 18857 11577
rect 6847 11495 6873 11521
rect 7911 11495 7937 11521
rect 10319 11495 10345 11521
rect 15807 11495 15833 11521
rect 16031 11495 16057 11521
rect 967 11439 993 11465
rect 9199 11439 9225 11465
rect 9647 11439 9673 11465
rect 20007 11439 20033 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 8415 11271 8441 11297
rect 14967 11271 14993 11297
rect 967 11215 993 11241
rect 12223 11215 12249 11241
rect 12503 11215 12529 11241
rect 14015 11215 14041 11241
rect 20007 11215 20033 11241
rect 2143 11159 2169 11185
rect 7911 11159 7937 11185
rect 8079 11159 8105 11185
rect 8247 11159 8273 11185
rect 8471 11159 8497 11185
rect 9591 11159 9617 11185
rect 9927 11159 9953 11185
rect 10039 11159 10065 11185
rect 10263 11159 10289 11185
rect 10711 11159 10737 11185
rect 12279 11159 12305 11185
rect 14127 11159 14153 11185
rect 14687 11159 14713 11185
rect 18831 11159 18857 11185
rect 8695 11103 8721 11129
rect 8807 11103 8833 11129
rect 11383 11103 11409 11129
rect 11831 11103 11857 11129
rect 12895 11103 12921 11129
rect 12951 11103 12977 11129
rect 14631 11103 14657 11129
rect 14743 11103 14769 11129
rect 8079 11047 8105 11073
rect 8415 11047 8441 11073
rect 8751 11047 8777 11073
rect 8975 11047 9001 11073
rect 9143 11047 9169 11073
rect 9311 11047 9337 11073
rect 10095 11047 10121 11073
rect 12727 11047 12753 11073
rect 13063 11047 13089 11073
rect 14295 11047 14321 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 7127 10879 7153 10905
rect 7743 10879 7769 10905
rect 11495 10879 11521 10905
rect 14407 10879 14433 10905
rect 7575 10823 7601 10849
rect 11607 10823 11633 10849
rect 6399 10767 6425 10793
rect 6567 10767 6593 10793
rect 6679 10767 6705 10793
rect 6791 10767 6817 10793
rect 6903 10767 6929 10793
rect 11327 10767 11353 10793
rect 11663 10767 11689 10793
rect 14183 10767 14209 10793
rect 4943 10711 4969 10737
rect 6007 10711 6033 10737
rect 6735 10711 6761 10737
rect 8807 10711 8833 10737
rect 12727 10711 12753 10737
rect 13791 10711 13817 10737
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 5895 10487 5921 10513
rect 10039 10487 10065 10513
rect 13567 10487 13593 10513
rect 13791 10487 13817 10513
rect 967 10431 993 10457
rect 5839 10431 5865 10457
rect 7967 10431 7993 10457
rect 9031 10431 9057 10457
rect 14519 10431 14545 10457
rect 20007 10431 20033 10457
rect 2087 10375 2113 10401
rect 7575 10375 7601 10401
rect 9367 10375 9393 10401
rect 10095 10375 10121 10401
rect 10207 10375 10233 10401
rect 10319 10375 10345 10401
rect 10655 10375 10681 10401
rect 13455 10375 13481 10401
rect 13679 10375 13705 10401
rect 14127 10375 14153 10401
rect 14799 10375 14825 10401
rect 14855 10375 14881 10401
rect 18831 10375 18857 10401
rect 9423 10319 9449 10345
rect 9759 10319 9785 10345
rect 12559 10319 12585 10345
rect 13847 10319 13873 10345
rect 14575 10319 14601 10345
rect 9591 10263 9617 10289
rect 14015 10263 14041 10289
rect 14687 10263 14713 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 8863 10095 8889 10121
rect 6175 10039 6201 10065
rect 9367 10039 9393 10065
rect 11271 10039 11297 10065
rect 2143 9983 2169 10009
rect 6287 9983 6313 10009
rect 6511 9983 6537 10009
rect 6623 9983 6649 10009
rect 6735 9983 6761 10009
rect 6847 9983 6873 10009
rect 8751 9983 8777 10009
rect 9815 9983 9841 10009
rect 10263 9983 10289 10009
rect 10655 9983 10681 10009
rect 11047 9983 11073 10009
rect 11327 9983 11353 10009
rect 11607 9983 11633 10009
rect 11831 9983 11857 10009
rect 12615 9983 12641 10009
rect 5727 9927 5753 9953
rect 6679 9927 6705 9953
rect 8415 9927 8441 9953
rect 9871 9927 9897 9953
rect 11439 9927 11465 9953
rect 14575 9927 14601 9953
rect 15471 9927 15497 9953
rect 967 9871 993 9897
rect 5783 9871 5809 9897
rect 11607 9871 11633 9897
rect 15415 9871 15441 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 6959 9703 6985 9729
rect 13511 9703 13537 9729
rect 967 9647 993 9673
rect 4831 9647 4857 9673
rect 5895 9647 5921 9673
rect 8639 9647 8665 9673
rect 9423 9647 9449 9673
rect 10431 9647 10457 9673
rect 12503 9647 12529 9673
rect 13399 9647 13425 9673
rect 16031 9647 16057 9673
rect 2143 9591 2169 9617
rect 6287 9591 6313 9617
rect 6679 9591 6705 9617
rect 6903 9591 6929 9617
rect 7071 9591 7097 9617
rect 7183 9591 7209 9617
rect 8975 9591 9001 9617
rect 9087 9591 9113 9617
rect 9647 9591 9673 9617
rect 9815 9591 9841 9617
rect 11159 9591 11185 9617
rect 11495 9591 11521 9617
rect 11663 9591 11689 9617
rect 12055 9591 12081 9617
rect 12279 9591 12305 9617
rect 12391 9591 12417 9617
rect 12559 9591 12585 9617
rect 12727 9591 12753 9617
rect 12895 9591 12921 9617
rect 13679 9591 13705 9617
rect 13791 9591 13817 9617
rect 14071 9591 14097 9617
rect 14183 9591 14209 9617
rect 14295 9591 14321 9617
rect 14575 9591 14601 9617
rect 9311 9535 9337 9561
rect 10767 9535 10793 9561
rect 10935 9535 10961 9561
rect 11271 9535 11297 9561
rect 11775 9535 11801 9561
rect 13063 9535 13089 9561
rect 13959 9535 13985 9561
rect 14967 9535 14993 9561
rect 6903 9479 6929 9505
rect 11663 9479 11689 9505
rect 14351 9479 14377 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 7743 9311 7769 9337
rect 9255 9311 9281 9337
rect 11831 9311 11857 9337
rect 12279 9311 12305 9337
rect 12223 9255 12249 9281
rect 13399 9255 13425 9281
rect 13679 9255 13705 9281
rect 5951 9199 5977 9225
rect 6343 9199 6369 9225
rect 6567 9199 6593 9225
rect 7911 9199 7937 9225
rect 9535 9199 9561 9225
rect 9759 9199 9785 9225
rect 10039 9199 10065 9225
rect 10431 9199 10457 9225
rect 10655 9199 10681 9225
rect 10879 9199 10905 9225
rect 11439 9199 11465 9225
rect 11775 9199 11801 9225
rect 12391 9199 12417 9225
rect 12951 9199 12977 9225
rect 13623 9199 13649 9225
rect 13791 9199 13817 9225
rect 14127 9199 14153 9225
rect 18943 9199 18969 9225
rect 4887 9143 4913 9169
rect 6511 9143 6537 9169
rect 6791 9143 6817 9169
rect 10263 9143 10289 9169
rect 11103 9143 11129 9169
rect 11271 9143 11297 9169
rect 11607 9143 11633 9169
rect 12839 9143 12865 9169
rect 13119 9143 13145 9169
rect 13455 9143 13481 9169
rect 14463 9143 14489 9169
rect 15527 9143 15553 9169
rect 15751 9143 15777 9169
rect 13287 9087 13313 9113
rect 20007 9087 20033 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 7743 8919 7769 8945
rect 9311 8919 9337 8945
rect 9535 8919 9561 8945
rect 9703 8919 9729 8945
rect 15079 8919 15105 8945
rect 967 8863 993 8889
rect 7407 8863 7433 8889
rect 7687 8863 7713 8889
rect 20007 8863 20033 8889
rect 2143 8807 2169 8833
rect 7239 8807 7265 8833
rect 7911 8807 7937 8833
rect 8079 8807 8105 8833
rect 8303 8807 8329 8833
rect 9367 8807 9393 8833
rect 9871 8807 9897 8833
rect 9927 8807 9953 8833
rect 10095 8807 10121 8833
rect 10767 8807 10793 8833
rect 10935 8807 10961 8833
rect 12671 8807 12697 8833
rect 12839 8807 12865 8833
rect 13007 8807 13033 8833
rect 14575 8807 14601 8833
rect 14687 8807 14713 8833
rect 14911 8807 14937 8833
rect 18831 8807 18857 8833
rect 8191 8751 8217 8777
rect 8863 8751 8889 8777
rect 9031 8751 9057 8777
rect 10655 8751 10681 8777
rect 15023 8751 15049 8777
rect 6455 8695 6481 8721
rect 7351 8695 7377 8721
rect 7911 8695 7937 8721
rect 8975 8695 9001 8721
rect 9311 8695 9337 8721
rect 9647 8695 9673 8721
rect 10767 8695 10793 8721
rect 12895 8695 12921 8721
rect 14295 8695 14321 8721
rect 14743 8695 14769 8721
rect 15079 8695 15105 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 9703 8527 9729 8553
rect 11047 8527 11073 8553
rect 11775 8527 11801 8553
rect 12839 8527 12865 8553
rect 7575 8471 7601 8497
rect 9311 8471 9337 8497
rect 10543 8471 10569 8497
rect 11383 8471 11409 8497
rect 12951 8471 12977 8497
rect 2143 8415 2169 8441
rect 7407 8415 7433 8441
rect 7743 8415 7769 8441
rect 9423 8415 9449 8441
rect 9759 8415 9785 8441
rect 10431 8415 10457 8441
rect 10879 8415 10905 8441
rect 11215 8415 11241 8441
rect 13007 8415 13033 8441
rect 13847 8415 13873 8441
rect 15527 8415 15553 8441
rect 18831 8415 18857 8441
rect 5951 8359 5977 8385
rect 7015 8359 7041 8385
rect 7631 8359 7657 8385
rect 8079 8359 8105 8385
rect 9871 8359 9897 8385
rect 11663 8359 11689 8385
rect 14239 8359 14265 8385
rect 15303 8359 15329 8385
rect 19951 8359 19977 8385
rect 967 8303 993 8329
rect 7799 8303 7825 8329
rect 9703 8303 9729 8329
rect 11831 8303 11857 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 7127 8135 7153 8161
rect 7183 8135 7209 8161
rect 7295 8135 7321 8161
rect 7351 8135 7377 8161
rect 9927 8135 9953 8161
rect 14183 8135 14209 8161
rect 7743 8079 7769 8105
rect 11327 8079 11353 8105
rect 12391 8079 12417 8105
rect 13007 8079 13033 8105
rect 20007 8079 20033 8105
rect 9255 8023 9281 8049
rect 9703 8023 9729 8049
rect 9871 8023 9897 8049
rect 12783 8023 12809 8049
rect 15023 8023 15049 8049
rect 18831 8023 18857 8049
rect 7631 7967 7657 7993
rect 7687 7967 7713 7993
rect 9367 7967 9393 7993
rect 9535 7967 9561 7993
rect 14183 7967 14209 7993
rect 14239 7967 14265 7993
rect 14519 7967 14545 7993
rect 14631 7967 14657 7993
rect 14687 7967 14713 7993
rect 15135 7911 15161 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 9983 7743 10009 7769
rect 11495 7743 11521 7769
rect 12111 7743 12137 7769
rect 14295 7743 14321 7769
rect 7015 7687 7041 7713
rect 7911 7687 7937 7713
rect 9703 7687 9729 7713
rect 10655 7687 10681 7713
rect 11775 7687 11801 7713
rect 13007 7687 13033 7713
rect 7351 7631 7377 7657
rect 9423 7631 9449 7657
rect 10151 7631 10177 7657
rect 10375 7631 10401 7657
rect 11607 7631 11633 7657
rect 11887 7631 11913 7657
rect 12671 7631 12697 7657
rect 5951 7575 5977 7601
rect 7631 7575 7657 7601
rect 9311 7575 9337 7601
rect 12167 7575 12193 7601
rect 14071 7575 14097 7601
rect 7855 7519 7881 7545
rect 11607 7519 11633 7545
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 8695 7295 8721 7321
rect 9255 7295 9281 7321
rect 10319 7295 10345 7321
rect 11495 7295 11521 7321
rect 12559 7295 12585 7321
rect 7239 7239 7265 7265
rect 8919 7239 8945 7265
rect 10711 7239 10737 7265
rect 11159 7239 11185 7265
rect 12839 7239 12865 7265
rect 7631 7183 7657 7209
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 8863 6959 8889 6985
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 12783 1807 12809 1833
rect 12279 1751 12305 1777
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8064 20600 8120 21000
rect 9408 20600 9464 21000
rect 9744 20600 9800 21000
rect 11088 20600 11144 21000
rect 11424 20600 11480 21000
rect 12096 20600 12152 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 8078 18354 8106 20600
rect 9422 19081 9450 20600
rect 9422 19055 9423 19081
rect 9449 19055 9450 19081
rect 9422 19049 9450 19055
rect 8974 19026 9002 19031
rect 8974 18979 9002 18998
rect 9310 19026 9338 19031
rect 8078 18321 8106 18326
rect 8694 18354 8722 18359
rect 8694 18307 8722 18326
rect 8190 18241 8218 18247
rect 8190 18215 8191 18241
rect 8217 18215 8218 18241
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 8190 15974 8218 18215
rect 8022 15946 8218 15974
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 8022 13538 8050 15946
rect 9310 14041 9338 18998
rect 9758 18746 9786 20600
rect 11102 19081 11130 20600
rect 11438 19138 11466 20600
rect 11438 19105 11466 19110
rect 11102 19055 11103 19081
rect 11129 19055 11130 19081
rect 11102 19049 11130 19055
rect 11886 19025 11914 19031
rect 11886 18999 11887 19025
rect 11913 18999 11914 19025
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 9758 18713 9786 18718
rect 10374 18746 10402 18751
rect 10374 18699 10402 18718
rect 9870 18634 9898 18639
rect 9310 14015 9311 14041
rect 9337 14015 9338 14041
rect 9310 14009 9338 14015
rect 9478 18633 9898 18634
rect 9478 18607 9871 18633
rect 9897 18607 9898 18633
rect 9478 18606 9898 18607
rect 9478 14042 9506 18606
rect 9870 18601 9898 18606
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 11494 14042 11522 14047
rect 9478 14041 9730 14042
rect 9478 14015 9479 14041
rect 9505 14015 9730 14041
rect 9478 14014 9730 14015
rect 8022 13510 8274 13538
rect 2086 13482 2114 13487
rect 7966 13481 7994 13487
rect 7966 13455 7967 13481
rect 7993 13455 7994 13481
rect 7966 13454 7994 13455
rect 966 13033 994 13039
rect 966 13007 967 13033
rect 993 13007 994 13033
rect 966 12810 994 13007
rect 966 12777 994 12782
rect 966 12025 994 12031
rect 966 11999 967 12025
rect 993 11999 994 12025
rect 966 11802 994 11999
rect 966 11769 994 11774
rect 966 11466 994 11471
rect 966 11419 994 11438
rect 966 11241 994 11247
rect 966 11215 967 11241
rect 993 11215 994 11241
rect 966 10794 994 11215
rect 966 10761 994 10766
rect 2086 10514 2114 13454
rect 7910 13426 7994 13454
rect 8022 13481 8050 13510
rect 8022 13455 8023 13481
rect 8049 13455 8050 13481
rect 8022 13449 8050 13455
rect 2142 13146 2170 13151
rect 2142 13099 2170 13118
rect 6062 13146 6090 13151
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 6062 12698 6090 13118
rect 6062 12305 6090 12670
rect 6846 13145 6874 13151
rect 6846 13119 6847 13145
rect 6873 13119 6874 13145
rect 6062 12279 6063 12305
rect 6089 12279 6090 12305
rect 6062 12273 6090 12279
rect 6454 12306 6482 12311
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 4998 12025 5026 12031
rect 4998 11999 4999 12025
rect 5025 11999 5026 12025
rect 2142 11970 2170 11975
rect 2142 11923 2170 11942
rect 4998 11914 5026 11999
rect 6454 11969 6482 12278
rect 6846 12306 6874 13119
rect 7182 13090 7210 13095
rect 7182 13043 7210 13062
rect 7910 12810 7938 13426
rect 8134 13425 8162 13431
rect 8134 13399 8135 13425
rect 8161 13399 8162 13425
rect 7910 12777 7938 12782
rect 7966 13090 7994 13095
rect 7350 12754 7378 12759
rect 7350 12707 7378 12726
rect 7574 12754 7602 12759
rect 7574 12707 7602 12726
rect 7182 12697 7210 12703
rect 7182 12671 7183 12697
rect 7209 12671 7210 12697
rect 7182 12642 7210 12671
rect 7238 12698 7266 12703
rect 7238 12651 7266 12670
rect 7462 12697 7490 12703
rect 7462 12671 7463 12697
rect 7489 12671 7490 12697
rect 7182 12609 7210 12614
rect 7462 12586 7490 12671
rect 7742 12698 7770 12703
rect 7910 12698 7938 12703
rect 7742 12697 7938 12698
rect 7742 12671 7743 12697
rect 7769 12671 7911 12697
rect 7937 12671 7938 12697
rect 7742 12670 7938 12671
rect 7742 12665 7770 12670
rect 7462 12553 7490 12558
rect 7518 12641 7546 12647
rect 7518 12615 7519 12641
rect 7545 12615 7546 12641
rect 7518 12474 7546 12615
rect 7126 12446 7546 12474
rect 7126 12417 7154 12446
rect 7126 12391 7127 12417
rect 7153 12391 7154 12417
rect 7126 12385 7154 12391
rect 7518 12361 7546 12367
rect 7518 12335 7519 12361
rect 7545 12335 7546 12361
rect 6846 12273 6874 12278
rect 7070 12306 7098 12311
rect 7070 12026 7098 12278
rect 7518 12306 7546 12335
rect 7518 12273 7546 12278
rect 7742 12306 7770 12311
rect 7070 12025 7154 12026
rect 7070 11999 7071 12025
rect 7097 11999 7154 12025
rect 7070 11998 7154 11999
rect 7070 11993 7098 11998
rect 6454 11943 6455 11969
rect 6481 11943 6482 11969
rect 6454 11937 6482 11943
rect 4998 11881 5026 11886
rect 6062 11914 6090 11919
rect 6790 11914 6818 11919
rect 6062 11913 6426 11914
rect 6062 11887 6063 11913
rect 6089 11887 6426 11913
rect 6062 11886 6426 11887
rect 6062 11881 6090 11886
rect 6398 11690 6426 11886
rect 6790 11867 6818 11886
rect 6846 11914 6874 11919
rect 7070 11914 7098 11919
rect 6846 11913 7070 11914
rect 6846 11887 6847 11913
rect 6873 11887 7070 11913
rect 6846 11886 7070 11887
rect 6846 11881 6874 11886
rect 6678 11857 6706 11863
rect 6678 11831 6679 11857
rect 6705 11831 6706 11857
rect 6454 11690 6482 11695
rect 6398 11689 6482 11690
rect 6398 11663 6455 11689
rect 6481 11663 6482 11689
rect 6398 11662 6482 11663
rect 6454 11657 6482 11662
rect 2142 11577 2170 11583
rect 2142 11551 2143 11577
rect 2169 11551 2170 11577
rect 2142 11522 2170 11551
rect 2142 11489 2170 11494
rect 6398 11577 6426 11583
rect 6398 11551 6399 11577
rect 6425 11551 6426 11577
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 6398 11298 6426 11551
rect 6398 11265 6426 11270
rect 6510 11577 6538 11583
rect 6510 11551 6511 11577
rect 6537 11551 6538 11577
rect 2142 11185 2170 11191
rect 2142 11159 2143 11185
rect 2169 11159 2170 11185
rect 2142 10738 2170 11159
rect 6398 10906 6426 10911
rect 6510 10906 6538 11551
rect 6678 11577 6706 11831
rect 6678 11551 6679 11577
rect 6705 11551 6706 11577
rect 6678 11545 6706 11551
rect 6846 11522 6874 11527
rect 6846 11475 6874 11494
rect 6902 10962 6930 11886
rect 7070 11881 7098 11886
rect 6846 10934 7042 10962
rect 6510 10878 6818 10906
rect 2142 10705 2170 10710
rect 4942 10794 4970 10799
rect 4942 10737 4970 10766
rect 6398 10793 6426 10878
rect 6398 10767 6399 10793
rect 6425 10767 6426 10793
rect 6398 10761 6426 10767
rect 6566 10794 6594 10799
rect 6566 10747 6594 10766
rect 6678 10793 6706 10799
rect 6678 10767 6679 10793
rect 6705 10767 6706 10793
rect 4942 10711 4943 10737
rect 4969 10711 4970 10737
rect 4942 10705 4970 10711
rect 5838 10738 5866 10743
rect 6006 10738 6034 10743
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 2086 10481 2114 10486
rect 966 10457 994 10463
rect 966 10431 967 10457
rect 993 10431 994 10457
rect 966 10122 994 10431
rect 5838 10457 5866 10710
rect 5894 10737 6034 10738
rect 5894 10711 6007 10737
rect 6033 10711 6034 10737
rect 5894 10710 6034 10711
rect 5894 10513 5922 10710
rect 6006 10705 6034 10710
rect 6678 10626 6706 10767
rect 6790 10794 6818 10878
rect 6790 10747 6818 10766
rect 6734 10738 6762 10743
rect 6734 10691 6762 10710
rect 6846 10682 6874 10934
rect 6790 10654 6874 10682
rect 6902 10850 6930 10855
rect 6902 10793 6930 10822
rect 6902 10767 6903 10793
rect 6929 10767 6930 10793
rect 6790 10626 6818 10654
rect 6678 10598 6818 10626
rect 5894 10487 5895 10513
rect 5921 10487 5922 10513
rect 5894 10481 5922 10487
rect 5838 10431 5839 10457
rect 5865 10431 5866 10457
rect 5838 10425 5866 10431
rect 966 10089 994 10094
rect 2086 10401 2114 10407
rect 2086 10375 2087 10401
rect 2113 10375 2114 10401
rect 966 9898 994 9903
rect 966 9851 994 9870
rect 2086 9898 2114 10375
rect 6902 10094 6930 10767
rect 6174 10066 6202 10071
rect 6174 10019 6202 10038
rect 6846 10066 6874 10071
rect 6902 10066 6986 10094
rect 2142 10010 2170 10015
rect 2142 9963 2170 9982
rect 6286 10010 6314 10015
rect 6510 10010 6538 10015
rect 6286 10009 6538 10010
rect 6286 9983 6287 10009
rect 6313 9983 6511 10009
rect 6537 9983 6538 10009
rect 6286 9982 6538 9983
rect 5726 9954 5754 9959
rect 5726 9907 5754 9926
rect 2086 9865 2114 9870
rect 4830 9898 4858 9903
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 966 9673 994 9679
rect 966 9647 967 9673
rect 993 9647 994 9673
rect 966 9450 994 9647
rect 4830 9673 4858 9870
rect 5782 9898 5810 9903
rect 6286 9898 6314 9982
rect 6510 9977 6538 9982
rect 6622 10009 6650 10015
rect 6622 9983 6623 10009
rect 6649 9983 6650 10009
rect 5782 9897 5922 9898
rect 5782 9871 5783 9897
rect 5809 9871 5922 9897
rect 5782 9870 5922 9871
rect 5782 9865 5810 9870
rect 4830 9647 4831 9673
rect 4857 9647 4858 9673
rect 4830 9641 4858 9647
rect 5894 9673 5922 9870
rect 6286 9865 6314 9870
rect 6622 9898 6650 9983
rect 6734 10010 6762 10015
rect 6734 9963 6762 9982
rect 6846 10009 6874 10038
rect 6846 9983 6847 10009
rect 6873 9983 6874 10009
rect 6678 9954 6706 9959
rect 6678 9907 6706 9926
rect 6622 9865 6650 9870
rect 5894 9647 5895 9673
rect 5921 9647 5922 9673
rect 5894 9641 5922 9647
rect 966 9417 994 9422
rect 2142 9617 2170 9623
rect 2142 9591 2143 9617
rect 2169 9591 2170 9617
rect 2142 9170 2170 9591
rect 6286 9618 6314 9623
rect 6678 9618 6706 9623
rect 6286 9617 6370 9618
rect 6286 9591 6287 9617
rect 6313 9591 6370 9617
rect 6286 9590 6370 9591
rect 6286 9585 6314 9590
rect 5950 9506 5978 9511
rect 5950 9225 5978 9478
rect 5950 9199 5951 9225
rect 5977 9199 5978 9225
rect 5950 9193 5978 9199
rect 6342 9225 6370 9590
rect 6342 9199 6343 9225
rect 6369 9199 6370 9225
rect 2142 9137 2170 9142
rect 4886 9170 4914 9175
rect 4886 9123 4914 9142
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 966 8889 994 8895
rect 966 8863 967 8889
rect 993 8863 994 8889
rect 966 8442 994 8863
rect 2142 8834 2170 8839
rect 2142 8787 2170 8806
rect 5950 8834 5978 8839
rect 966 8409 994 8414
rect 2142 8442 2170 8447
rect 2142 8395 2170 8414
rect 5894 8442 5922 8447
rect 966 8329 994 8335
rect 966 8303 967 8329
rect 993 8303 994 8329
rect 966 8106 994 8303
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 966 8073 994 8078
rect 5894 7994 5922 8414
rect 5950 8385 5978 8806
rect 6342 8722 6370 9199
rect 6566 9617 6706 9618
rect 6566 9591 6679 9617
rect 6705 9591 6706 9617
rect 6566 9590 6706 9591
rect 6566 9225 6594 9590
rect 6678 9585 6706 9590
rect 6846 9562 6874 9983
rect 6958 9730 6986 10066
rect 7014 9898 7042 10934
rect 7126 10906 7154 11998
rect 7742 11858 7770 12278
rect 7742 11825 7770 11830
rect 7798 11410 7826 12670
rect 7910 12665 7938 12670
rect 7966 12642 7994 13062
rect 8078 12754 8106 12759
rect 8134 12754 8162 13399
rect 8246 13089 8274 13510
rect 8302 13537 8330 13543
rect 8302 13511 8303 13537
rect 8329 13511 8330 13537
rect 8302 13482 8330 13511
rect 8638 13482 8666 13487
rect 8302 13454 8442 13482
rect 8246 13063 8247 13089
rect 8273 13063 8274 13089
rect 8246 13057 8274 13063
rect 8078 12753 8162 12754
rect 8078 12727 8079 12753
rect 8105 12727 8162 12753
rect 8078 12726 8162 12727
rect 8246 12810 8274 12815
rect 8246 12753 8274 12782
rect 8246 12727 8247 12753
rect 8273 12727 8274 12753
rect 8078 12721 8106 12726
rect 8246 12721 8274 12727
rect 8078 12642 8106 12647
rect 7966 12641 8106 12642
rect 7966 12615 8079 12641
rect 8105 12615 8106 12641
rect 7966 12614 8106 12615
rect 8078 12609 8106 12614
rect 8414 12641 8442 13454
rect 8638 13481 9058 13482
rect 8638 13455 8639 13481
rect 8665 13455 9058 13481
rect 8638 13454 9058 13455
rect 8638 13449 8666 13454
rect 8414 12615 8415 12641
rect 8441 12615 8442 12641
rect 7798 11377 7826 11382
rect 7854 12530 7882 12535
rect 7854 11914 7882 12502
rect 8414 12362 8442 12615
rect 7966 11914 7994 11919
rect 7854 11913 7994 11914
rect 7854 11887 7967 11913
rect 7993 11887 7994 11913
rect 7854 11886 7994 11887
rect 7126 10859 7154 10878
rect 7630 10906 7658 10911
rect 7574 10850 7602 10855
rect 7574 10803 7602 10822
rect 7574 10402 7602 10407
rect 7630 10402 7658 10878
rect 7742 10906 7770 10911
rect 7742 10859 7770 10878
rect 7574 10401 7658 10402
rect 7574 10375 7575 10401
rect 7601 10375 7658 10401
rect 7574 10374 7658 10375
rect 7574 10369 7602 10374
rect 7014 9865 7042 9870
rect 7182 10010 7210 10015
rect 6958 9729 7154 9730
rect 6958 9703 6959 9729
rect 6985 9703 7154 9729
rect 6958 9702 7154 9703
rect 6958 9697 6986 9702
rect 6902 9618 6930 9637
rect 6902 9585 6930 9590
rect 7070 9617 7098 9623
rect 7070 9591 7071 9617
rect 7097 9591 7098 9617
rect 6846 9529 6874 9534
rect 7070 9562 7098 9591
rect 7070 9529 7098 9534
rect 6902 9506 6930 9511
rect 6902 9459 6930 9478
rect 6566 9199 6567 9225
rect 6593 9199 6594 9225
rect 6566 9193 6594 9199
rect 6510 9170 6538 9175
rect 6510 9123 6538 9142
rect 6790 9169 6818 9175
rect 6790 9143 6791 9169
rect 6817 9143 6818 9169
rect 6454 8722 6482 8727
rect 6342 8721 6482 8722
rect 6342 8695 6455 8721
rect 6481 8695 6482 8721
rect 6342 8694 6482 8695
rect 6454 8442 6482 8694
rect 6510 8442 6538 8447
rect 6454 8414 6510 8442
rect 6510 8409 6538 8414
rect 6790 8442 6818 9143
rect 7126 9002 7154 9702
rect 7182 9617 7210 9982
rect 7182 9591 7183 9617
rect 7209 9591 7210 9617
rect 7182 9338 7210 9591
rect 7182 9305 7210 9310
rect 7742 9618 7770 9623
rect 7854 9618 7882 11886
rect 7966 11881 7994 11886
rect 8022 11857 8050 11863
rect 8022 11831 8023 11857
rect 8049 11831 8050 11857
rect 7910 11522 7938 11527
rect 8022 11522 8050 11831
rect 7910 11521 7994 11522
rect 7910 11495 7911 11521
rect 7937 11495 7994 11521
rect 7910 11494 7994 11495
rect 7910 11489 7938 11494
rect 7910 11410 7938 11415
rect 7910 11185 7938 11382
rect 7966 11242 7994 11494
rect 8022 11489 8050 11494
rect 8134 11857 8162 11863
rect 8134 11831 8135 11857
rect 8161 11831 8162 11857
rect 7966 11214 8050 11242
rect 7910 11159 7911 11185
rect 7937 11159 7938 11185
rect 7910 11153 7938 11159
rect 7966 11074 7994 11079
rect 8022 11074 8050 11214
rect 8078 11186 8106 11191
rect 8134 11186 8162 11831
rect 8358 11858 8386 11863
rect 8414 11858 8442 12334
rect 8862 13145 8890 13151
rect 8862 13119 8863 13145
rect 8889 13119 8890 13145
rect 8806 11970 8834 11975
rect 8806 11913 8834 11942
rect 8806 11887 8807 11913
rect 8833 11887 8834 11913
rect 8386 11857 8442 11858
rect 8386 11831 8415 11857
rect 8441 11831 8442 11857
rect 8386 11830 8442 11831
rect 8078 11185 8162 11186
rect 8078 11159 8079 11185
rect 8105 11159 8162 11185
rect 8078 11158 8162 11159
rect 8246 11802 8274 11807
rect 8246 11185 8274 11774
rect 8302 11578 8330 11583
rect 8358 11578 8386 11830
rect 8414 11825 8442 11830
rect 8638 11857 8666 11863
rect 8638 11831 8639 11857
rect 8665 11831 8666 11857
rect 8638 11802 8666 11831
rect 8638 11769 8666 11774
rect 8750 11857 8778 11863
rect 8750 11831 8751 11857
rect 8777 11831 8778 11857
rect 8302 11577 8386 11578
rect 8302 11551 8303 11577
rect 8329 11551 8386 11577
rect 8302 11550 8386 11551
rect 8302 11545 8330 11550
rect 8246 11159 8247 11185
rect 8273 11159 8274 11185
rect 8078 11153 8106 11158
rect 8246 11153 8274 11159
rect 8078 11074 8106 11079
rect 8022 11073 8106 11074
rect 8022 11047 8079 11073
rect 8105 11047 8106 11073
rect 8022 11046 8106 11047
rect 7966 10457 7994 11046
rect 8078 11041 8106 11046
rect 8358 10738 8386 11550
rect 8414 11746 8442 11751
rect 8414 11298 8442 11718
rect 8694 11634 8722 11639
rect 8694 11410 8722 11606
rect 8694 11377 8722 11382
rect 8414 11251 8442 11270
rect 8470 11186 8498 11191
rect 8470 11139 8498 11158
rect 8694 11186 8722 11191
rect 8750 11186 8778 11831
rect 8806 11466 8834 11887
rect 8862 11746 8890 13119
rect 9030 13090 9058 13454
rect 9422 13258 9450 13263
rect 9198 13257 9450 13258
rect 9198 13231 9423 13257
rect 9449 13231 9450 13257
rect 9198 13230 9450 13231
rect 9086 13202 9114 13207
rect 9086 13155 9114 13174
rect 9142 13202 9170 13207
rect 9198 13202 9226 13230
rect 9422 13225 9450 13230
rect 9142 13201 9226 13202
rect 9142 13175 9143 13201
rect 9169 13175 9226 13201
rect 9142 13174 9226 13175
rect 9478 13201 9506 14014
rect 9702 13593 9730 14014
rect 11382 14014 11494 14042
rect 11214 13986 11242 13991
rect 10934 13985 11242 13986
rect 10934 13959 11215 13985
rect 11241 13959 11242 13985
rect 10934 13958 11242 13959
rect 10486 13818 10514 13823
rect 9702 13567 9703 13593
rect 9729 13567 9730 13593
rect 9702 13561 9730 13567
rect 10430 13790 10486 13818
rect 9926 13426 9954 13431
rect 9478 13175 9479 13201
rect 9505 13175 9506 13201
rect 9142 13169 9170 13174
rect 9478 13169 9506 13175
rect 9814 13425 9954 13426
rect 9814 13399 9927 13425
rect 9953 13399 9954 13425
rect 9814 13398 9954 13399
rect 9254 13145 9282 13151
rect 9254 13119 9255 13145
rect 9281 13119 9282 13145
rect 9086 13090 9114 13095
rect 9030 13089 9114 13090
rect 9030 13063 9087 13089
rect 9113 13063 9114 13089
rect 9030 13062 9114 13063
rect 9086 13057 9114 13062
rect 9254 12697 9282 13119
rect 9366 13146 9394 13151
rect 9310 12810 9338 12815
rect 9310 12763 9338 12782
rect 9254 12671 9255 12697
rect 9281 12671 9282 12697
rect 9198 11970 9226 11975
rect 9254 11970 9282 12671
rect 9366 12754 9394 13118
rect 9366 12641 9394 12726
rect 9814 13146 9842 13398
rect 9926 13393 9954 13398
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9982 13146 10010 13151
rect 9814 13145 10010 13146
rect 9814 13119 9983 13145
rect 10009 13119 10010 13145
rect 9814 13118 10010 13119
rect 9814 13089 9842 13118
rect 9982 13113 10010 13118
rect 9814 13063 9815 13089
rect 9841 13063 9842 13089
rect 9478 12698 9506 12703
rect 9478 12651 9506 12670
rect 9366 12615 9367 12641
rect 9393 12615 9394 12641
rect 9366 12138 9394 12615
rect 9814 12642 9842 13063
rect 10374 13089 10402 13095
rect 10374 13063 10375 13089
rect 10401 13063 10402 13089
rect 10318 12866 10346 12871
rect 10374 12866 10402 13063
rect 10318 12865 10402 12866
rect 10318 12839 10319 12865
rect 10345 12839 10402 12865
rect 10318 12838 10402 12839
rect 10318 12833 10346 12838
rect 10318 12754 10346 12759
rect 9590 12418 9618 12423
rect 9366 12110 9562 12138
rect 9226 11942 9282 11970
rect 9198 11937 9226 11942
rect 8862 11713 8890 11718
rect 9086 11633 9114 11639
rect 9086 11607 9087 11633
rect 9113 11607 9114 11633
rect 8862 11578 8890 11583
rect 9086 11578 9114 11607
rect 8862 11577 8946 11578
rect 8862 11551 8863 11577
rect 8889 11551 8946 11577
rect 8862 11550 8946 11551
rect 8862 11545 8890 11550
rect 8806 11438 8890 11466
rect 8750 11158 8834 11186
rect 8694 11129 8722 11158
rect 8694 11103 8695 11129
rect 8721 11103 8722 11129
rect 8694 11097 8722 11103
rect 8806 11129 8834 11158
rect 8806 11103 8807 11129
rect 8833 11103 8834 11129
rect 8414 11073 8442 11079
rect 8414 11047 8415 11073
rect 8441 11047 8442 11073
rect 8414 10850 8442 11047
rect 8750 11074 8778 11079
rect 8750 11027 8778 11046
rect 8806 10850 8834 11103
rect 8414 10817 8442 10822
rect 8638 10822 8834 10850
rect 8414 10738 8442 10743
rect 8358 10710 8414 10738
rect 7966 10431 7967 10457
rect 7993 10431 7994 10457
rect 7966 10425 7994 10431
rect 8414 9954 8442 10710
rect 7770 9590 7882 9618
rect 8358 9953 8442 9954
rect 8358 9927 8415 9953
rect 8441 9927 8442 9953
rect 8358 9926 8442 9927
rect 7742 9337 7770 9590
rect 7742 9311 7743 9337
rect 7769 9311 7770 9337
rect 7742 9305 7770 9311
rect 7966 9338 7994 9343
rect 7910 9225 7938 9231
rect 7910 9199 7911 9225
rect 7937 9199 7938 9225
rect 7126 8974 7210 9002
rect 7014 8498 7042 8503
rect 6790 8409 6818 8414
rect 6958 8470 7014 8498
rect 5950 8359 5951 8385
rect 5977 8359 5978 8385
rect 5950 8353 5978 8359
rect 5894 7602 5922 7966
rect 6958 7714 6986 8470
rect 7014 8465 7042 8470
rect 7014 8385 7042 8391
rect 7014 8359 7015 8385
rect 7041 8359 7042 8385
rect 7014 8162 7042 8359
rect 7182 8386 7210 8974
rect 7742 8946 7770 8951
rect 7910 8946 7938 9199
rect 7742 8945 7938 8946
rect 7742 8919 7743 8945
rect 7769 8919 7938 8945
rect 7742 8918 7938 8919
rect 7742 8913 7770 8918
rect 7406 8890 7434 8895
rect 7406 8843 7434 8862
rect 7686 8890 7714 8895
rect 7238 8834 7266 8839
rect 7238 8787 7266 8806
rect 7350 8721 7378 8727
rect 7350 8695 7351 8721
rect 7377 8695 7378 8721
rect 7126 8162 7154 8167
rect 7014 8161 7154 8162
rect 7014 8135 7127 8161
rect 7153 8135 7154 8161
rect 7014 8134 7154 8135
rect 7126 8129 7154 8134
rect 7182 8161 7210 8358
rect 7182 8135 7183 8161
rect 7209 8135 7210 8161
rect 7182 8129 7210 8135
rect 7294 8610 7322 8615
rect 7294 8161 7322 8582
rect 7294 8135 7295 8161
rect 7321 8135 7322 8161
rect 7294 8129 7322 8135
rect 7350 8161 7378 8695
rect 7574 8498 7602 8503
rect 7574 8451 7602 8470
rect 7350 8135 7351 8161
rect 7377 8135 7378 8161
rect 7350 8129 7378 8135
rect 7406 8442 7434 8447
rect 7014 7714 7042 7719
rect 6958 7713 7042 7714
rect 6958 7687 7015 7713
rect 7041 7687 7042 7713
rect 6958 7686 7042 7687
rect 7014 7681 7042 7686
rect 7350 7658 7378 7663
rect 7406 7658 7434 8414
rect 7630 8386 7658 8391
rect 7630 8339 7658 8358
rect 7686 8274 7714 8862
rect 7910 8833 7938 8918
rect 7910 8807 7911 8833
rect 7937 8807 7938 8833
rect 7910 8801 7938 8807
rect 7910 8722 7938 8727
rect 7742 8721 7938 8722
rect 7742 8695 7911 8721
rect 7937 8695 7938 8721
rect 7742 8694 7938 8695
rect 7742 8441 7770 8694
rect 7910 8689 7938 8694
rect 7742 8415 7743 8441
rect 7769 8415 7770 8441
rect 7742 8409 7770 8415
rect 7798 8329 7826 8335
rect 7798 8303 7799 8329
rect 7825 8303 7826 8329
rect 7686 8246 7770 8274
rect 7742 8105 7770 8246
rect 7742 8079 7743 8105
rect 7769 8079 7770 8105
rect 7742 8073 7770 8079
rect 7630 7994 7658 7999
rect 7630 7947 7658 7966
rect 7686 7994 7714 7999
rect 7798 7994 7826 8303
rect 7686 7993 7826 7994
rect 7686 7967 7687 7993
rect 7713 7967 7826 7993
rect 7686 7966 7826 7967
rect 7686 7961 7714 7966
rect 7910 7714 7938 7719
rect 7966 7714 7994 9310
rect 8078 8833 8106 8839
rect 8078 8807 8079 8833
rect 8105 8807 8106 8833
rect 8078 8554 8106 8807
rect 8302 8834 8330 8839
rect 8302 8787 8330 8806
rect 8190 8778 8218 8783
rect 8190 8731 8218 8750
rect 8078 8521 8106 8526
rect 7938 7686 7994 7714
rect 8078 8386 8106 8391
rect 8358 8386 8386 9926
rect 8414 9921 8442 9926
rect 8638 9673 8666 10822
rect 8806 10738 8834 10743
rect 8806 10691 8834 10710
rect 8862 10121 8890 11438
rect 8918 10906 8946 11550
rect 9086 11545 9114 11550
rect 9142 11578 9170 11583
rect 9310 11578 9338 11583
rect 9142 11577 9338 11578
rect 9142 11551 9143 11577
rect 9169 11551 9311 11577
rect 9337 11551 9338 11577
rect 9142 11550 9338 11551
rect 9142 11186 9170 11550
rect 9310 11545 9338 11550
rect 9478 11577 9506 11583
rect 9478 11551 9479 11577
rect 9505 11551 9506 11577
rect 9478 11522 9506 11551
rect 9478 11489 9506 11494
rect 9198 11465 9226 11471
rect 9198 11439 9199 11465
rect 9225 11439 9226 11465
rect 9198 11410 9226 11439
rect 9198 11377 9226 11382
rect 9142 11153 9170 11158
rect 8918 10514 8946 10878
rect 8918 10481 8946 10486
rect 8974 11073 9002 11079
rect 8974 11047 8975 11073
rect 9001 11047 9002 11073
rect 8974 10850 9002 11047
rect 8974 10178 9002 10822
rect 9142 11073 9170 11079
rect 9142 11047 9143 11073
rect 9169 11047 9170 11073
rect 9030 10570 9058 10575
rect 9030 10457 9058 10542
rect 9030 10431 9031 10457
rect 9057 10431 9058 10457
rect 9030 10425 9058 10431
rect 9030 10178 9058 10183
rect 8974 10150 9030 10178
rect 8862 10095 8863 10121
rect 8889 10095 8890 10121
rect 8862 10089 8890 10095
rect 8638 9647 8639 9673
rect 8665 9647 8666 9673
rect 8638 9641 8666 9647
rect 8750 10009 8778 10015
rect 8750 9983 8751 10009
rect 8777 9983 8778 10009
rect 8750 9562 8778 9983
rect 8974 9674 9002 9679
rect 8974 9617 9002 9646
rect 8974 9591 8975 9617
rect 9001 9591 9002 9617
rect 8974 9585 9002 9591
rect 8750 8890 8778 9534
rect 8750 8857 8778 8862
rect 8862 8778 8890 8783
rect 8862 8731 8890 8750
rect 9030 8778 9058 10150
rect 9142 9842 9170 11047
rect 9310 11073 9338 11079
rect 9310 11047 9311 11073
rect 9337 11047 9338 11073
rect 9310 10570 9338 11047
rect 9338 10542 9506 10570
rect 9310 10537 9338 10542
rect 9366 10401 9394 10407
rect 9366 10375 9367 10401
rect 9393 10375 9394 10401
rect 9366 10346 9394 10375
rect 9142 9809 9170 9814
rect 9254 10318 9394 10346
rect 9422 10345 9450 10351
rect 9422 10319 9423 10345
rect 9449 10319 9450 10345
rect 9254 10066 9282 10318
rect 9366 10178 9394 10183
rect 9422 10178 9450 10319
rect 9394 10150 9450 10178
rect 9366 10145 9394 10150
rect 9478 10122 9506 10542
rect 9534 10290 9562 12110
rect 9590 12081 9618 12390
rect 9646 12362 9674 12367
rect 9814 12362 9842 12614
rect 10262 12698 10290 12703
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9674 12334 9842 12362
rect 9646 12315 9674 12334
rect 9590 12055 9591 12081
rect 9617 12055 9618 12081
rect 9590 12049 9618 12055
rect 10038 12305 10066 12311
rect 10038 12279 10039 12305
rect 10065 12279 10066 12305
rect 9646 11970 9674 11975
rect 9926 11970 9954 11975
rect 9646 11923 9674 11942
rect 9814 11969 9954 11970
rect 9814 11943 9927 11969
rect 9953 11943 9954 11969
rect 9814 11942 9954 11943
rect 9590 11633 9618 11639
rect 9590 11607 9591 11633
rect 9617 11607 9618 11633
rect 9590 11354 9618 11607
rect 9646 11466 9674 11471
rect 9646 11419 9674 11438
rect 9590 11326 9786 11354
rect 9590 11186 9618 11191
rect 9590 11185 9730 11186
rect 9590 11159 9591 11185
rect 9617 11159 9730 11185
rect 9590 11158 9730 11159
rect 9590 11153 9618 11158
rect 9590 10290 9618 10295
rect 9534 10289 9618 10290
rect 9534 10263 9591 10289
rect 9617 10263 9618 10289
rect 9534 10262 9618 10263
rect 9590 10257 9618 10262
rect 9422 10094 9506 10122
rect 9254 9730 9282 10038
rect 9366 10065 9394 10071
rect 9366 10039 9367 10065
rect 9393 10039 9394 10065
rect 9366 9786 9394 10039
rect 9366 9753 9394 9758
rect 9254 9697 9282 9702
rect 9422 9674 9450 10094
rect 9366 9673 9450 9674
rect 9366 9647 9423 9673
rect 9449 9647 9450 9673
rect 9366 9646 9450 9647
rect 9086 9618 9114 9623
rect 9198 9618 9226 9623
rect 9086 9617 9198 9618
rect 9086 9591 9087 9617
rect 9113 9591 9198 9617
rect 9086 9590 9198 9591
rect 9086 9585 9114 9590
rect 9198 9226 9226 9590
rect 9310 9562 9338 9567
rect 9310 9515 9338 9534
rect 9366 9450 9394 9646
rect 9422 9641 9450 9646
rect 9534 9954 9562 9959
rect 9254 9422 9506 9450
rect 9254 9337 9282 9422
rect 9254 9311 9255 9337
rect 9281 9311 9282 9337
rect 9254 9305 9282 9311
rect 9366 9226 9394 9231
rect 9198 9198 9338 9226
rect 9310 8945 9338 9198
rect 9310 8919 9311 8945
rect 9337 8919 9338 8945
rect 9310 8913 9338 8919
rect 9366 8946 9394 9198
rect 9478 9058 9506 9422
rect 9534 9225 9562 9926
rect 9702 9674 9730 11158
rect 9758 10794 9786 11326
rect 9758 10761 9786 10766
rect 9814 11298 9842 11942
rect 9926 11937 9954 11942
rect 10038 11858 10066 12279
rect 10262 11970 10290 12670
rect 10318 12697 10346 12726
rect 10374 12754 10402 12759
rect 10430 12754 10458 13790
rect 10486 13785 10514 13790
rect 10878 13538 10906 13543
rect 10878 13491 10906 13510
rect 10374 12753 10458 12754
rect 10374 12727 10375 12753
rect 10401 12727 10458 12753
rect 10374 12726 10458 12727
rect 10374 12721 10402 12726
rect 10318 12671 10319 12697
rect 10345 12671 10346 12697
rect 10318 12665 10346 12671
rect 10934 12698 10962 13958
rect 11214 13953 11242 13958
rect 11270 13929 11298 13935
rect 11270 13903 11271 13929
rect 11297 13903 11298 13929
rect 11214 13817 11242 13823
rect 11214 13791 11215 13817
rect 11241 13791 11242 13817
rect 11214 13593 11242 13791
rect 11270 13762 11298 13903
rect 11270 13729 11298 13734
rect 11214 13567 11215 13593
rect 11241 13567 11242 13593
rect 11214 13561 11242 13567
rect 11382 13454 11410 14014
rect 11494 13995 11522 14014
rect 11550 13930 11578 13935
rect 11550 13929 11746 13930
rect 11550 13903 11551 13929
rect 11577 13903 11746 13929
rect 11550 13902 11746 13903
rect 11550 13897 11578 13902
rect 11494 13818 11522 13823
rect 11494 13771 11522 13790
rect 11550 13762 11578 13767
rect 11578 13734 11690 13762
rect 11550 13729 11578 13734
rect 11382 13426 11466 13454
rect 11438 13089 11466 13426
rect 11662 13257 11690 13734
rect 11662 13231 11663 13257
rect 11689 13231 11690 13257
rect 11662 13225 11690 13231
rect 11718 13146 11746 13902
rect 11774 13594 11802 13599
rect 11774 13257 11802 13566
rect 11774 13231 11775 13257
rect 11801 13231 11802 13257
rect 11774 13225 11802 13231
rect 11830 13146 11858 13151
rect 11718 13145 11858 13146
rect 11718 13119 11831 13145
rect 11857 13119 11858 13145
rect 11718 13118 11858 13119
rect 11438 13063 11439 13089
rect 11465 13063 11466 13089
rect 11438 13057 11466 13063
rect 11830 12754 11858 13118
rect 10934 12665 10962 12670
rect 11662 12726 11830 12754
rect 11214 12642 11242 12647
rect 11214 12595 11242 12614
rect 11270 12474 11298 12479
rect 11102 12446 11270 12474
rect 11102 12305 11130 12446
rect 11270 12427 11298 12446
rect 11662 12473 11690 12726
rect 11830 12721 11858 12726
rect 11662 12447 11663 12473
rect 11689 12447 11690 12473
rect 11662 12441 11690 12447
rect 11886 12474 11914 18999
rect 12110 18746 12138 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 12110 18713 12138 18718
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 12278 14042 12306 18999
rect 13118 18746 13146 18751
rect 13118 18699 13146 18718
rect 12278 14009 12306 14014
rect 12614 18633 12642 18639
rect 12614 18607 12615 18633
rect 12641 18607 12642 18633
rect 12278 13594 12306 13599
rect 12278 13547 12306 13566
rect 12614 13594 12642 18607
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 12614 13561 12642 13566
rect 20006 13593 20034 13599
rect 20006 13567 20007 13593
rect 20033 13567 20034 13593
rect 12502 13538 12530 13543
rect 12502 13491 12530 13510
rect 13006 13538 13034 13543
rect 13006 13454 13034 13510
rect 18942 13537 18970 13543
rect 18942 13511 18943 13537
rect 18969 13511 18970 13537
rect 13006 13426 13090 13454
rect 11886 12441 11914 12446
rect 13062 13145 13090 13426
rect 13062 13119 13063 13145
rect 13089 13119 13090 13145
rect 12054 12418 12082 12423
rect 12054 12371 12082 12390
rect 13006 12418 13034 12423
rect 11382 12362 11410 12367
rect 11102 12279 11103 12305
rect 11129 12279 11130 12305
rect 11102 12273 11130 12279
rect 11270 12361 11410 12362
rect 11270 12335 11383 12361
rect 11409 12335 11410 12361
rect 11270 12334 11410 12335
rect 11214 12249 11242 12255
rect 11214 12223 11215 12249
rect 11241 12223 11242 12249
rect 10318 11970 10346 11975
rect 10262 11969 10346 11970
rect 10262 11943 10319 11969
rect 10345 11943 10346 11969
rect 10262 11942 10346 11943
rect 10038 11830 10122 11858
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9758 10345 9786 10351
rect 9758 10319 9759 10345
rect 9785 10319 9786 10345
rect 9758 10010 9786 10319
rect 9814 10122 9842 11270
rect 9926 11634 9954 11639
rect 9926 11185 9954 11606
rect 9926 11159 9927 11185
rect 9953 11159 9954 11185
rect 9926 11153 9954 11159
rect 10038 11466 10066 11471
rect 10038 11185 10066 11438
rect 10038 11159 10039 11185
rect 10065 11159 10066 11185
rect 10038 11153 10066 11159
rect 10094 11073 10122 11830
rect 10262 11802 10290 11807
rect 10206 11690 10234 11695
rect 10206 11633 10234 11662
rect 10206 11607 10207 11633
rect 10233 11607 10234 11633
rect 10206 11410 10234 11607
rect 10206 11377 10234 11382
rect 10262 11185 10290 11774
rect 10318 11521 10346 11942
rect 10766 11969 10794 11975
rect 10766 11943 10767 11969
rect 10793 11943 10794 11969
rect 10318 11495 10319 11521
rect 10345 11495 10346 11521
rect 10318 11489 10346 11495
rect 10374 11913 10402 11919
rect 10374 11887 10375 11913
rect 10401 11887 10402 11913
rect 10374 11354 10402 11887
rect 10654 11634 10682 11639
rect 10374 11321 10402 11326
rect 10430 11578 10458 11583
rect 10262 11159 10263 11185
rect 10289 11159 10290 11185
rect 10262 11153 10290 11159
rect 10430 11186 10458 11550
rect 10430 11153 10458 11158
rect 10542 11577 10570 11583
rect 10542 11551 10543 11577
rect 10569 11551 10570 11577
rect 10542 11522 10570 11551
rect 10094 11047 10095 11073
rect 10121 11047 10122 11073
rect 10094 11041 10122 11047
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 10094 10962 10122 10967
rect 10038 10514 10066 10519
rect 10038 10467 10066 10486
rect 10094 10401 10122 10934
rect 10542 10962 10570 11494
rect 10542 10929 10570 10934
rect 10654 10962 10682 11606
rect 10710 11186 10738 11191
rect 10766 11186 10794 11943
rect 10990 11969 11018 11975
rect 10990 11943 10991 11969
rect 11017 11943 11018 11969
rect 10990 11634 11018 11943
rect 10990 11601 11018 11606
rect 11046 11857 11074 11863
rect 11046 11831 11047 11857
rect 11073 11831 11074 11857
rect 10710 11185 11018 11186
rect 10710 11159 10711 11185
rect 10737 11159 11018 11185
rect 10710 11158 11018 11159
rect 10710 11153 10738 11158
rect 10654 10929 10682 10934
rect 10934 10962 10962 10967
rect 10094 10375 10095 10401
rect 10121 10375 10122 10401
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9814 10094 9898 10122
rect 9758 9977 9786 9982
rect 9814 10009 9842 10015
rect 9814 9983 9815 10009
rect 9841 9983 9842 10009
rect 9814 9954 9842 9983
rect 9814 9921 9842 9926
rect 9870 9953 9898 10094
rect 9870 9927 9871 9953
rect 9897 9927 9898 9953
rect 9870 9921 9898 9927
rect 9814 9842 9842 9847
rect 9534 9199 9535 9225
rect 9561 9199 9562 9225
rect 9534 9114 9562 9199
rect 9646 9617 9674 9623
rect 9646 9591 9647 9617
rect 9673 9591 9674 9617
rect 9646 9226 9674 9591
rect 9702 9338 9730 9646
rect 9702 9305 9730 9310
rect 9758 9814 9814 9842
rect 9646 9193 9674 9198
rect 9758 9225 9786 9814
rect 9814 9809 9842 9814
rect 9758 9199 9759 9225
rect 9785 9199 9786 9225
rect 9758 9193 9786 9199
rect 9814 9617 9842 9623
rect 9814 9591 9815 9617
rect 9841 9591 9842 9617
rect 9534 9086 9786 9114
rect 9478 9030 9562 9058
rect 9366 8833 9394 8918
rect 9534 8945 9562 9030
rect 9534 8919 9535 8945
rect 9561 8919 9562 8945
rect 9534 8913 9562 8919
rect 9702 8946 9730 8951
rect 9702 8899 9730 8918
rect 9366 8807 9367 8833
rect 9393 8807 9394 8833
rect 9366 8801 9394 8807
rect 9030 8731 9058 8750
rect 8974 8722 9002 8727
rect 9254 8722 9282 8727
rect 8974 8675 9002 8694
rect 9198 8694 9254 8722
rect 8078 8385 8386 8386
rect 8078 8359 8079 8385
rect 8105 8359 8386 8385
rect 8078 8358 8386 8359
rect 7910 7667 7938 7686
rect 7350 7657 7434 7658
rect 7350 7631 7351 7657
rect 7377 7631 7434 7657
rect 7350 7630 7434 7631
rect 5950 7602 5978 7607
rect 5894 7601 5978 7602
rect 5894 7575 5951 7601
rect 5977 7575 5978 7601
rect 5894 7574 5978 7575
rect 5950 7569 5978 7574
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 7238 7266 7266 7271
rect 7350 7266 7378 7630
rect 7630 7601 7658 7607
rect 7630 7575 7631 7601
rect 7657 7575 7658 7601
rect 7630 7574 7658 7575
rect 7630 7546 7714 7574
rect 7238 7265 7350 7266
rect 7238 7239 7239 7265
rect 7265 7239 7350 7265
rect 7238 7238 7350 7239
rect 7238 7233 7266 7238
rect 7350 7233 7378 7238
rect 7686 7266 7714 7546
rect 7686 7233 7714 7238
rect 7854 7545 7882 7551
rect 7854 7519 7855 7545
rect 7881 7519 7882 7545
rect 7630 7209 7658 7215
rect 7630 7183 7631 7209
rect 7657 7183 7658 7209
rect 7630 7154 7658 7183
rect 7854 7154 7882 7519
rect 8078 7266 8106 8358
rect 8694 7602 8722 7607
rect 8694 7321 8722 7574
rect 8694 7295 8695 7321
rect 8721 7295 8722 7321
rect 8694 7289 8722 7295
rect 9198 7322 9226 8694
rect 9254 8689 9282 8694
rect 9310 8722 9338 8727
rect 9310 8721 9450 8722
rect 9310 8695 9311 8721
rect 9337 8695 9450 8721
rect 9310 8694 9450 8695
rect 9310 8689 9338 8694
rect 9310 8498 9338 8503
rect 9310 8451 9338 8470
rect 9422 8442 9450 8694
rect 9646 8721 9674 8727
rect 9646 8695 9647 8721
rect 9673 8695 9674 8721
rect 9646 8610 9674 8695
rect 9646 8577 9674 8582
rect 9702 8554 9730 8559
rect 9702 8507 9730 8526
rect 9422 8395 9450 8414
rect 9758 8441 9786 9086
rect 9814 8610 9842 9591
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9926 9338 9954 9343
rect 9926 9170 9954 9310
rect 10038 9226 10066 9231
rect 10038 9179 10066 9198
rect 9870 8834 9898 8839
rect 9870 8787 9898 8806
rect 9926 8833 9954 9142
rect 10094 9114 10122 10375
rect 10206 10401 10234 10407
rect 10206 10375 10207 10401
rect 10233 10375 10234 10401
rect 10206 10066 10234 10375
rect 10318 10401 10346 10407
rect 10318 10375 10319 10401
rect 10345 10375 10346 10401
rect 10262 10066 10290 10071
rect 10206 10038 10262 10066
rect 10094 9081 10122 9086
rect 10150 10010 10178 10015
rect 9926 8807 9927 8833
rect 9953 8807 9954 8833
rect 9926 8801 9954 8807
rect 10094 8833 10122 8839
rect 10094 8807 10095 8833
rect 10121 8807 10122 8833
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9814 8577 9842 8582
rect 9758 8415 9759 8441
rect 9785 8415 9786 8441
rect 9758 8409 9786 8415
rect 9870 8386 9898 8391
rect 9870 8339 9898 8358
rect 10094 8386 10122 8807
rect 10094 8353 10122 8358
rect 10150 8722 10178 9982
rect 10262 10009 10290 10038
rect 10262 9983 10263 10009
rect 10289 9983 10290 10009
rect 10262 9977 10290 9983
rect 10318 9954 10346 10375
rect 10318 9921 10346 9926
rect 10430 10402 10458 10407
rect 10430 9673 10458 10374
rect 10654 10402 10682 10407
rect 10654 10355 10682 10374
rect 10654 10010 10682 10015
rect 10654 9963 10682 9982
rect 10430 9647 10431 9673
rect 10457 9647 10458 9673
rect 10430 9641 10458 9647
rect 10598 9730 10626 9735
rect 10262 9450 10290 9455
rect 10262 9169 10290 9422
rect 10262 9143 10263 9169
rect 10289 9143 10290 9169
rect 10262 9137 10290 9143
rect 10430 9225 10458 9231
rect 10430 9199 10431 9225
rect 10457 9199 10458 9225
rect 10430 9170 10458 9199
rect 10598 9226 10626 9702
rect 10766 9561 10794 9567
rect 10766 9535 10767 9561
rect 10793 9535 10794 9561
rect 10654 9226 10682 9231
rect 10598 9225 10682 9226
rect 10598 9199 10655 9225
rect 10681 9199 10682 9225
rect 10598 9198 10682 9199
rect 10654 9193 10682 9198
rect 10430 9137 10458 9142
rect 10766 9114 10794 9535
rect 10934 9561 10962 10934
rect 10990 10010 11018 11158
rect 11046 11018 11074 11831
rect 11214 11802 11242 12223
rect 11214 11769 11242 11774
rect 11046 10985 11074 10990
rect 11270 10178 11298 12334
rect 11382 12329 11410 12334
rect 11550 12361 11578 12367
rect 11550 12335 11551 12361
rect 11577 12335 11578 12361
rect 11550 11634 11578 12335
rect 11774 12361 11802 12367
rect 11998 12362 12026 12367
rect 11774 12335 11775 12361
rect 11801 12335 11802 12361
rect 11606 11970 11634 11975
rect 11606 11923 11634 11942
rect 11774 11914 11802 12335
rect 11774 11881 11802 11886
rect 11886 12361 12026 12362
rect 11886 12335 11999 12361
rect 12025 12335 12026 12361
rect 11886 12334 12026 12335
rect 11886 11690 11914 12334
rect 11998 12329 12026 12334
rect 12166 12361 12194 12367
rect 12166 12335 12167 12361
rect 12193 12335 12194 12361
rect 11942 11914 11970 11919
rect 11942 11913 12082 11914
rect 11942 11887 11943 11913
rect 11969 11887 12082 11913
rect 11942 11886 12082 11887
rect 11942 11881 11970 11886
rect 11914 11662 11970 11690
rect 11886 11657 11914 11662
rect 11382 11129 11410 11135
rect 11382 11103 11383 11129
rect 11409 11103 11410 11129
rect 11382 10962 11410 11103
rect 11382 10929 11410 10934
rect 11494 10906 11522 10911
rect 11550 10906 11578 11606
rect 11886 11577 11914 11583
rect 11886 11551 11887 11577
rect 11913 11551 11914 11577
rect 11494 10905 11578 10906
rect 11494 10879 11495 10905
rect 11521 10879 11578 10905
rect 11494 10878 11578 10879
rect 11606 11158 11858 11186
rect 11494 10873 11522 10878
rect 11606 10849 11634 11158
rect 11830 11129 11858 11158
rect 11830 11103 11831 11129
rect 11857 11103 11858 11129
rect 11830 11097 11858 11103
rect 11606 10823 11607 10849
rect 11633 10823 11634 10849
rect 11326 10793 11354 10799
rect 11326 10767 11327 10793
rect 11353 10767 11354 10793
rect 11326 10346 11354 10767
rect 11326 10313 11354 10318
rect 11214 10150 11298 10178
rect 11046 10010 11074 10015
rect 10990 10009 11074 10010
rect 10990 9983 11047 10009
rect 11073 9983 11074 10009
rect 10990 9982 11074 9983
rect 10990 9842 11018 9982
rect 11046 9977 11074 9982
rect 10990 9809 11018 9814
rect 10934 9535 10935 9561
rect 10961 9535 10962 9561
rect 10934 9338 10962 9535
rect 10766 9081 10794 9086
rect 10822 9310 10962 9338
rect 11158 9617 11186 9623
rect 11158 9591 11159 9617
rect 11185 9591 11186 9617
rect 10766 8890 10794 8895
rect 10766 8833 10794 8862
rect 10766 8807 10767 8833
rect 10793 8807 10794 8833
rect 10766 8801 10794 8807
rect 10654 8778 10682 8783
rect 10654 8731 10682 8750
rect 9702 8329 9730 8335
rect 9702 8303 9703 8329
rect 9729 8303 9730 8329
rect 9534 8274 9562 8279
rect 9254 8050 9282 8055
rect 9254 8049 9338 8050
rect 9254 8023 9255 8049
rect 9281 8023 9338 8049
rect 9254 8022 9338 8023
rect 9254 8017 9282 8022
rect 9310 7602 9338 8022
rect 9366 7994 9394 7999
rect 9366 7947 9394 7966
rect 9534 7993 9562 8246
rect 9534 7967 9535 7993
rect 9561 7967 9562 7993
rect 9534 7714 9562 7967
rect 9534 7681 9562 7686
rect 9702 8049 9730 8303
rect 10150 8274 10178 8694
rect 10766 8722 10794 8727
rect 10766 8675 10794 8694
rect 10430 8554 10458 8559
rect 10430 8441 10458 8526
rect 10430 8415 10431 8441
rect 10457 8415 10458 8441
rect 10430 8409 10458 8415
rect 10542 8497 10570 8503
rect 10542 8471 10543 8497
rect 10569 8471 10570 8497
rect 10542 8386 10570 8471
rect 10542 8353 10570 8358
rect 9926 8246 10178 8274
rect 9926 8161 9954 8246
rect 9926 8135 9927 8161
rect 9953 8135 9954 8161
rect 9926 8129 9954 8135
rect 9870 8050 9898 8055
rect 9702 8023 9703 8049
rect 9729 8023 9730 8049
rect 9702 7713 9730 8023
rect 9814 8022 9870 8050
rect 9814 7770 9842 8022
rect 9870 8003 9898 8022
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9982 7770 10010 7775
rect 9814 7769 10010 7770
rect 9814 7743 9983 7769
rect 10009 7743 10010 7769
rect 9814 7742 10010 7743
rect 9982 7737 10010 7742
rect 9702 7687 9703 7713
rect 9729 7687 9730 7713
rect 9702 7681 9730 7687
rect 10654 7714 10682 7719
rect 10822 7714 10850 9310
rect 11158 9282 11186 9591
rect 11046 9254 11186 9282
rect 10878 9226 10906 9231
rect 11046 9226 11074 9254
rect 10878 9225 11074 9226
rect 10878 9199 10879 9225
rect 10905 9199 11074 9225
rect 10878 9198 11074 9199
rect 10878 8946 10906 9198
rect 11102 9170 11130 9175
rect 11102 9123 11130 9142
rect 11214 9058 11242 10150
rect 11270 10066 11298 10071
rect 11270 10019 11298 10038
rect 11326 10009 11354 10015
rect 11606 10010 11634 10823
rect 11326 9983 11327 10009
rect 11353 9983 11354 10009
rect 11326 9954 11354 9983
rect 11550 10009 11634 10010
rect 11550 9983 11607 10009
rect 11633 9983 11634 10009
rect 11550 9982 11634 9983
rect 11326 9921 11354 9926
rect 11438 9954 11466 9959
rect 11438 9907 11466 9926
rect 11494 9618 11522 9623
rect 11494 9571 11522 9590
rect 11270 9561 11298 9567
rect 11270 9535 11271 9561
rect 11297 9535 11298 9561
rect 11270 9506 11298 9535
rect 11270 9473 11298 9478
rect 11438 9226 11466 9231
rect 11438 9179 11466 9198
rect 11270 9169 11298 9175
rect 11270 9143 11271 9169
rect 11297 9143 11298 9169
rect 11270 9114 11298 9143
rect 11550 9114 11578 9982
rect 11606 9977 11634 9982
rect 11662 11018 11690 11023
rect 11662 10793 11690 10990
rect 11662 10767 11663 10793
rect 11689 10767 11690 10793
rect 11662 10010 11690 10767
rect 11690 9982 11746 10010
rect 11662 9977 11690 9982
rect 11606 9898 11634 9903
rect 11606 9851 11634 9870
rect 11662 9842 11690 9847
rect 11662 9617 11690 9814
rect 11718 9786 11746 9982
rect 11718 9753 11746 9758
rect 11830 10009 11858 10015
rect 11830 9983 11831 10009
rect 11857 9983 11858 10009
rect 11830 9674 11858 9983
rect 11886 9842 11914 11551
rect 11886 9809 11914 9814
rect 11830 9641 11858 9646
rect 11942 9618 11970 11662
rect 12054 11689 12082 11886
rect 12054 11663 12055 11689
rect 12081 11663 12082 11689
rect 12054 11657 12082 11663
rect 11998 11634 12026 11639
rect 11998 11587 12026 11606
rect 12166 11633 12194 12335
rect 13006 12082 13034 12390
rect 13062 12362 13090 13119
rect 14630 13146 14658 13151
rect 13398 13090 13426 13095
rect 14182 13090 14210 13095
rect 13398 13089 13482 13090
rect 13398 13063 13399 13089
rect 13425 13063 13482 13089
rect 13398 13062 13482 13063
rect 13398 13057 13426 13062
rect 13454 12753 13482 13062
rect 13454 12727 13455 12753
rect 13481 12727 13482 12753
rect 13454 12721 13482 12727
rect 13622 12782 14042 12810
rect 13622 12753 13650 12782
rect 13622 12727 13623 12753
rect 13649 12727 13650 12753
rect 13622 12721 13650 12727
rect 14014 12754 14042 12782
rect 14070 12754 14098 12759
rect 14014 12753 14098 12754
rect 14014 12727 14071 12753
rect 14097 12727 14098 12753
rect 14014 12726 14098 12727
rect 14070 12721 14098 12726
rect 13958 12698 13986 12703
rect 13958 12651 13986 12670
rect 14182 12697 14210 13062
rect 14462 13090 14490 13095
rect 14462 13043 14490 13062
rect 14238 12754 14266 12759
rect 14238 12707 14266 12726
rect 14574 12754 14602 12759
rect 14574 12707 14602 12726
rect 14182 12671 14183 12697
rect 14209 12671 14210 12697
rect 14182 12665 14210 12671
rect 14630 12697 14658 13118
rect 18830 13146 18858 13151
rect 18830 13099 18858 13118
rect 14630 12671 14631 12697
rect 14657 12671 14658 12697
rect 13566 12641 13594 12647
rect 13566 12615 13567 12641
rect 13593 12615 13594 12641
rect 13062 12329 13090 12334
rect 13342 12362 13370 12367
rect 13006 12025 13034 12054
rect 13006 11999 13007 12025
rect 13033 11999 13034 12025
rect 13006 11993 13034 11999
rect 13230 11970 13258 11975
rect 13342 11970 13370 12334
rect 13258 11942 13370 11970
rect 13230 11923 13258 11942
rect 12166 11607 12167 11633
rect 12193 11607 12194 11633
rect 12166 11601 12194 11607
rect 12222 11354 12250 11359
rect 12222 11242 12250 11326
rect 12950 11298 12978 11303
rect 12222 11195 12250 11214
rect 12502 11241 12530 11247
rect 12502 11215 12503 11241
rect 12529 11215 12530 11241
rect 12278 11186 12306 11191
rect 12278 11139 12306 11158
rect 12502 11186 12530 11215
rect 12502 11153 12530 11158
rect 12894 11242 12922 11247
rect 12894 11129 12922 11214
rect 12894 11103 12895 11129
rect 12921 11103 12922 11129
rect 12726 11074 12754 11079
rect 12726 11073 12866 11074
rect 12726 11047 12727 11073
rect 12753 11047 12866 11073
rect 12726 11046 12866 11047
rect 12726 11041 12754 11046
rect 12726 10738 12754 10743
rect 12502 10402 12530 10407
rect 12278 10066 12306 10071
rect 12054 9618 12082 9623
rect 11662 9591 11663 9617
rect 11689 9591 11690 9617
rect 11662 9585 11690 9591
rect 11886 9590 11970 9618
rect 11998 9590 12054 9618
rect 11774 9562 11802 9567
rect 11886 9562 11914 9590
rect 11774 9561 11914 9562
rect 11774 9535 11775 9561
rect 11801 9535 11914 9561
rect 11774 9534 11914 9535
rect 11662 9505 11690 9511
rect 11662 9479 11663 9505
rect 11689 9479 11690 9505
rect 11270 9086 11578 9114
rect 10878 8913 10906 8918
rect 10934 9030 11242 9058
rect 10934 8833 10962 9030
rect 10934 8807 10935 8833
rect 10961 8807 10962 8833
rect 10934 8801 10962 8807
rect 11046 8553 11074 9030
rect 11046 8527 11047 8553
rect 11073 8527 11074 8553
rect 11046 8498 11074 8527
rect 11046 8465 11074 8470
rect 11326 8890 11354 8895
rect 11326 8554 11354 8862
rect 10878 8441 10906 8447
rect 10878 8415 10879 8441
rect 10905 8415 10906 8441
rect 10878 8386 10906 8415
rect 11214 8442 11242 8447
rect 11214 8395 11242 8414
rect 10878 8353 10906 8358
rect 11326 8105 11354 8526
rect 11326 8079 11327 8105
rect 11353 8079 11354 8105
rect 11326 8073 11354 8079
rect 11382 8497 11410 8503
rect 11382 8471 11383 8497
rect 11409 8471 11410 8497
rect 10654 7713 10850 7714
rect 10654 7687 10655 7713
rect 10681 7687 10850 7713
rect 10654 7686 10850 7687
rect 10654 7681 10682 7686
rect 9422 7658 9450 7663
rect 9422 7611 9450 7630
rect 10150 7658 10178 7663
rect 10374 7658 10402 7663
rect 10150 7657 10402 7658
rect 10150 7631 10151 7657
rect 10177 7631 10375 7657
rect 10401 7631 10402 7657
rect 10150 7630 10402 7631
rect 10150 7625 10178 7630
rect 9310 7569 9338 7574
rect 9254 7322 9282 7327
rect 9198 7321 9282 7322
rect 9198 7295 9255 7321
rect 9281 7295 9282 7321
rect 9198 7294 9282 7295
rect 9254 7289 9282 7294
rect 10318 7321 10346 7630
rect 10374 7625 10402 7630
rect 11382 7658 11410 8471
rect 11494 7770 11522 7775
rect 11382 7625 11410 7630
rect 11438 7769 11522 7770
rect 11438 7743 11495 7769
rect 11521 7743 11522 7769
rect 11438 7742 11522 7743
rect 10318 7295 10319 7321
rect 10345 7295 10346 7321
rect 10318 7289 10346 7295
rect 11438 7322 11466 7742
rect 11494 7737 11522 7742
rect 11550 7546 11578 9086
rect 11606 9169 11634 9175
rect 11606 9143 11607 9169
rect 11633 9143 11634 9169
rect 11606 9114 11634 9143
rect 11606 9081 11634 9086
rect 11662 8385 11690 9479
rect 11774 9450 11802 9534
rect 11998 9506 12026 9590
rect 12054 9571 12082 9590
rect 12278 9617 12306 10038
rect 12278 9591 12279 9617
rect 12305 9591 12306 9617
rect 11774 9417 11802 9422
rect 11830 9478 12026 9506
rect 12222 9562 12250 9567
rect 11830 9337 11858 9478
rect 11830 9311 11831 9337
rect 11857 9311 11858 9337
rect 11830 9305 11858 9311
rect 12222 9281 12250 9534
rect 12278 9337 12306 9591
rect 12390 9730 12418 9735
rect 12390 9617 12418 9702
rect 12502 9673 12530 10374
rect 12558 10346 12586 10351
rect 12586 10318 12642 10346
rect 12558 10299 12586 10318
rect 12502 9647 12503 9673
rect 12529 9647 12530 9673
rect 12502 9641 12530 9647
rect 12558 10010 12586 10015
rect 12390 9591 12391 9617
rect 12417 9591 12418 9617
rect 12390 9585 12418 9591
rect 12558 9617 12586 9982
rect 12614 10009 12642 10318
rect 12614 9983 12615 10009
rect 12641 9983 12642 10009
rect 12614 9977 12642 9983
rect 12558 9591 12559 9617
rect 12585 9591 12586 9617
rect 12558 9585 12586 9591
rect 12726 9617 12754 10710
rect 12726 9591 12727 9617
rect 12753 9591 12754 9617
rect 12726 9585 12754 9591
rect 12838 9618 12866 11046
rect 12894 10738 12922 11103
rect 12950 11130 12978 11270
rect 12950 11083 12978 11102
rect 13566 11130 13594 12615
rect 13790 12641 13818 12647
rect 13790 12615 13791 12641
rect 13817 12615 13818 12641
rect 13734 12418 13762 12423
rect 13790 12418 13818 12615
rect 13734 12417 13818 12418
rect 13734 12391 13735 12417
rect 13761 12391 13818 12417
rect 13734 12390 13818 12391
rect 13902 12641 13930 12647
rect 13902 12615 13903 12641
rect 13929 12615 13930 12641
rect 13734 12385 13762 12390
rect 13566 11097 13594 11102
rect 13062 11073 13090 11079
rect 13062 11047 13063 11073
rect 13089 11047 13090 11073
rect 12894 10710 13034 10738
rect 12894 9618 12922 9623
rect 12866 9617 12922 9618
rect 12866 9591 12895 9617
rect 12921 9591 12922 9617
rect 12866 9590 12922 9591
rect 12838 9571 12866 9590
rect 12894 9585 12922 9590
rect 12278 9311 12279 9337
rect 12305 9311 12306 9337
rect 12278 9305 12306 9311
rect 12222 9255 12223 9281
rect 12249 9255 12250 9281
rect 12222 9249 12250 9255
rect 11774 9225 11802 9231
rect 11774 9199 11775 9225
rect 11801 9199 11802 9225
rect 11774 8890 11802 9199
rect 12390 9226 12418 9231
rect 12390 9179 12418 9198
rect 12950 9226 12978 9231
rect 12950 9179 12978 9198
rect 12838 9170 12866 9175
rect 11774 8857 11802 8862
rect 12782 9169 12866 9170
rect 12782 9143 12839 9169
rect 12865 9143 12866 9169
rect 12782 9142 12866 9143
rect 12782 9114 12810 9142
rect 12838 9137 12866 9142
rect 12670 8834 12698 8839
rect 12782 8834 12810 9086
rect 12698 8806 12810 8834
rect 12838 8833 12866 8839
rect 12838 8807 12839 8833
rect 12865 8807 12866 8833
rect 12670 8787 12698 8806
rect 11774 8722 11802 8727
rect 11774 8554 11802 8694
rect 11662 8359 11663 8385
rect 11689 8359 11690 8385
rect 11662 8353 11690 8359
rect 11718 8553 11802 8554
rect 11718 8527 11775 8553
rect 11801 8527 11802 8553
rect 11718 8526 11802 8527
rect 11606 7658 11634 7663
rect 11718 7658 11746 8526
rect 11774 8521 11802 8526
rect 12838 8553 12866 8807
rect 13006 8833 13034 10710
rect 13062 10514 13090 11047
rect 13790 10738 13818 10743
rect 13790 10737 13874 10738
rect 13790 10711 13791 10737
rect 13817 10711 13874 10737
rect 13790 10710 13874 10711
rect 13790 10705 13818 10710
rect 13062 10481 13090 10486
rect 13566 10514 13594 10519
rect 13790 10514 13818 10519
rect 13566 10467 13594 10486
rect 13622 10513 13818 10514
rect 13622 10487 13791 10513
rect 13817 10487 13818 10513
rect 13622 10486 13818 10487
rect 13846 10514 13874 10710
rect 13902 10682 13930 12615
rect 14350 12362 14378 12367
rect 14182 11634 14210 11639
rect 14182 11587 14210 11606
rect 14070 11578 14098 11583
rect 14070 11531 14098 11550
rect 14350 11578 14378 12334
rect 14630 12250 14658 12671
rect 14686 13089 14714 13095
rect 14686 13063 14687 13089
rect 14713 13063 14714 13089
rect 14686 12362 14714 13063
rect 18942 13090 18970 13511
rect 20006 13146 20034 13567
rect 20006 13113 20034 13118
rect 18942 13057 18970 13062
rect 20006 13033 20034 13039
rect 20006 13007 20007 13033
rect 20033 13007 20034 13033
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 20006 12810 20034 13007
rect 20006 12777 20034 12782
rect 14742 12698 14770 12703
rect 14742 12651 14770 12670
rect 14686 12329 14714 12334
rect 15022 12362 15050 12367
rect 15022 12315 15050 12334
rect 14798 12305 14826 12311
rect 14798 12279 14799 12305
rect 14825 12279 14826 12305
rect 14798 12250 14826 12279
rect 14630 12222 14826 12250
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 18830 11970 18858 11975
rect 18830 11923 18858 11942
rect 20006 11802 20034 11999
rect 20006 11769 20034 11774
rect 14742 11634 14770 11639
rect 14742 11587 14770 11606
rect 14966 11578 14994 11583
rect 14350 11577 14434 11578
rect 14350 11551 14351 11577
rect 14377 11551 14434 11577
rect 14350 11550 14434 11551
rect 14350 11545 14378 11550
rect 14406 11522 14434 11550
rect 14014 11242 14042 11247
rect 14014 11195 14042 11214
rect 14126 11186 14154 11191
rect 14126 11139 14154 11158
rect 14294 11074 14322 11079
rect 14294 11027 14322 11046
rect 14406 10906 14434 11494
rect 14966 11297 14994 11550
rect 18830 11578 18858 11583
rect 18830 11531 18858 11550
rect 14966 11271 14967 11297
rect 14993 11271 14994 11297
rect 14966 11265 14994 11271
rect 15806 11521 15834 11527
rect 15806 11495 15807 11521
rect 15833 11495 15834 11521
rect 15806 11466 15834 11495
rect 16030 11522 16058 11527
rect 16030 11475 16058 11494
rect 15806 11242 15834 11438
rect 20006 11466 20034 11471
rect 20006 11419 20034 11438
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 14182 10905 14434 10906
rect 14182 10879 14407 10905
rect 14433 10879 14434 10905
rect 14182 10878 14434 10879
rect 14182 10793 14210 10878
rect 14182 10767 14183 10793
rect 14209 10767 14210 10793
rect 14182 10761 14210 10767
rect 13902 10654 14210 10682
rect 13846 10486 13986 10514
rect 13454 10402 13482 10407
rect 13454 10355 13482 10374
rect 13622 10094 13650 10486
rect 13790 10481 13818 10486
rect 13398 10066 13426 10071
rect 13062 9842 13090 9847
rect 13062 9561 13090 9814
rect 13398 9842 13426 10038
rect 13398 9673 13426 9814
rect 13398 9647 13399 9673
rect 13425 9647 13426 9673
rect 13398 9641 13426 9647
rect 13454 10066 13650 10094
rect 13678 10401 13706 10407
rect 13678 10375 13679 10401
rect 13705 10375 13706 10401
rect 13678 10094 13706 10375
rect 13846 10345 13874 10351
rect 13846 10319 13847 10345
rect 13873 10319 13874 10345
rect 13846 10178 13874 10319
rect 13958 10290 13986 10486
rect 14126 10402 14154 10407
rect 14070 10401 14154 10402
rect 14070 10375 14127 10401
rect 14153 10375 14154 10401
rect 14070 10374 14154 10375
rect 14014 10290 14042 10295
rect 13958 10289 14042 10290
rect 13958 10263 14015 10289
rect 14041 10263 14042 10289
rect 13958 10262 14042 10263
rect 14014 10257 14042 10262
rect 14070 10178 14098 10374
rect 14126 10369 14154 10374
rect 14182 10402 14210 10654
rect 13846 10150 14098 10178
rect 14182 10094 14210 10374
rect 13678 10066 14098 10094
rect 13062 9535 13063 9561
rect 13089 9535 13090 9561
rect 13062 9529 13090 9535
rect 13398 9281 13426 9287
rect 13398 9255 13399 9281
rect 13425 9255 13426 9281
rect 13118 9170 13146 9175
rect 13118 9123 13146 9142
rect 13006 8807 13007 8833
rect 13033 8807 13034 8833
rect 13006 8801 13034 8807
rect 13286 9113 13314 9119
rect 13286 9087 13287 9113
rect 13313 9087 13314 9113
rect 12894 8721 12922 8727
rect 12894 8695 12895 8721
rect 12921 8695 12922 8721
rect 12894 8610 12922 8695
rect 12894 8582 13146 8610
rect 12838 8527 12839 8553
rect 12865 8527 12866 8553
rect 12838 8521 12866 8527
rect 12950 8498 12978 8503
rect 12950 8451 12978 8470
rect 12894 8442 12922 8447
rect 12894 8386 12922 8414
rect 13006 8441 13034 8447
rect 13006 8415 13007 8441
rect 13033 8415 13034 8441
rect 13006 8386 13034 8415
rect 12894 8358 13034 8386
rect 13062 8442 13090 8447
rect 11830 8330 11858 8335
rect 11830 8329 12418 8330
rect 11830 8303 11831 8329
rect 11857 8303 12418 8329
rect 11830 8302 12418 8303
rect 11830 8297 11858 8302
rect 12390 8105 12418 8302
rect 13006 8106 13034 8111
rect 13062 8106 13090 8414
rect 12390 8079 12391 8105
rect 12417 8079 12418 8105
rect 12390 8073 12418 8079
rect 12782 8105 13090 8106
rect 12782 8079 13007 8105
rect 13033 8079 13090 8105
rect 12782 8078 13090 8079
rect 12782 8050 12810 8078
rect 13006 8073 13034 8078
rect 12670 8049 12810 8050
rect 12670 8023 12783 8049
rect 12809 8023 12810 8049
rect 12670 8022 12810 8023
rect 12110 7770 12138 7775
rect 11774 7769 12138 7770
rect 11774 7743 12111 7769
rect 12137 7743 12138 7769
rect 11774 7742 12138 7743
rect 11774 7713 11802 7742
rect 12110 7737 12138 7742
rect 11774 7687 11775 7713
rect 11801 7687 11802 7713
rect 11774 7681 11802 7687
rect 11606 7657 11746 7658
rect 11606 7631 11607 7657
rect 11633 7631 11746 7657
rect 11606 7630 11746 7631
rect 11886 7658 11914 7663
rect 11606 7625 11634 7630
rect 11886 7611 11914 7630
rect 12670 7657 12698 8022
rect 12782 8017 12810 8022
rect 13118 7994 13146 8582
rect 13286 8274 13314 9087
rect 13398 8554 13426 9255
rect 13454 9169 13482 10066
rect 13510 9954 13538 9959
rect 13510 9729 13538 9926
rect 13510 9703 13511 9729
rect 13537 9703 13538 9729
rect 13510 9697 13538 9703
rect 13678 9618 13706 9623
rect 13790 9618 13818 9623
rect 13678 9617 13818 9618
rect 13678 9591 13679 9617
rect 13705 9591 13791 9617
rect 13817 9591 13818 9617
rect 13678 9590 13818 9591
rect 13678 9585 13706 9590
rect 13790 9585 13818 9590
rect 14070 9617 14098 10066
rect 14070 9591 14071 9617
rect 14097 9591 14098 9617
rect 13958 9561 13986 9567
rect 13958 9535 13959 9561
rect 13985 9535 13986 9561
rect 13958 9506 13986 9535
rect 13958 9473 13986 9478
rect 13790 9338 13818 9343
rect 13678 9281 13706 9287
rect 13678 9255 13679 9281
rect 13705 9255 13706 9281
rect 13622 9226 13650 9231
rect 13622 9179 13650 9198
rect 13454 9143 13455 9169
rect 13481 9143 13482 9169
rect 13454 9137 13482 9143
rect 13678 9114 13706 9255
rect 13790 9225 13818 9310
rect 13790 9199 13791 9225
rect 13817 9199 13818 9225
rect 13790 9193 13818 9199
rect 14014 9338 14042 9343
rect 13678 9081 13706 9086
rect 13398 8521 13426 8526
rect 13958 8778 13986 8783
rect 13958 8498 13986 8750
rect 13846 8442 13874 8447
rect 13846 8395 13874 8414
rect 13286 8241 13314 8246
rect 13006 7966 13146 7994
rect 13006 7713 13034 7966
rect 13006 7687 13007 7713
rect 13033 7687 13034 7713
rect 13006 7681 13034 7687
rect 12670 7631 12671 7657
rect 12697 7631 12698 7657
rect 12166 7601 12194 7607
rect 12166 7575 12167 7601
rect 12193 7575 12194 7601
rect 11606 7546 11634 7551
rect 11550 7545 11634 7546
rect 11550 7519 11607 7545
rect 11633 7519 11634 7545
rect 11550 7518 11634 7519
rect 11606 7513 11634 7518
rect 11494 7322 11522 7327
rect 11438 7321 11522 7322
rect 11438 7295 11495 7321
rect 11521 7295 11522 7321
rect 11438 7294 11522 7295
rect 12166 7322 12194 7575
rect 12558 7322 12586 7327
rect 12166 7321 12586 7322
rect 12166 7295 12559 7321
rect 12585 7295 12586 7321
rect 12166 7294 12586 7295
rect 11494 7289 11522 7294
rect 8918 7266 8946 7271
rect 8078 7233 8106 7238
rect 8862 7238 8918 7266
rect 7630 7126 7882 7154
rect 8862 6985 8890 7238
rect 8918 7219 8946 7238
rect 10710 7266 10738 7271
rect 10710 7219 10738 7238
rect 11158 7266 11186 7271
rect 11158 7219 11186 7238
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 8862 6959 8863 6985
rect 8889 6959 8890 6985
rect 8862 6953 8890 6959
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 12558 4214 12586 7294
rect 12670 7266 12698 7631
rect 13958 7602 13986 8470
rect 14014 8050 14042 9310
rect 14070 9170 14098 9591
rect 14126 10066 14210 10094
rect 14126 9506 14154 10066
rect 14406 9954 14434 10878
rect 14518 11214 14714 11242
rect 14518 10457 14546 11214
rect 14686 11185 14714 11214
rect 15806 11209 15834 11214
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 14686 11159 14687 11185
rect 14713 11159 14714 11185
rect 14686 11153 14714 11159
rect 18830 11185 18858 11191
rect 18830 11159 18831 11185
rect 18857 11159 18858 11185
rect 14518 10431 14519 10457
rect 14545 10431 14546 10457
rect 14518 10425 14546 10431
rect 14630 11129 14658 11135
rect 14630 11103 14631 11129
rect 14657 11103 14658 11129
rect 14574 10345 14602 10351
rect 14574 10319 14575 10345
rect 14601 10319 14602 10345
rect 14574 10066 14602 10319
rect 14574 10033 14602 10038
rect 14574 9954 14602 9959
rect 14406 9953 14602 9954
rect 14406 9927 14575 9953
rect 14601 9927 14602 9953
rect 14406 9926 14602 9927
rect 14294 9898 14322 9903
rect 14126 9473 14154 9478
rect 14182 9617 14210 9623
rect 14182 9591 14183 9617
rect 14209 9591 14210 9617
rect 14070 8834 14098 9142
rect 14070 8801 14098 8806
rect 14126 9226 14154 9231
rect 14126 8722 14154 9198
rect 14182 8834 14210 9591
rect 14294 9617 14322 9870
rect 14294 9591 14295 9617
rect 14321 9591 14322 9617
rect 14294 9585 14322 9591
rect 14574 9617 14602 9926
rect 14574 9591 14575 9617
rect 14601 9591 14602 9617
rect 14350 9562 14378 9567
rect 14350 9505 14378 9534
rect 14350 9479 14351 9505
rect 14377 9479 14378 9505
rect 14350 9473 14378 9479
rect 14574 9226 14602 9591
rect 14630 9338 14658 11103
rect 14742 11129 14770 11135
rect 14742 11103 14743 11129
rect 14769 11103 14770 11129
rect 14742 11074 14770 11103
rect 14742 11041 14770 11046
rect 14798 11130 14826 11135
rect 14798 10401 14826 11102
rect 18830 10738 18858 11159
rect 20006 10794 20034 11215
rect 20006 10761 20034 10766
rect 18830 10705 18858 10710
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 20006 10457 20034 10463
rect 20006 10431 20007 10457
rect 20033 10431 20034 10457
rect 14798 10375 14799 10401
rect 14825 10375 14826 10401
rect 14798 10369 14826 10375
rect 14854 10402 14882 10407
rect 14854 10355 14882 10374
rect 18830 10401 18858 10407
rect 18830 10375 18831 10401
rect 18857 10375 18858 10401
rect 14630 9305 14658 9310
rect 14686 10289 14714 10295
rect 14686 10263 14687 10289
rect 14713 10263 14714 10289
rect 14686 9954 14714 10263
rect 14574 9193 14602 9198
rect 14462 9170 14490 9175
rect 14462 9169 14546 9170
rect 14462 9143 14463 9169
rect 14489 9143 14546 9169
rect 14462 9142 14546 9143
rect 14462 9137 14490 9142
rect 14182 8806 14378 8834
rect 14294 8722 14322 8727
rect 14126 8721 14322 8722
rect 14126 8695 14295 8721
rect 14321 8695 14322 8721
rect 14126 8694 14322 8695
rect 14294 8442 14322 8694
rect 14350 8554 14378 8806
rect 14518 8722 14546 9142
rect 14574 8834 14602 8839
rect 14574 8787 14602 8806
rect 14686 8833 14714 9926
rect 15470 9953 15498 9959
rect 15470 9927 15471 9953
rect 15497 9927 15498 9953
rect 15414 9898 15442 9903
rect 15414 9851 15442 9870
rect 15470 9674 15498 9927
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 15470 9641 15498 9646
rect 16030 9674 16058 9679
rect 16030 9627 16058 9646
rect 18830 9674 18858 10375
rect 20006 10122 20034 10431
rect 20006 10089 20034 10094
rect 18830 9641 18858 9646
rect 14966 9562 14994 9567
rect 14966 9515 14994 9534
rect 18942 9225 18970 9231
rect 18942 9199 18943 9225
rect 18969 9199 18970 9225
rect 15526 9169 15554 9175
rect 15526 9143 15527 9169
rect 15553 9143 15554 9169
rect 15078 8945 15106 8951
rect 15078 8919 15079 8945
rect 15105 8919 15106 8945
rect 15078 8890 15106 8919
rect 14966 8862 15106 8890
rect 14686 8807 14687 8833
rect 14713 8807 14714 8833
rect 14686 8801 14714 8807
rect 14910 8834 14938 8839
rect 14966 8834 14994 8862
rect 14910 8833 14994 8834
rect 14910 8807 14911 8833
rect 14937 8807 14994 8833
rect 14910 8806 14994 8807
rect 14910 8801 14938 8806
rect 15022 8777 15050 8783
rect 15022 8751 15023 8777
rect 15049 8751 15050 8777
rect 14742 8722 14770 8727
rect 14518 8721 14770 8722
rect 14518 8695 14743 8721
rect 14769 8695 14770 8721
rect 14518 8694 14770 8695
rect 14742 8689 14770 8694
rect 14350 8521 14378 8526
rect 14686 8554 14714 8559
rect 14238 8385 14266 8391
rect 14238 8359 14239 8385
rect 14265 8359 14266 8385
rect 14182 8162 14210 8167
rect 14238 8162 14266 8359
rect 14182 8161 14266 8162
rect 14182 8135 14183 8161
rect 14209 8135 14266 8161
rect 14182 8134 14266 8135
rect 14182 8129 14210 8134
rect 14014 8022 14210 8050
rect 14182 7993 14210 8022
rect 14182 7967 14183 7993
rect 14209 7967 14210 7993
rect 14182 7961 14210 7967
rect 14238 7994 14266 7999
rect 14238 7947 14266 7966
rect 14294 7769 14322 8414
rect 14630 8050 14658 8055
rect 14518 7994 14546 7999
rect 14518 7947 14546 7966
rect 14630 7993 14658 8022
rect 14630 7967 14631 7993
rect 14657 7967 14658 7993
rect 14630 7961 14658 7967
rect 14686 7993 14714 8526
rect 15022 8554 15050 8751
rect 15078 8721 15106 8727
rect 15078 8695 15079 8721
rect 15105 8695 15106 8721
rect 15078 8666 15106 8695
rect 15078 8633 15106 8638
rect 15526 8666 15554 9143
rect 15526 8633 15554 8638
rect 15750 9169 15778 9175
rect 15750 9143 15751 9169
rect 15777 9143 15778 9169
rect 15022 8521 15050 8526
rect 15526 8442 15554 8447
rect 15750 8442 15778 9143
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 18942 8666 18970 9199
rect 20006 9114 20034 9119
rect 20006 9067 20034 9086
rect 18942 8633 18970 8638
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 15554 8414 15778 8442
rect 18830 8441 18858 8447
rect 18830 8415 18831 8441
rect 18857 8415 18858 8441
rect 15526 8395 15554 8414
rect 15022 8386 15050 8391
rect 15022 8050 15050 8358
rect 15302 8386 15330 8391
rect 15302 8339 15330 8358
rect 18830 8386 18858 8415
rect 20006 8442 20034 8863
rect 20006 8409 20034 8414
rect 18830 8353 18858 8358
rect 19950 8385 19978 8391
rect 19950 8359 19951 8385
rect 19977 8359 19978 8385
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 19950 8106 19978 8359
rect 19950 8073 19978 8078
rect 20006 8105 20034 8111
rect 20006 8079 20007 8105
rect 20033 8079 20034 8105
rect 15022 8003 15050 8022
rect 18830 8050 18858 8055
rect 18830 8003 18858 8022
rect 14686 7967 14687 7993
rect 14713 7967 14714 7993
rect 14294 7743 14295 7769
rect 14321 7743 14322 7769
rect 14294 7737 14322 7743
rect 14686 7658 14714 7967
rect 15134 7938 15162 7943
rect 15134 7891 15162 7910
rect 20006 7770 20034 8079
rect 20006 7737 20034 7742
rect 14686 7625 14714 7630
rect 14070 7602 14098 7607
rect 13958 7601 14098 7602
rect 13958 7575 14071 7601
rect 14097 7575 14098 7601
rect 13958 7574 14098 7575
rect 14070 7569 14098 7574
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 12670 7233 12698 7238
rect 12838 7266 12866 7271
rect 12838 7219 12866 7238
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 12278 4186 12586 4214
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 12110 1834 12138 1839
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 12110 400 12138 1806
rect 12278 1777 12306 4186
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1745 12306 1751
rect 12096 0 12152 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 8974 19025 9002 19026
rect 8974 18999 8975 19025
rect 8975 18999 9001 19025
rect 9001 18999 9002 19025
rect 8974 18998 9002 18999
rect 9310 18998 9338 19026
rect 8078 18326 8106 18354
rect 8694 18353 8722 18354
rect 8694 18327 8695 18353
rect 8695 18327 8721 18353
rect 8721 18327 8722 18353
rect 8694 18326 8722 18327
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 11438 19110 11466 19138
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 9758 18718 9786 18746
rect 10374 18745 10402 18746
rect 10374 18719 10375 18745
rect 10375 18719 10401 18745
rect 10401 18719 10402 18745
rect 10374 18718 10402 18719
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 2086 13454 2114 13482
rect 966 12782 994 12810
rect 966 11774 994 11802
rect 966 11465 994 11466
rect 966 11439 967 11465
rect 967 11439 993 11465
rect 993 11439 994 11465
rect 966 11438 994 11439
rect 966 10766 994 10794
rect 2142 13145 2170 13146
rect 2142 13119 2143 13145
rect 2143 13119 2169 13145
rect 2169 13119 2170 13145
rect 2142 13118 2170 13119
rect 6062 13118 6090 13146
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 6062 12670 6090 12698
rect 6454 12278 6482 12306
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 2142 11969 2170 11970
rect 2142 11943 2143 11969
rect 2143 11943 2169 11969
rect 2169 11943 2170 11969
rect 2142 11942 2170 11943
rect 7182 13089 7210 13090
rect 7182 13063 7183 13089
rect 7183 13063 7209 13089
rect 7209 13063 7210 13089
rect 7182 13062 7210 13063
rect 7910 12782 7938 12810
rect 7966 13062 7994 13090
rect 7350 12753 7378 12754
rect 7350 12727 7351 12753
rect 7351 12727 7377 12753
rect 7377 12727 7378 12753
rect 7350 12726 7378 12727
rect 7574 12753 7602 12754
rect 7574 12727 7575 12753
rect 7575 12727 7601 12753
rect 7601 12727 7602 12753
rect 7574 12726 7602 12727
rect 7238 12697 7266 12698
rect 7238 12671 7239 12697
rect 7239 12671 7265 12697
rect 7265 12671 7266 12697
rect 7238 12670 7266 12671
rect 7182 12614 7210 12642
rect 7462 12558 7490 12586
rect 6846 12278 6874 12306
rect 7070 12278 7098 12306
rect 7518 12278 7546 12306
rect 7742 12305 7770 12306
rect 7742 12279 7743 12305
rect 7743 12279 7769 12305
rect 7769 12279 7770 12305
rect 7742 12278 7770 12279
rect 4998 11886 5026 11914
rect 6790 11913 6818 11914
rect 6790 11887 6791 11913
rect 6791 11887 6817 11913
rect 6817 11887 6818 11913
rect 6790 11886 6818 11887
rect 7070 11886 7098 11914
rect 2142 11494 2170 11522
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 6398 11270 6426 11298
rect 6398 10878 6426 10906
rect 6846 11521 6874 11522
rect 6846 11495 6847 11521
rect 6847 11495 6873 11521
rect 6873 11495 6874 11521
rect 6846 11494 6874 11495
rect 2142 10710 2170 10738
rect 4942 10766 4970 10794
rect 6566 10793 6594 10794
rect 6566 10767 6567 10793
rect 6567 10767 6593 10793
rect 6593 10767 6594 10793
rect 6566 10766 6594 10767
rect 5838 10710 5866 10738
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 2086 10486 2114 10514
rect 6790 10793 6818 10794
rect 6790 10767 6791 10793
rect 6791 10767 6817 10793
rect 6817 10767 6818 10793
rect 6790 10766 6818 10767
rect 6734 10737 6762 10738
rect 6734 10711 6735 10737
rect 6735 10711 6761 10737
rect 6761 10711 6762 10737
rect 6734 10710 6762 10711
rect 6902 10822 6930 10850
rect 966 10094 994 10122
rect 966 9897 994 9898
rect 966 9871 967 9897
rect 967 9871 993 9897
rect 993 9871 994 9897
rect 966 9870 994 9871
rect 6174 10065 6202 10066
rect 6174 10039 6175 10065
rect 6175 10039 6201 10065
rect 6201 10039 6202 10065
rect 6174 10038 6202 10039
rect 6846 10038 6874 10066
rect 2142 10009 2170 10010
rect 2142 9983 2143 10009
rect 2143 9983 2169 10009
rect 2169 9983 2170 10009
rect 2142 9982 2170 9983
rect 5726 9953 5754 9954
rect 5726 9927 5727 9953
rect 5727 9927 5753 9953
rect 5753 9927 5754 9953
rect 5726 9926 5754 9927
rect 2086 9870 2114 9898
rect 4830 9870 4858 9898
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 6286 9870 6314 9898
rect 6734 10009 6762 10010
rect 6734 9983 6735 10009
rect 6735 9983 6761 10009
rect 6761 9983 6762 10009
rect 6734 9982 6762 9983
rect 6678 9953 6706 9954
rect 6678 9927 6679 9953
rect 6679 9927 6705 9953
rect 6705 9927 6706 9953
rect 6678 9926 6706 9927
rect 6622 9870 6650 9898
rect 966 9422 994 9450
rect 5950 9478 5978 9506
rect 2142 9142 2170 9170
rect 4886 9169 4914 9170
rect 4886 9143 4887 9169
rect 4887 9143 4913 9169
rect 4913 9143 4914 9169
rect 4886 9142 4914 9143
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 2142 8833 2170 8834
rect 2142 8807 2143 8833
rect 2143 8807 2169 8833
rect 2169 8807 2170 8833
rect 2142 8806 2170 8807
rect 5950 8806 5978 8834
rect 966 8414 994 8442
rect 2142 8441 2170 8442
rect 2142 8415 2143 8441
rect 2143 8415 2169 8441
rect 2169 8415 2170 8441
rect 2142 8414 2170 8415
rect 5894 8414 5922 8442
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 966 8078 994 8106
rect 7742 11830 7770 11858
rect 8246 12782 8274 12810
rect 7798 11382 7826 11410
rect 7854 12502 7882 12530
rect 8414 12334 8442 12362
rect 7126 10905 7154 10906
rect 7126 10879 7127 10905
rect 7127 10879 7153 10905
rect 7153 10879 7154 10905
rect 7126 10878 7154 10879
rect 7630 10878 7658 10906
rect 7574 10849 7602 10850
rect 7574 10823 7575 10849
rect 7575 10823 7601 10849
rect 7601 10823 7602 10849
rect 7574 10822 7602 10823
rect 7742 10905 7770 10906
rect 7742 10879 7743 10905
rect 7743 10879 7769 10905
rect 7769 10879 7770 10905
rect 7742 10878 7770 10879
rect 7014 9870 7042 9898
rect 7182 9982 7210 10010
rect 6902 9617 6930 9618
rect 6902 9591 6903 9617
rect 6903 9591 6929 9617
rect 6929 9591 6930 9617
rect 6902 9590 6930 9591
rect 6846 9534 6874 9562
rect 7070 9534 7098 9562
rect 6902 9505 6930 9506
rect 6902 9479 6903 9505
rect 6903 9479 6929 9505
rect 6929 9479 6930 9505
rect 6902 9478 6930 9479
rect 6510 9169 6538 9170
rect 6510 9143 6511 9169
rect 6511 9143 6537 9169
rect 6537 9143 6538 9169
rect 6510 9142 6538 9143
rect 6510 8414 6538 8442
rect 7182 9310 7210 9338
rect 7910 11382 7938 11410
rect 8022 11494 8050 11522
rect 7966 11046 7994 11074
rect 8806 11942 8834 11970
rect 8358 11830 8386 11858
rect 8246 11774 8274 11802
rect 8638 11774 8666 11802
rect 8414 11718 8442 11746
rect 8694 11633 8722 11634
rect 8694 11607 8695 11633
rect 8695 11607 8721 11633
rect 8721 11607 8722 11633
rect 8694 11606 8722 11607
rect 8694 11382 8722 11410
rect 8414 11297 8442 11298
rect 8414 11271 8415 11297
rect 8415 11271 8441 11297
rect 8441 11271 8442 11297
rect 8414 11270 8442 11271
rect 8470 11185 8498 11186
rect 8470 11159 8471 11185
rect 8471 11159 8497 11185
rect 8497 11159 8498 11185
rect 8470 11158 8498 11159
rect 8694 11158 8722 11186
rect 9086 13201 9114 13202
rect 9086 13175 9087 13201
rect 9087 13175 9113 13201
rect 9113 13175 9114 13201
rect 9086 13174 9114 13175
rect 11494 14041 11522 14042
rect 11494 14015 11495 14041
rect 11495 14015 11521 14041
rect 11521 14015 11522 14041
rect 11494 14014 11522 14015
rect 10486 13790 10514 13818
rect 9366 13118 9394 13146
rect 9310 12809 9338 12810
rect 9310 12783 9311 12809
rect 9311 12783 9337 12809
rect 9337 12783 9338 12809
rect 9310 12782 9338 12783
rect 9366 12726 9394 12754
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9478 12697 9506 12698
rect 9478 12671 9479 12697
rect 9479 12671 9505 12697
rect 9505 12671 9506 12697
rect 9478 12670 9506 12671
rect 10318 12726 10346 12754
rect 9814 12614 9842 12642
rect 9590 12390 9618 12418
rect 9198 11942 9226 11970
rect 8862 11718 8890 11746
rect 8750 11073 8778 11074
rect 8750 11047 8751 11073
rect 8751 11047 8777 11073
rect 8777 11047 8778 11073
rect 8750 11046 8778 11047
rect 8414 10822 8442 10850
rect 8414 10710 8442 10738
rect 7742 9590 7770 9618
rect 7966 9310 7994 9338
rect 6790 8414 6818 8442
rect 7014 8470 7042 8498
rect 5894 7966 5922 7994
rect 7406 8889 7434 8890
rect 7406 8863 7407 8889
rect 7407 8863 7433 8889
rect 7433 8863 7434 8889
rect 7406 8862 7434 8863
rect 7686 8889 7714 8890
rect 7686 8863 7687 8889
rect 7687 8863 7713 8889
rect 7713 8863 7714 8889
rect 7686 8862 7714 8863
rect 7238 8833 7266 8834
rect 7238 8807 7239 8833
rect 7239 8807 7265 8833
rect 7265 8807 7266 8833
rect 7238 8806 7266 8807
rect 7182 8358 7210 8386
rect 7294 8582 7322 8610
rect 7574 8497 7602 8498
rect 7574 8471 7575 8497
rect 7575 8471 7601 8497
rect 7601 8471 7602 8497
rect 7574 8470 7602 8471
rect 7406 8441 7434 8442
rect 7406 8415 7407 8441
rect 7407 8415 7433 8441
rect 7433 8415 7434 8441
rect 7406 8414 7434 8415
rect 7630 8385 7658 8386
rect 7630 8359 7631 8385
rect 7631 8359 7657 8385
rect 7657 8359 7658 8385
rect 7630 8358 7658 8359
rect 7630 7993 7658 7994
rect 7630 7967 7631 7993
rect 7631 7967 7657 7993
rect 7657 7967 7658 7993
rect 7630 7966 7658 7967
rect 8302 8833 8330 8834
rect 8302 8807 8303 8833
rect 8303 8807 8329 8833
rect 8329 8807 8330 8833
rect 8302 8806 8330 8807
rect 8190 8777 8218 8778
rect 8190 8751 8191 8777
rect 8191 8751 8217 8777
rect 8217 8751 8218 8777
rect 8190 8750 8218 8751
rect 8078 8526 8106 8554
rect 7910 7713 7938 7714
rect 7910 7687 7911 7713
rect 7911 7687 7937 7713
rect 7937 7687 7938 7713
rect 7910 7686 7938 7687
rect 8806 10737 8834 10738
rect 8806 10711 8807 10737
rect 8807 10711 8833 10737
rect 8833 10711 8834 10737
rect 8806 10710 8834 10711
rect 9086 11550 9114 11578
rect 9478 11494 9506 11522
rect 9198 11382 9226 11410
rect 9142 11158 9170 11186
rect 8918 10878 8946 10906
rect 8918 10486 8946 10514
rect 8974 10822 9002 10850
rect 9030 10542 9058 10570
rect 9030 10150 9058 10178
rect 8974 9646 9002 9674
rect 8750 9534 8778 9562
rect 8750 8862 8778 8890
rect 8862 8777 8890 8778
rect 8862 8751 8863 8777
rect 8863 8751 8889 8777
rect 8889 8751 8890 8777
rect 8862 8750 8890 8751
rect 9310 10542 9338 10570
rect 9142 9814 9170 9842
rect 9366 10150 9394 10178
rect 10262 12670 10290 12698
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9646 12361 9674 12362
rect 9646 12335 9647 12361
rect 9647 12335 9673 12361
rect 9673 12335 9674 12361
rect 9646 12334 9674 12335
rect 9646 11969 9674 11970
rect 9646 11943 9647 11969
rect 9647 11943 9673 11969
rect 9673 11943 9674 11969
rect 9646 11942 9674 11943
rect 9646 11465 9674 11466
rect 9646 11439 9647 11465
rect 9647 11439 9673 11465
rect 9673 11439 9674 11465
rect 9646 11438 9674 11439
rect 9254 10038 9282 10066
rect 9366 9758 9394 9786
rect 9254 9702 9282 9730
rect 9198 9590 9226 9618
rect 9310 9561 9338 9562
rect 9310 9535 9311 9561
rect 9311 9535 9337 9561
rect 9337 9535 9338 9561
rect 9310 9534 9338 9535
rect 9534 9926 9562 9954
rect 9366 9198 9394 9226
rect 9758 10766 9786 10794
rect 10878 13537 10906 13538
rect 10878 13511 10879 13537
rect 10879 13511 10905 13537
rect 10905 13511 10906 13537
rect 10878 13510 10906 13511
rect 11270 13734 11298 13762
rect 11494 13817 11522 13818
rect 11494 13791 11495 13817
rect 11495 13791 11521 13817
rect 11521 13791 11522 13817
rect 11494 13790 11522 13791
rect 11550 13734 11578 13762
rect 11774 13566 11802 13594
rect 10934 12670 10962 12698
rect 11830 12726 11858 12754
rect 11214 12641 11242 12642
rect 11214 12615 11215 12641
rect 11215 12615 11241 12641
rect 11241 12615 11242 12641
rect 11214 12614 11242 12615
rect 11270 12473 11298 12474
rect 11270 12447 11271 12473
rect 11271 12447 11297 12473
rect 11297 12447 11298 12473
rect 11270 12446 11298 12447
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 12110 18718 12138 18746
rect 13118 18745 13146 18746
rect 13118 18719 13119 18745
rect 13119 18719 13145 18745
rect 13145 18719 13146 18745
rect 13118 18718 13146 18719
rect 12278 14014 12306 14042
rect 12278 13593 12306 13594
rect 12278 13567 12279 13593
rect 12279 13567 12305 13593
rect 12305 13567 12306 13593
rect 12278 13566 12306 13567
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 12614 13566 12642 13594
rect 12502 13537 12530 13538
rect 12502 13511 12503 13537
rect 12503 13511 12529 13537
rect 12529 13511 12530 13537
rect 12502 13510 12530 13511
rect 13006 13510 13034 13538
rect 11886 12446 11914 12474
rect 12054 12417 12082 12418
rect 12054 12391 12055 12417
rect 12055 12391 12081 12417
rect 12081 12391 12082 12417
rect 12054 12390 12082 12391
rect 13006 12390 13034 12418
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 9814 11270 9842 11298
rect 9926 11606 9954 11634
rect 10038 11438 10066 11466
rect 10262 11774 10290 11802
rect 10206 11662 10234 11690
rect 10206 11382 10234 11410
rect 10654 11633 10682 11634
rect 10654 11607 10655 11633
rect 10655 11607 10681 11633
rect 10681 11607 10682 11633
rect 10654 11606 10682 11607
rect 10374 11326 10402 11354
rect 10430 11577 10458 11578
rect 10430 11551 10431 11577
rect 10431 11551 10457 11577
rect 10457 11551 10458 11577
rect 10430 11550 10458 11551
rect 10430 11158 10458 11186
rect 10542 11494 10570 11522
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 10094 10934 10122 10962
rect 10038 10513 10066 10514
rect 10038 10487 10039 10513
rect 10039 10487 10065 10513
rect 10065 10487 10066 10513
rect 10038 10486 10066 10487
rect 10542 10934 10570 10962
rect 10990 11606 11018 11634
rect 10654 10934 10682 10962
rect 10934 10934 10962 10962
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9758 9982 9786 10010
rect 9814 9926 9842 9954
rect 9702 9646 9730 9674
rect 9702 9310 9730 9338
rect 9814 9814 9842 9842
rect 9646 9198 9674 9226
rect 9366 8918 9394 8946
rect 9702 8945 9730 8946
rect 9702 8919 9703 8945
rect 9703 8919 9729 8945
rect 9729 8919 9730 8945
rect 9702 8918 9730 8919
rect 9030 8777 9058 8778
rect 9030 8751 9031 8777
rect 9031 8751 9057 8777
rect 9057 8751 9058 8777
rect 9030 8750 9058 8751
rect 8974 8721 9002 8722
rect 8974 8695 8975 8721
rect 8975 8695 9001 8721
rect 9001 8695 9002 8721
rect 8974 8694 9002 8695
rect 9254 8694 9282 8722
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 7350 7238 7378 7266
rect 7686 7238 7714 7266
rect 8694 7574 8722 7602
rect 9310 8497 9338 8498
rect 9310 8471 9311 8497
rect 9311 8471 9337 8497
rect 9337 8471 9338 8497
rect 9310 8470 9338 8471
rect 9646 8582 9674 8610
rect 9702 8553 9730 8554
rect 9702 8527 9703 8553
rect 9703 8527 9729 8553
rect 9729 8527 9730 8553
rect 9702 8526 9730 8527
rect 9422 8441 9450 8442
rect 9422 8415 9423 8441
rect 9423 8415 9449 8441
rect 9449 8415 9450 8441
rect 9422 8414 9450 8415
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9926 9310 9954 9338
rect 10038 9225 10066 9226
rect 10038 9199 10039 9225
rect 10039 9199 10065 9225
rect 10065 9199 10066 9225
rect 10038 9198 10066 9199
rect 9926 9142 9954 9170
rect 9870 8833 9898 8834
rect 9870 8807 9871 8833
rect 9871 8807 9897 8833
rect 9897 8807 9898 8833
rect 9870 8806 9898 8807
rect 10262 10038 10290 10066
rect 10094 9086 10122 9114
rect 10150 9982 10178 10010
rect 9814 8582 9842 8610
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 9870 8385 9898 8386
rect 9870 8359 9871 8385
rect 9871 8359 9897 8385
rect 9897 8359 9898 8385
rect 9870 8358 9898 8359
rect 10094 8358 10122 8386
rect 10318 9926 10346 9954
rect 10430 10374 10458 10402
rect 10654 10401 10682 10402
rect 10654 10375 10655 10401
rect 10655 10375 10681 10401
rect 10681 10375 10682 10401
rect 10654 10374 10682 10375
rect 10654 10009 10682 10010
rect 10654 9983 10655 10009
rect 10655 9983 10681 10009
rect 10681 9983 10682 10009
rect 10654 9982 10682 9983
rect 10598 9702 10626 9730
rect 10262 9422 10290 9450
rect 10430 9142 10458 9170
rect 11214 11774 11242 11802
rect 11046 10990 11074 11018
rect 11606 11969 11634 11970
rect 11606 11943 11607 11969
rect 11607 11943 11633 11969
rect 11633 11943 11634 11969
rect 11606 11942 11634 11943
rect 11774 11886 11802 11914
rect 11886 11662 11914 11690
rect 11550 11606 11578 11634
rect 11382 10934 11410 10962
rect 11326 10318 11354 10346
rect 10990 9814 11018 9842
rect 10766 9086 10794 9114
rect 10766 8862 10794 8890
rect 10654 8777 10682 8778
rect 10654 8751 10655 8777
rect 10655 8751 10681 8777
rect 10681 8751 10682 8777
rect 10654 8750 10682 8751
rect 10150 8694 10178 8722
rect 9534 8246 9562 8274
rect 9366 7993 9394 7994
rect 9366 7967 9367 7993
rect 9367 7967 9393 7993
rect 9393 7967 9394 7993
rect 9366 7966 9394 7967
rect 9534 7686 9562 7714
rect 10766 8721 10794 8722
rect 10766 8695 10767 8721
rect 10767 8695 10793 8721
rect 10793 8695 10794 8721
rect 10766 8694 10794 8695
rect 10430 8526 10458 8554
rect 10542 8358 10570 8386
rect 9870 8049 9898 8050
rect 9870 8023 9871 8049
rect 9871 8023 9897 8049
rect 9897 8023 9898 8049
rect 9870 8022 9898 8023
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 11102 9169 11130 9170
rect 11102 9143 11103 9169
rect 11103 9143 11129 9169
rect 11129 9143 11130 9169
rect 11102 9142 11130 9143
rect 11270 10065 11298 10066
rect 11270 10039 11271 10065
rect 11271 10039 11297 10065
rect 11297 10039 11298 10065
rect 11270 10038 11298 10039
rect 11326 9926 11354 9954
rect 11438 9953 11466 9954
rect 11438 9927 11439 9953
rect 11439 9927 11465 9953
rect 11465 9927 11466 9953
rect 11438 9926 11466 9927
rect 11494 9617 11522 9618
rect 11494 9591 11495 9617
rect 11495 9591 11521 9617
rect 11521 9591 11522 9617
rect 11494 9590 11522 9591
rect 11270 9478 11298 9506
rect 11438 9225 11466 9226
rect 11438 9199 11439 9225
rect 11439 9199 11465 9225
rect 11465 9199 11466 9225
rect 11438 9198 11466 9199
rect 11662 10990 11690 11018
rect 11662 9982 11690 10010
rect 11606 9897 11634 9898
rect 11606 9871 11607 9897
rect 11607 9871 11633 9897
rect 11633 9871 11634 9897
rect 11606 9870 11634 9871
rect 11662 9814 11690 9842
rect 11718 9758 11746 9786
rect 11886 9814 11914 9842
rect 11830 9646 11858 9674
rect 11998 11633 12026 11634
rect 11998 11607 11999 11633
rect 11999 11607 12025 11633
rect 12025 11607 12026 11633
rect 11998 11606 12026 11607
rect 14630 13118 14658 13146
rect 14182 13062 14210 13090
rect 13958 12697 13986 12698
rect 13958 12671 13959 12697
rect 13959 12671 13985 12697
rect 13985 12671 13986 12697
rect 13958 12670 13986 12671
rect 14462 13089 14490 13090
rect 14462 13063 14463 13089
rect 14463 13063 14489 13089
rect 14489 13063 14490 13089
rect 14462 13062 14490 13063
rect 14238 12753 14266 12754
rect 14238 12727 14239 12753
rect 14239 12727 14265 12753
rect 14265 12727 14266 12753
rect 14238 12726 14266 12727
rect 14574 12753 14602 12754
rect 14574 12727 14575 12753
rect 14575 12727 14601 12753
rect 14601 12727 14602 12753
rect 14574 12726 14602 12727
rect 18830 13145 18858 13146
rect 18830 13119 18831 13145
rect 18831 13119 18857 13145
rect 18857 13119 18858 13145
rect 18830 13118 18858 13119
rect 13062 12334 13090 12362
rect 13342 12361 13370 12362
rect 13342 12335 13343 12361
rect 13343 12335 13369 12361
rect 13369 12335 13370 12361
rect 13342 12334 13370 12335
rect 13006 12054 13034 12082
rect 13230 11969 13258 11970
rect 13230 11943 13231 11969
rect 13231 11943 13257 11969
rect 13257 11943 13258 11969
rect 13230 11942 13258 11943
rect 12222 11326 12250 11354
rect 12950 11270 12978 11298
rect 12222 11241 12250 11242
rect 12222 11215 12223 11241
rect 12223 11215 12249 11241
rect 12249 11215 12250 11241
rect 12222 11214 12250 11215
rect 12278 11185 12306 11186
rect 12278 11159 12279 11185
rect 12279 11159 12305 11185
rect 12305 11159 12306 11185
rect 12278 11158 12306 11159
rect 12502 11158 12530 11186
rect 12894 11214 12922 11242
rect 12726 10737 12754 10738
rect 12726 10711 12727 10737
rect 12727 10711 12753 10737
rect 12753 10711 12754 10737
rect 12726 10710 12754 10711
rect 12502 10374 12530 10402
rect 12278 10038 12306 10066
rect 12054 9617 12082 9618
rect 12054 9591 12055 9617
rect 12055 9591 12081 9617
rect 12081 9591 12082 9617
rect 12054 9590 12082 9591
rect 10878 8918 10906 8946
rect 11046 8470 11074 8498
rect 11326 8862 11354 8890
rect 11326 8526 11354 8554
rect 11214 8441 11242 8442
rect 11214 8415 11215 8441
rect 11215 8415 11241 8441
rect 11241 8415 11242 8441
rect 11214 8414 11242 8415
rect 10878 8358 10906 8386
rect 9422 7657 9450 7658
rect 9422 7631 9423 7657
rect 9423 7631 9449 7657
rect 9449 7631 9450 7657
rect 9422 7630 9450 7631
rect 9310 7601 9338 7602
rect 9310 7575 9311 7601
rect 9311 7575 9337 7601
rect 9337 7575 9338 7601
rect 9310 7574 9338 7575
rect 11382 7630 11410 7658
rect 11606 9086 11634 9114
rect 11774 9422 11802 9450
rect 12222 9534 12250 9562
rect 12390 9702 12418 9730
rect 12558 10345 12586 10346
rect 12558 10319 12559 10345
rect 12559 10319 12585 10345
rect 12585 10319 12586 10345
rect 12558 10318 12586 10319
rect 12558 9982 12586 10010
rect 12950 11129 12978 11130
rect 12950 11103 12951 11129
rect 12951 11103 12977 11129
rect 12977 11103 12978 11129
rect 12950 11102 12978 11103
rect 13566 11102 13594 11130
rect 12838 9590 12866 9618
rect 12390 9225 12418 9226
rect 12390 9199 12391 9225
rect 12391 9199 12417 9225
rect 12417 9199 12418 9225
rect 12390 9198 12418 9199
rect 12950 9225 12978 9226
rect 12950 9199 12951 9225
rect 12951 9199 12977 9225
rect 12977 9199 12978 9225
rect 12950 9198 12978 9199
rect 11774 8862 11802 8890
rect 12782 9086 12810 9114
rect 12670 8833 12698 8834
rect 12670 8807 12671 8833
rect 12671 8807 12697 8833
rect 12697 8807 12698 8833
rect 12670 8806 12698 8807
rect 11774 8694 11802 8722
rect 13062 10486 13090 10514
rect 13566 10513 13594 10514
rect 13566 10487 13567 10513
rect 13567 10487 13593 10513
rect 13593 10487 13594 10513
rect 13566 10486 13594 10487
rect 14350 12334 14378 12362
rect 14182 11633 14210 11634
rect 14182 11607 14183 11633
rect 14183 11607 14209 11633
rect 14209 11607 14210 11633
rect 14182 11606 14210 11607
rect 14070 11577 14098 11578
rect 14070 11551 14071 11577
rect 14071 11551 14097 11577
rect 14097 11551 14098 11577
rect 14070 11550 14098 11551
rect 20006 13118 20034 13146
rect 18942 13062 18970 13090
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 20006 12782 20034 12810
rect 14742 12697 14770 12698
rect 14742 12671 14743 12697
rect 14743 12671 14769 12697
rect 14769 12671 14770 12697
rect 14742 12670 14770 12671
rect 14686 12334 14714 12362
rect 15022 12361 15050 12362
rect 15022 12335 15023 12361
rect 15023 12335 15049 12361
rect 15049 12335 15050 12361
rect 15022 12334 15050 12335
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 18830 11969 18858 11970
rect 18830 11943 18831 11969
rect 18831 11943 18857 11969
rect 18857 11943 18858 11969
rect 18830 11942 18858 11943
rect 20006 11774 20034 11802
rect 14742 11633 14770 11634
rect 14742 11607 14743 11633
rect 14743 11607 14769 11633
rect 14769 11607 14770 11633
rect 14742 11606 14770 11607
rect 14406 11494 14434 11522
rect 14014 11241 14042 11242
rect 14014 11215 14015 11241
rect 14015 11215 14041 11241
rect 14041 11215 14042 11241
rect 14014 11214 14042 11215
rect 14126 11185 14154 11186
rect 14126 11159 14127 11185
rect 14127 11159 14153 11185
rect 14153 11159 14154 11185
rect 14126 11158 14154 11159
rect 14294 11073 14322 11074
rect 14294 11047 14295 11073
rect 14295 11047 14321 11073
rect 14321 11047 14322 11073
rect 14294 11046 14322 11047
rect 14966 11550 14994 11578
rect 18830 11577 18858 11578
rect 18830 11551 18831 11577
rect 18831 11551 18857 11577
rect 18857 11551 18858 11577
rect 18830 11550 18858 11551
rect 16030 11521 16058 11522
rect 16030 11495 16031 11521
rect 16031 11495 16057 11521
rect 16057 11495 16058 11521
rect 16030 11494 16058 11495
rect 15806 11438 15834 11466
rect 20006 11465 20034 11466
rect 20006 11439 20007 11465
rect 20007 11439 20033 11465
rect 20033 11439 20034 11465
rect 20006 11438 20034 11439
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 13454 10401 13482 10402
rect 13454 10375 13455 10401
rect 13455 10375 13481 10401
rect 13481 10375 13482 10401
rect 13454 10374 13482 10375
rect 13398 10038 13426 10066
rect 13062 9814 13090 9842
rect 13398 9814 13426 9842
rect 14182 10374 14210 10402
rect 13118 9169 13146 9170
rect 13118 9143 13119 9169
rect 13119 9143 13145 9169
rect 13145 9143 13146 9169
rect 13118 9142 13146 9143
rect 12950 8497 12978 8498
rect 12950 8471 12951 8497
rect 12951 8471 12977 8497
rect 12977 8471 12978 8497
rect 12950 8470 12978 8471
rect 12894 8414 12922 8442
rect 13062 8414 13090 8442
rect 11886 7657 11914 7658
rect 11886 7631 11887 7657
rect 11887 7631 11913 7657
rect 11913 7631 11914 7657
rect 11886 7630 11914 7631
rect 13510 9926 13538 9954
rect 13958 9478 13986 9506
rect 13790 9310 13818 9338
rect 13622 9225 13650 9226
rect 13622 9199 13623 9225
rect 13623 9199 13649 9225
rect 13649 9199 13650 9225
rect 13622 9198 13650 9199
rect 14014 9310 14042 9338
rect 13678 9086 13706 9114
rect 13398 8526 13426 8554
rect 13958 8750 13986 8778
rect 13958 8470 13986 8498
rect 13846 8441 13874 8442
rect 13846 8415 13847 8441
rect 13847 8415 13873 8441
rect 13873 8415 13874 8441
rect 13846 8414 13874 8415
rect 13286 8246 13314 8274
rect 8078 7238 8106 7266
rect 8918 7265 8946 7266
rect 8918 7239 8919 7265
rect 8919 7239 8945 7265
rect 8945 7239 8946 7265
rect 8918 7238 8946 7239
rect 10710 7265 10738 7266
rect 10710 7239 10711 7265
rect 10711 7239 10737 7265
rect 10737 7239 10738 7265
rect 10710 7238 10738 7239
rect 11158 7265 11186 7266
rect 11158 7239 11159 7265
rect 11159 7239 11185 7265
rect 11185 7239 11186 7265
rect 11158 7238 11186 7239
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 15806 11214 15834 11242
rect 14574 10038 14602 10066
rect 14294 9870 14322 9898
rect 14126 9478 14154 9506
rect 14070 9142 14098 9170
rect 14070 8806 14098 8834
rect 14126 9225 14154 9226
rect 14126 9199 14127 9225
rect 14127 9199 14153 9225
rect 14153 9199 14154 9225
rect 14126 9198 14154 9199
rect 14350 9534 14378 9562
rect 14742 11046 14770 11074
rect 14798 11102 14826 11130
rect 20006 10766 20034 10794
rect 18830 10710 18858 10738
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 14854 10401 14882 10402
rect 14854 10375 14855 10401
rect 14855 10375 14881 10401
rect 14881 10375 14882 10401
rect 14854 10374 14882 10375
rect 14630 9310 14658 9338
rect 14686 9926 14714 9954
rect 14574 9198 14602 9226
rect 14574 8833 14602 8834
rect 14574 8807 14575 8833
rect 14575 8807 14601 8833
rect 14601 8807 14602 8833
rect 14574 8806 14602 8807
rect 15414 9897 15442 9898
rect 15414 9871 15415 9897
rect 15415 9871 15441 9897
rect 15441 9871 15442 9897
rect 15414 9870 15442 9871
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 15470 9646 15498 9674
rect 16030 9673 16058 9674
rect 16030 9647 16031 9673
rect 16031 9647 16057 9673
rect 16057 9647 16058 9673
rect 16030 9646 16058 9647
rect 20006 10094 20034 10122
rect 18830 9646 18858 9674
rect 14966 9561 14994 9562
rect 14966 9535 14967 9561
rect 14967 9535 14993 9561
rect 14993 9535 14994 9561
rect 14966 9534 14994 9535
rect 14350 8526 14378 8554
rect 14686 8526 14714 8554
rect 14294 8414 14322 8442
rect 14238 7993 14266 7994
rect 14238 7967 14239 7993
rect 14239 7967 14265 7993
rect 14265 7967 14266 7993
rect 14238 7966 14266 7967
rect 14630 8022 14658 8050
rect 14518 7993 14546 7994
rect 14518 7967 14519 7993
rect 14519 7967 14545 7993
rect 14545 7967 14546 7993
rect 14518 7966 14546 7967
rect 15078 8638 15106 8666
rect 15526 8638 15554 8666
rect 15022 8526 15050 8554
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 20006 9113 20034 9114
rect 20006 9087 20007 9113
rect 20007 9087 20033 9113
rect 20033 9087 20034 9113
rect 20006 9086 20034 9087
rect 18942 8638 18970 8666
rect 15526 8441 15554 8442
rect 15526 8415 15527 8441
rect 15527 8415 15553 8441
rect 15553 8415 15554 8441
rect 15526 8414 15554 8415
rect 15022 8358 15050 8386
rect 15302 8385 15330 8386
rect 15302 8359 15303 8385
rect 15303 8359 15329 8385
rect 15329 8359 15330 8385
rect 15302 8358 15330 8359
rect 20006 8414 20034 8442
rect 18830 8358 18858 8386
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 19950 8078 19978 8106
rect 15022 8049 15050 8050
rect 15022 8023 15023 8049
rect 15023 8023 15049 8049
rect 15049 8023 15050 8049
rect 15022 8022 15050 8023
rect 18830 8049 18858 8050
rect 18830 8023 18831 8049
rect 18831 8023 18857 8049
rect 18857 8023 18858 8049
rect 18830 8022 18858 8023
rect 15134 7937 15162 7938
rect 15134 7911 15135 7937
rect 15135 7911 15161 7937
rect 15161 7911 15162 7937
rect 15134 7910 15162 7911
rect 20006 7742 20034 7770
rect 14686 7630 14714 7658
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 12670 7238 12698 7266
rect 12838 7265 12866 7266
rect 12838 7239 12839 7265
rect 12839 7239 12865 7265
rect 12865 7239 12866 7265
rect 12838 7238 12866 7239
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 12110 1806 12138 1834
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 11433 19110 11438 19138
rect 11466 19110 12782 19138
rect 12810 19110 12815 19138
rect 8969 18998 8974 19026
rect 9002 18998 9310 19026
rect 9338 18998 9343 19026
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 9753 18718 9758 18746
rect 9786 18718 10374 18746
rect 10402 18718 10407 18746
rect 12105 18718 12110 18746
rect 12138 18718 13118 18746
rect 13146 18718 13151 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 8073 18326 8078 18354
rect 8106 18326 8694 18354
rect 8722 18326 8727 18354
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 11489 14014 11494 14042
rect 11522 14014 12278 14042
rect 12306 14014 12311 14042
rect 10481 13790 10486 13818
rect 10514 13790 11494 13818
rect 11522 13790 11527 13818
rect 11265 13734 11270 13762
rect 11298 13734 11550 13762
rect 11578 13734 11583 13762
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 11769 13566 11774 13594
rect 11802 13566 12278 13594
rect 12306 13566 12614 13594
rect 12642 13566 12647 13594
rect 10873 13510 10878 13538
rect 10906 13510 12502 13538
rect 12530 13510 13006 13538
rect 13034 13510 13039 13538
rect 0 13482 400 13496
rect 0 13454 2086 13482
rect 2114 13454 2119 13482
rect 0 13440 400 13454
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 9081 13174 9086 13202
rect 9114 13174 9394 13202
rect 9366 13146 9394 13174
rect 20600 13146 21000 13160
rect 2137 13118 2142 13146
rect 2170 13118 6062 13146
rect 6090 13118 6095 13146
rect 9361 13118 9366 13146
rect 9394 13118 9399 13146
rect 14625 13118 14630 13146
rect 14658 13118 18830 13146
rect 18858 13118 18863 13146
rect 20001 13118 20006 13146
rect 20034 13118 21000 13146
rect 20600 13104 21000 13118
rect 7177 13062 7182 13090
rect 7210 13062 7966 13090
rect 7994 13062 7999 13090
rect 14177 13062 14182 13090
rect 14210 13062 14462 13090
rect 14490 13062 18942 13090
rect 18970 13062 18975 13090
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 0 12810 400 12824
rect 20600 12810 21000 12824
rect 0 12782 966 12810
rect 994 12782 999 12810
rect 7854 12782 7910 12810
rect 7938 12782 7943 12810
rect 8241 12782 8246 12810
rect 8274 12782 9310 12810
rect 9338 12782 9343 12810
rect 20001 12782 20006 12810
rect 20034 12782 21000 12810
rect 0 12768 400 12782
rect 7345 12726 7350 12754
rect 7378 12726 7574 12754
rect 7602 12726 7607 12754
rect 6057 12670 6062 12698
rect 6090 12670 7238 12698
rect 7266 12670 7271 12698
rect 7854 12642 7882 12782
rect 20600 12768 21000 12782
rect 9361 12726 9366 12754
rect 9394 12726 10318 12754
rect 10346 12726 10351 12754
rect 11825 12726 11830 12754
rect 11858 12726 14238 12754
rect 14266 12726 14574 12754
rect 14602 12726 14607 12754
rect 9473 12670 9478 12698
rect 9506 12670 10262 12698
rect 10290 12670 10934 12698
rect 10962 12670 10967 12698
rect 13953 12670 13958 12698
rect 13986 12670 14742 12698
rect 14770 12670 14775 12698
rect 7177 12614 7182 12642
rect 7210 12614 7882 12642
rect 9809 12614 9814 12642
rect 9842 12614 11214 12642
rect 11242 12614 11247 12642
rect 7457 12558 7462 12586
rect 7490 12558 7574 12586
rect 7546 12418 7574 12558
rect 7854 12530 7882 12614
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 7849 12502 7854 12530
rect 7882 12502 7887 12530
rect 11265 12446 11270 12474
rect 11298 12446 11886 12474
rect 11914 12446 11919 12474
rect 7546 12390 9590 12418
rect 9618 12390 9623 12418
rect 12049 12390 12054 12418
rect 12082 12390 13006 12418
rect 13034 12390 13039 12418
rect 8409 12334 8414 12362
rect 8442 12334 9646 12362
rect 9674 12334 9679 12362
rect 13057 12334 13062 12362
rect 13090 12334 13342 12362
rect 13370 12334 14350 12362
rect 14378 12334 14686 12362
rect 14714 12334 15022 12362
rect 15050 12334 15055 12362
rect 6449 12278 6454 12306
rect 6482 12278 6846 12306
rect 6874 12278 7070 12306
rect 7098 12278 7518 12306
rect 7546 12278 7742 12306
rect 7770 12278 7775 12306
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 13001 12054 13006 12082
rect 13034 12054 15974 12082
rect 15946 11970 15974 12054
rect 2137 11942 2142 11970
rect 2170 11942 4214 11970
rect 8801 11942 8806 11970
rect 8834 11942 9198 11970
rect 9226 11942 9646 11970
rect 9674 11942 9679 11970
rect 11601 11942 11606 11970
rect 11634 11942 13230 11970
rect 13258 11942 13263 11970
rect 15946 11942 18830 11970
rect 18858 11942 18863 11970
rect 4186 11914 4214 11942
rect 4186 11886 4998 11914
rect 5026 11886 6790 11914
rect 6818 11886 6823 11914
rect 7065 11886 7070 11914
rect 7098 11886 11774 11914
rect 11802 11886 11807 11914
rect 7737 11830 7742 11858
rect 7770 11830 8358 11858
rect 8386 11830 8391 11858
rect 0 11802 400 11816
rect 20600 11802 21000 11816
rect 0 11774 966 11802
rect 994 11774 999 11802
rect 8241 11774 8246 11802
rect 8274 11774 8638 11802
rect 8666 11774 8671 11802
rect 10257 11774 10262 11802
rect 10290 11774 11214 11802
rect 11242 11774 11247 11802
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 0 11760 400 11774
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 20600 11760 21000 11774
rect 8409 11718 8414 11746
rect 8442 11718 8862 11746
rect 8890 11718 8895 11746
rect 10201 11662 10206 11690
rect 10234 11662 11886 11690
rect 11914 11662 11919 11690
rect 8689 11606 8694 11634
rect 8722 11606 9926 11634
rect 9954 11606 9959 11634
rect 10649 11606 10654 11634
rect 10682 11606 10990 11634
rect 11018 11606 11023 11634
rect 11545 11606 11550 11634
rect 11578 11606 11998 11634
rect 12026 11606 12031 11634
rect 14177 11606 14182 11634
rect 14210 11606 14742 11634
rect 14770 11606 14775 11634
rect 9081 11550 9086 11578
rect 9114 11550 10430 11578
rect 10458 11550 10463 11578
rect 14065 11550 14070 11578
rect 14098 11550 14966 11578
rect 14994 11550 14999 11578
rect 18825 11550 18830 11578
rect 18858 11550 18863 11578
rect 2137 11494 2142 11522
rect 2170 11494 6846 11522
rect 6874 11494 8022 11522
rect 8050 11494 8055 11522
rect 9473 11494 9478 11522
rect 9506 11494 10542 11522
rect 10570 11494 10575 11522
rect 14401 11494 14406 11522
rect 14434 11494 16030 11522
rect 16058 11494 16063 11522
rect 0 11466 400 11480
rect 18830 11466 18858 11550
rect 20600 11466 21000 11480
rect 0 11438 966 11466
rect 994 11438 999 11466
rect 9641 11438 9646 11466
rect 9674 11438 10038 11466
rect 10066 11438 10071 11466
rect 15801 11438 15806 11466
rect 15834 11438 18858 11466
rect 20001 11438 20006 11466
rect 20034 11438 21000 11466
rect 0 11424 400 11438
rect 20600 11424 21000 11438
rect 7793 11382 7798 11410
rect 7826 11382 7910 11410
rect 7938 11382 8694 11410
rect 8722 11382 8727 11410
rect 9193 11382 9198 11410
rect 9226 11382 10206 11410
rect 10234 11382 10239 11410
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 10369 11326 10374 11354
rect 10402 11326 12222 11354
rect 12250 11326 12255 11354
rect 6393 11270 6398 11298
rect 6426 11270 8414 11298
rect 8442 11270 8447 11298
rect 9809 11270 9814 11298
rect 9842 11270 12950 11298
rect 12978 11270 12983 11298
rect 12217 11214 12222 11242
rect 12250 11214 12894 11242
rect 12922 11214 12927 11242
rect 14009 11214 14014 11242
rect 14042 11214 15806 11242
rect 15834 11214 15839 11242
rect 8465 11158 8470 11186
rect 8498 11158 8694 11186
rect 8722 11158 9142 11186
rect 9170 11158 9175 11186
rect 10425 11158 10430 11186
rect 10458 11158 12278 11186
rect 12306 11158 12502 11186
rect 12530 11158 14126 11186
rect 14154 11158 14159 11186
rect 12945 11102 12950 11130
rect 12978 11102 13566 11130
rect 13594 11102 14798 11130
rect 14826 11102 14831 11130
rect 7961 11046 7966 11074
rect 7994 11046 8750 11074
rect 8778 11046 8783 11074
rect 14289 11046 14294 11074
rect 14322 11046 14742 11074
rect 14770 11046 14775 11074
rect 11041 10990 11046 11018
rect 11074 10990 11662 11018
rect 11690 10990 11695 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 10089 10934 10094 10962
rect 10122 10934 10542 10962
rect 10570 10934 10575 10962
rect 10649 10934 10654 10962
rect 10682 10934 10934 10962
rect 10962 10934 11382 10962
rect 11410 10934 11415 10962
rect 6393 10878 6398 10906
rect 6426 10878 7126 10906
rect 7154 10878 7630 10906
rect 7658 10878 7663 10906
rect 7737 10878 7742 10906
rect 7770 10878 8918 10906
rect 8946 10878 8951 10906
rect 6897 10822 6902 10850
rect 6930 10822 7574 10850
rect 7602 10822 7607 10850
rect 8409 10822 8414 10850
rect 8442 10822 8974 10850
rect 9002 10822 9007 10850
rect 0 10794 400 10808
rect 20600 10794 21000 10808
rect 0 10766 966 10794
rect 994 10766 999 10794
rect 4186 10766 4942 10794
rect 4970 10766 6566 10794
rect 6594 10766 6599 10794
rect 6785 10766 6790 10794
rect 6818 10766 9310 10794
rect 9338 10766 9758 10794
rect 9786 10766 9791 10794
rect 20001 10766 20006 10794
rect 20034 10766 21000 10794
rect 0 10752 400 10766
rect 4186 10738 4214 10766
rect 20600 10752 21000 10766
rect 2137 10710 2142 10738
rect 2170 10710 4214 10738
rect 5833 10710 5838 10738
rect 5866 10710 6734 10738
rect 6762 10710 6767 10738
rect 8409 10710 8414 10738
rect 8442 10710 8806 10738
rect 8834 10710 8839 10738
rect 12721 10710 12726 10738
rect 12754 10710 18830 10738
rect 18858 10710 18863 10738
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 9025 10542 9030 10570
rect 9058 10542 9310 10570
rect 9338 10542 9343 10570
rect 2081 10486 2086 10514
rect 2114 10486 4214 10514
rect 8913 10486 8918 10514
rect 8946 10486 10038 10514
rect 10066 10486 10071 10514
rect 13057 10486 13062 10514
rect 13090 10486 13566 10514
rect 13594 10486 13599 10514
rect 4186 10402 4214 10486
rect 4186 10374 10430 10402
rect 10458 10374 10654 10402
rect 10682 10374 10687 10402
rect 12497 10374 12502 10402
rect 12530 10374 13454 10402
rect 13482 10374 13487 10402
rect 14177 10374 14182 10402
rect 14210 10374 14854 10402
rect 14882 10374 14887 10402
rect 11321 10318 11326 10346
rect 11354 10318 12558 10346
rect 12586 10318 12591 10346
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 9025 10150 9030 10178
rect 9058 10150 9366 10178
rect 9394 10150 9399 10178
rect 0 10122 400 10136
rect 20600 10122 21000 10136
rect 0 10094 966 10122
rect 994 10094 999 10122
rect 20001 10094 20006 10122
rect 20034 10094 21000 10122
rect 0 10080 400 10094
rect 20600 10080 21000 10094
rect 4186 10038 6174 10066
rect 6202 10038 6207 10066
rect 6841 10038 6846 10066
rect 6874 10038 9254 10066
rect 9282 10038 9287 10066
rect 10257 10038 10262 10066
rect 10290 10038 11270 10066
rect 11298 10038 12278 10066
rect 12306 10038 12311 10066
rect 13393 10038 13398 10066
rect 13426 10038 14574 10066
rect 14602 10038 14607 10066
rect 4186 10010 4214 10038
rect 2137 9982 2142 10010
rect 2170 9982 4214 10010
rect 6729 9982 6734 10010
rect 6762 9982 7182 10010
rect 7210 9982 7215 10010
rect 9753 9982 9758 10010
rect 9786 9982 10150 10010
rect 10178 9982 10654 10010
rect 10682 9982 10687 10010
rect 11657 9982 11662 10010
rect 11690 9982 12558 10010
rect 12586 9982 12591 10010
rect 5721 9926 5726 9954
rect 5754 9926 6678 9954
rect 6706 9926 6711 9954
rect 9529 9926 9534 9954
rect 9562 9926 9814 9954
rect 9842 9926 10318 9954
rect 10346 9926 11326 9954
rect 11354 9926 11359 9954
rect 11433 9926 11438 9954
rect 11466 9926 13510 9954
rect 13538 9926 14686 9954
rect 14714 9926 14719 9954
rect 961 9870 966 9898
rect 994 9870 999 9898
rect 2081 9870 2086 9898
rect 2114 9870 4830 9898
rect 4858 9870 6286 9898
rect 6314 9870 6319 9898
rect 6617 9870 6622 9898
rect 6650 9870 7014 9898
rect 7042 9870 11606 9898
rect 11634 9870 11639 9898
rect 14289 9870 14294 9898
rect 14322 9870 15414 9898
rect 15442 9870 15447 9898
rect 0 9786 400 9800
rect 966 9786 994 9870
rect 9137 9814 9142 9842
rect 9170 9814 9814 9842
rect 9842 9814 10990 9842
rect 11018 9814 11023 9842
rect 11657 9814 11662 9842
rect 11690 9814 11886 9842
rect 11914 9814 13062 9842
rect 13090 9814 13398 9842
rect 13426 9814 13431 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 0 9758 994 9786
rect 9361 9758 9366 9786
rect 9394 9758 11718 9786
rect 11746 9758 11751 9786
rect 0 9744 400 9758
rect 9249 9702 9254 9730
rect 9282 9702 10598 9730
rect 10626 9702 12390 9730
rect 12418 9702 12423 9730
rect 8969 9646 8974 9674
rect 9002 9646 9702 9674
rect 9730 9646 9735 9674
rect 11825 9646 11830 9674
rect 11858 9646 11863 9674
rect 15465 9646 15470 9674
rect 15498 9646 16030 9674
rect 16058 9646 18830 9674
rect 18858 9646 18863 9674
rect 11830 9618 11858 9646
rect 6897 9590 6902 9618
rect 6930 9590 7742 9618
rect 7770 9590 7775 9618
rect 9193 9590 9198 9618
rect 9226 9590 11494 9618
rect 11522 9590 11527 9618
rect 11830 9590 12054 9618
rect 12082 9590 12838 9618
rect 12866 9590 12871 9618
rect 11494 9562 11522 9590
rect 6841 9534 6846 9562
rect 6874 9534 7070 9562
rect 7098 9534 7103 9562
rect 8745 9534 8750 9562
rect 8778 9534 9310 9562
rect 9338 9534 9343 9562
rect 11494 9534 12222 9562
rect 12250 9534 12255 9562
rect 14345 9534 14350 9562
rect 14378 9534 14966 9562
rect 14994 9534 14999 9562
rect 5945 9478 5950 9506
rect 5978 9478 6902 9506
rect 6930 9478 6935 9506
rect 11265 9478 11270 9506
rect 11298 9478 13958 9506
rect 13986 9478 14126 9506
rect 14154 9478 14159 9506
rect 0 9450 400 9464
rect 0 9422 966 9450
rect 994 9422 999 9450
rect 10257 9422 10262 9450
rect 10290 9422 11774 9450
rect 11802 9422 11807 9450
rect 0 9408 400 9422
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 7177 9310 7182 9338
rect 7210 9310 7966 9338
rect 7994 9310 7999 9338
rect 9697 9310 9702 9338
rect 9730 9310 9926 9338
rect 9954 9310 9959 9338
rect 13785 9310 13790 9338
rect 13818 9310 14014 9338
rect 14042 9310 14630 9338
rect 14658 9310 14663 9338
rect 9361 9198 9366 9226
rect 9394 9198 9646 9226
rect 9674 9198 10038 9226
rect 10066 9198 11438 9226
rect 11466 9198 11471 9226
rect 12385 9198 12390 9226
rect 12418 9198 12950 9226
rect 12978 9198 13622 9226
rect 13650 9198 13655 9226
rect 14121 9198 14126 9226
rect 14154 9198 14574 9226
rect 14602 9198 14607 9226
rect 2137 9142 2142 9170
rect 2170 9142 4886 9170
rect 4914 9142 6510 9170
rect 6538 9142 6543 9170
rect 9921 9142 9926 9170
rect 9954 9142 10430 9170
rect 10458 9142 11102 9170
rect 11130 9142 11135 9170
rect 13113 9142 13118 9170
rect 13146 9142 14070 9170
rect 14098 9142 14103 9170
rect 20600 9114 21000 9128
rect 10089 9086 10094 9114
rect 10122 9086 10766 9114
rect 10794 9086 11606 9114
rect 11634 9086 11639 9114
rect 12777 9086 12782 9114
rect 12810 9086 13678 9114
rect 13706 9086 13711 9114
rect 20001 9086 20006 9114
rect 20034 9086 21000 9114
rect 20600 9072 21000 9086
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 9347 8918 9366 8946
rect 9394 8918 9399 8946
rect 9697 8918 9702 8946
rect 9730 8918 10878 8946
rect 10906 8918 10911 8946
rect 7401 8862 7406 8890
rect 7434 8862 7686 8890
rect 7714 8862 8750 8890
rect 8778 8862 8783 8890
rect 9305 8862 9310 8890
rect 9338 8862 10766 8890
rect 10794 8862 10799 8890
rect 11321 8862 11326 8890
rect 11354 8862 11774 8890
rect 11802 8862 11807 8890
rect 2137 8806 2142 8834
rect 2170 8806 5950 8834
rect 5978 8806 7238 8834
rect 7266 8806 7271 8834
rect 8297 8806 8302 8834
rect 8330 8806 9870 8834
rect 9898 8806 12670 8834
rect 12698 8806 12703 8834
rect 14065 8806 14070 8834
rect 14098 8806 14574 8834
rect 14602 8806 14607 8834
rect 15946 8806 18830 8834
rect 18858 8806 18863 8834
rect 15946 8778 15974 8806
rect 8185 8750 8190 8778
rect 8218 8750 8862 8778
rect 8890 8750 8895 8778
rect 9025 8750 9030 8778
rect 9058 8750 10654 8778
rect 10682 8750 10687 8778
rect 13953 8750 13958 8778
rect 13986 8750 15974 8778
rect 8969 8694 8974 8722
rect 9002 8694 9254 8722
rect 9282 8694 10150 8722
rect 10178 8694 10183 8722
rect 10761 8694 10766 8722
rect 10794 8694 11774 8722
rect 11802 8694 11807 8722
rect 15073 8638 15078 8666
rect 15106 8638 15526 8666
rect 15554 8638 18942 8666
rect 18970 8638 18975 8666
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 7289 8582 7294 8610
rect 7322 8582 7574 8610
rect 9641 8582 9646 8610
rect 9674 8582 9814 8610
rect 9842 8582 9847 8610
rect 7546 8554 7574 8582
rect 9814 8554 9842 8582
rect 7546 8526 8078 8554
rect 8106 8526 9702 8554
rect 9730 8526 9735 8554
rect 9814 8526 10430 8554
rect 10458 8526 11326 8554
rect 11354 8526 11359 8554
rect 12838 8526 13398 8554
rect 13426 8526 13431 8554
rect 14345 8526 14350 8554
rect 14378 8526 14686 8554
rect 14714 8526 15022 8554
rect 15050 8526 15055 8554
rect 7009 8470 7014 8498
rect 7042 8470 7574 8498
rect 7602 8470 7607 8498
rect 9291 8470 9310 8498
rect 9338 8470 9343 8498
rect 11041 8470 11046 8498
rect 11074 8470 12250 8498
rect 0 8442 400 8456
rect 12222 8442 12250 8470
rect 12838 8442 12866 8526
rect 12945 8470 12950 8498
rect 12978 8470 13958 8498
rect 13986 8470 13991 8498
rect 20600 8442 21000 8456
rect 0 8414 966 8442
rect 994 8414 999 8442
rect 2137 8414 2142 8442
rect 2170 8414 5894 8442
rect 5922 8414 5927 8442
rect 6505 8414 6510 8442
rect 6538 8414 6790 8442
rect 6818 8414 7406 8442
rect 7434 8414 7439 8442
rect 9403 8414 9422 8442
rect 9450 8414 9455 8442
rect 10878 8414 11214 8442
rect 11242 8414 11247 8442
rect 12222 8414 12894 8442
rect 12922 8414 12927 8442
rect 13057 8414 13062 8442
rect 13090 8414 13846 8442
rect 13874 8414 14294 8442
rect 14322 8414 15526 8442
rect 15554 8414 15559 8442
rect 20001 8414 20006 8442
rect 20034 8414 21000 8442
rect 0 8400 400 8414
rect 10878 8386 10906 8414
rect 20600 8400 21000 8414
rect 7177 8358 7182 8386
rect 7210 8358 7630 8386
rect 7658 8358 7663 8386
rect 9865 8358 9870 8386
rect 9898 8358 10094 8386
rect 10122 8358 10542 8386
rect 10570 8358 10878 8386
rect 10906 8358 10911 8386
rect 15017 8358 15022 8386
rect 15050 8358 15302 8386
rect 15330 8358 18830 8386
rect 18858 8358 18863 8386
rect 9529 8246 9534 8274
rect 9562 8246 13286 8274
rect 13314 8246 13319 8274
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 0 8106 400 8120
rect 20600 8106 21000 8120
rect 0 8078 966 8106
rect 994 8078 999 8106
rect 19945 8078 19950 8106
rect 19978 8078 21000 8106
rect 0 8064 400 8078
rect 20600 8064 21000 8078
rect 9417 8022 9422 8050
rect 9450 8022 9870 8050
rect 9898 8022 9903 8050
rect 14625 8022 14630 8050
rect 14658 8022 15022 8050
rect 15050 8022 15055 8050
rect 15946 8022 18830 8050
rect 18858 8022 18863 8050
rect 5889 7966 5894 7994
rect 5922 7966 7630 7994
rect 7658 7966 7663 7994
rect 9347 7966 9366 7994
rect 9394 7966 9399 7994
rect 14233 7966 14238 7994
rect 14266 7966 14518 7994
rect 14546 7966 14551 7994
rect 15946 7938 15974 8022
rect 15129 7910 15134 7938
rect 15162 7910 15974 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 20600 7770 21000 7784
rect 20001 7742 20006 7770
rect 20034 7742 21000 7770
rect 20600 7728 21000 7742
rect 7905 7686 7910 7714
rect 7938 7686 9534 7714
rect 9562 7686 9567 7714
rect 9403 7630 9422 7658
rect 9450 7630 9455 7658
rect 11377 7630 11382 7658
rect 11410 7630 11886 7658
rect 11914 7630 14686 7658
rect 14714 7630 14719 7658
rect 8689 7574 8694 7602
rect 8722 7574 9310 7602
rect 9338 7574 9343 7602
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 7345 7238 7350 7266
rect 7378 7238 7686 7266
rect 7714 7238 8078 7266
rect 8106 7238 8918 7266
rect 8946 7238 10710 7266
rect 10738 7238 10743 7266
rect 11153 7238 11158 7266
rect 11186 7238 12670 7266
rect 12698 7238 12838 7266
rect 12866 7238 12871 7266
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 12105 1806 12110 1834
rect 12138 1806 12782 1834
rect 12810 1806 12815 1834
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 9310 10766 9338 10794
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9366 8918 9394 8946
rect 9310 8862 9338 8890
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 9310 8470 9338 8498
rect 9422 8414 9450 8442
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9422 8022 9450 8050
rect 9366 7966 9394 7994
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 9422 7630 9450 7658
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 9310 10794 9338 10799
rect 9310 8890 9338 10766
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9310 8498 9338 8862
rect 9310 8465 9338 8470
rect 9366 8946 9394 8951
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 9366 7994 9394 8918
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9366 7961 9394 7966
rect 9422 8442 9450 8447
rect 9422 8050 9450 8414
rect 9422 7658 9450 8022
rect 9422 7625 9450 7630
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10248 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_
timestamp 1698175906
transform -1 0 9576 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1698175906
transform 1 0 9128 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11368 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11704 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12824 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9240 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _119_
timestamp 1698175906
transform -1 0 10584 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9296 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9296 0 -1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _122_
timestamp 1698175906
transform 1 0 10304 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698175906
transform 1 0 10808 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _124_
timestamp 1698175906
transform 1 0 11032 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _125_
timestamp 1698175906
transform 1 0 10304 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _126_
timestamp 1698175906
transform -1 0 10136 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11200 0 1 11760
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _128_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11760 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _129_
timestamp 1698175906
transform -1 0 11592 0 -1 12544
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _130_
timestamp 1698175906
transform 1 0 11928 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _131_
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _132_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10416 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8960 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _134_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10304 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9072 0 -1 7840
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _136_
timestamp 1698175906
transform -1 0 9800 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _137_
timestamp 1698175906
transform 1 0 9464 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _138_
timestamp 1698175906
transform -1 0 11032 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _139_
timestamp 1698175906
transform -1 0 12040 0 -1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _140_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6440 0 -1 10192
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _141_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5656 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform 1 0 11928 0 -1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _143_
timestamp 1698175906
transform 1 0 12824 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _144_
timestamp 1698175906
transform -1 0 12264 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _145_
timestamp 1698175906
transform 1 0 9800 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _146_
timestamp 1698175906
transform -1 0 8008 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _147_
timestamp 1698175906
transform -1 0 9464 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _148_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9240 0 1 9408
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _149_
timestamp 1698175906
transform -1 0 8904 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _150_
timestamp 1698175906
transform -1 0 9240 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _151_
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _152_
timestamp 1698175906
transform -1 0 11872 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _153_
timestamp 1698175906
transform 1 0 11592 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _154_
timestamp 1698175906
transform -1 0 12264 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _155_
timestamp 1698175906
transform 1 0 11144 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _156_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11984 0 -1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _157_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698175906
transform 1 0 14952 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _159_
timestamp 1698175906
transform -1 0 10472 0 1 8624
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform 1 0 12152 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _161_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12768 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _162_
timestamp 1698175906
transform -1 0 14952 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _163_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9688 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _164_
timestamp 1698175906
transform -1 0 11928 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _165_
timestamp 1698175906
transform -1 0 11928 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _166_
timestamp 1698175906
transform -1 0 11368 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _167_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9016 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _168_
timestamp 1698175906
transform -1 0 14336 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _169_
timestamp 1698175906
transform -1 0 13720 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _170_
timestamp 1698175906
transform -1 0 13104 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _171_
timestamp 1698175906
transform -1 0 12376 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _172_
timestamp 1698175906
transform -1 0 13048 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _173_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9968 0 1 10192
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _174_
timestamp 1698175906
transform -1 0 11648 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _175_
timestamp 1698175906
transform -1 0 10472 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _176_
timestamp 1698175906
transform -1 0 11312 0 1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _178_
timestamp 1698175906
transform -1 0 14056 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _179_
timestamp 1698175906
transform 1 0 13216 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _180_
timestamp 1698175906
transform 1 0 12824 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _181_
timestamp 1698175906
transform 1 0 12376 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _182_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13384 0 1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _183_
timestamp 1698175906
transform -1 0 14280 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _184_
timestamp 1698175906
transform 1 0 13552 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _185_
timestamp 1698175906
transform -1 0 14784 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _186_
timestamp 1698175906
transform -1 0 14336 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _187_
timestamp 1698175906
transform -1 0 15568 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _188_
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _189_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13776 0 1 9408
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _190_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15008 0 1 10192
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _191_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13944 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _192_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _193_
timestamp 1698175906
transform 1 0 13944 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _194_
timestamp 1698175906
transform -1 0 8568 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _195_
timestamp 1698175906
transform -1 0 6944 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _196_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6328 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _197_
timestamp 1698175906
transform -1 0 7840 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _198_
timestamp 1698175906
transform 1 0 6496 0 -1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _199_
timestamp 1698175906
transform 1 0 5768 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _200_
timestamp 1698175906
transform -1 0 9576 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _201_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10080 0 1 9408
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _202_
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _203_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9352 0 -1 13328
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _204_
timestamp 1698175906
transform -1 0 9128 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _205_
timestamp 1698175906
transform 1 0 9576 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _206_
timestamp 1698175906
transform 1 0 7616 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _207_
timestamp 1698175906
transform -1 0 8400 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _208_
timestamp 1698175906
transform -1 0 7840 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _209_
timestamp 1698175906
transform -1 0 7952 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _210_
timestamp 1698175906
transform -1 0 8008 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _211_
timestamp 1698175906
transform 1 0 6440 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _212_
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _213_
timestamp 1698175906
transform -1 0 7504 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _214_
timestamp 1698175906
transform -1 0 7504 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _215_
timestamp 1698175906
transform 1 0 7896 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _216_
timestamp 1698175906
transform -1 0 8904 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _217_
timestamp 1698175906
transform -1 0 8288 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _218_
timestamp 1698175906
transform 1 0 7112 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _219_
timestamp 1698175906
transform -1 0 10472 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _220_
timestamp 1698175906
transform 1 0 7392 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _221_
timestamp 1698175906
transform 1 0 7896 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _222_
timestamp 1698175906
transform 1 0 9184 0 1 12544
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _223_
timestamp 1698175906
transform -1 0 8288 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9576 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform -1 0 6384 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 11480 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform 1 0 8792 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 7168 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 7504 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform -1 0 12880 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 11032 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 14000 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform 1 0 10752 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 12936 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform 1 0 9912 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 13272 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698175906
transform -1 0 14280 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform 1 0 13776 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _240_
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _241_
timestamp 1698175906
transform 1 0 14280 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _242_
timestamp 1698175906
transform -1 0 6552 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _243_
timestamp 1698175906
transform -1 0 6496 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _244_
timestamp 1698175906
transform 1 0 8176 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _245_
timestamp 1698175906
transform -1 0 7504 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _246_
timestamp 1698175906
transform -1 0 6440 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _247_
timestamp 1698175906
transform -1 0 7504 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _248_
timestamp 1698175906
transform -1 0 8400 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _249_
timestamp 1698175906
transform -1 0 7616 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _250_
timestamp 1698175906
transform 1 0 6720 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _251_
timestamp 1698175906
transform 1 0 14896 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _252_
timestamp 1698175906
transform -1 0 6440 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _253_
timestamp 1698175906
transform -1 0 9576 0 -1 14112
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11200 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 6776 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 13216 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 10696 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform -1 0 8904 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 8400 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 12992 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform -1 0 12880 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 15736 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 12488 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 14672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 14280 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform 1 0 9800 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 15008 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform 1 0 14392 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform 1 0 15512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__CLK
timestamp 1698175906
transform 1 0 14280 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__CLK
timestamp 1698175906
transform 1 0 16016 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__CLK
timestamp 1698175906
transform 1 0 7056 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__CLK
timestamp 1698175906
transform 1 0 7112 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__CLK
timestamp 1698175906
transform 1 0 9912 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__CLK
timestamp 1698175906
transform 1 0 7616 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__CLK
timestamp 1698175906
transform 1 0 6440 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__CLK
timestamp 1698175906
transform 1 0 8064 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__CLK
timestamp 1698175906
transform 1 0 8400 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__CLK
timestamp 1698175906
transform 1 0 7728 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__CLK
timestamp 1698175906
transform 1 0 8400 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 11424 0 -1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 12208 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 16128 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 10248 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_144
timestamp 1698175906
transform 1 0 8736 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_147
timestamp 1698175906
transform 1 0 8904 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_179 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10696 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_195 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11592 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_203
timestamp 1698175906
transform 1 0 12040 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1698175906
transform 1 0 12264 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 12376 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_115
timestamp 1698175906
transform 1 0 7112 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 10416 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_181
timestamp 1698175906
transform 1 0 10808 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_214
timestamp 1698175906
transform 1 0 12656 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_218
timestamp 1698175906
transform 1 0 12880 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_234
timestamp 1698175906
transform 1 0 13776 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_242
timestamp 1698175906
transform 1 0 14224 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 14336 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_88
timestamp 1698175906
transform 1 0 5600 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_92
timestamp 1698175906
transform 1 0 5824 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_122
timestamp 1698175906
transform 1 0 7504 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_126
timestamp 1698175906
transform 1 0 7728 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_131
timestamp 1698175906
transform 1 0 8008 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698175906
transform 1 0 8456 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_163
timestamp 1698175906
transform 1 0 9800 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_171
timestamp 1698175906
transform 1 0 10248 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_180
timestamp 1698175906
transform 1 0 10752 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_188
timestamp 1698175906
transform 1 0 11200 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_202
timestamp 1698175906
transform 1 0 11984 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698175906
transform 1 0 12264 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 12376 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_241
timestamp 1698175906
transform 1 0 14168 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_245
timestamp 1698175906
transform 1 0 14392 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698175906
transform 1 0 16184 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 16296 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_111
timestamp 1698175906
transform 1 0 6888 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_113
timestamp 1698175906
transform 1 0 7000 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_128
timestamp 1698175906
transform 1 0 7840 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_144
timestamp 1698175906
transform 1 0 8736 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_148
timestamp 1698175906
transform 1 0 8960 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_150
timestamp 1698175906
transform 1 0 9072 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_167
timestamp 1698175906
transform 1 0 10024 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_185
timestamp 1698175906
transform 1 0 11032 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_218
timestamp 1698175906
transform 1 0 12880 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_222
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_238
timestamp 1698175906
transform 1 0 14000 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 14336 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_252
timestamp 1698175906
transform 1 0 14784 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_260
timestamp 1698175906
transform 1 0 15232 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_292
timestamp 1698175906
transform 1 0 17024 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_308
timestamp 1698175906
transform 1 0 17920 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_312
timestamp 1698175906
transform 1 0 18144 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1698175906
transform 1 0 18256 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 18648 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 2240 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 4032 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 4480 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_88
timestamp 1698175906
transform 1 0 5600 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_92
timestamp 1698175906
transform 1 0 5824 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_130
timestamp 1698175906
transform 1 0 7952 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_134
timestamp 1698175906
transform 1 0 8176 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698175906
transform 1 0 8400 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_150
timestamp 1698175906
transform 1 0 9072 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_152
timestamp 1698175906
transform 1 0 9184 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_167
timestamp 1698175906
transform 1 0 10024 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_171
timestamp 1698175906
transform 1 0 10248 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_178
timestamp 1698175906
transform 1 0 10640 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_180
timestamp 1698175906
transform 1 0 10752 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_193
timestamp 1698175906
transform 1 0 11480 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_201
timestamp 1698175906
transform 1 0 11928 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 12376 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_216
timestamp 1698175906
transform 1 0 12768 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_222
timestamp 1698175906
transform 1 0 13104 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_230
timestamp 1698175906
transform 1 0 13552 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_263
timestamp 1698175906
transform 1 0 15400 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_267
timestamp 1698175906
transform 1 0 15624 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_275
timestamp 1698175906
transform 1 0 16072 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 16296 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_115
timestamp 1698175906
transform 1 0 7112 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_122
timestamp 1698175906
transform 1 0 7504 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_138
timestamp 1698175906
transform 1 0 8400 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_151
timestamp 1698175906
transform 1 0 9128 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_185
timestamp 1698175906
transform 1 0 11032 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_201
timestamp 1698175906
transform 1 0 11928 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_209
timestamp 1698175906
transform 1 0 12376 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_221
timestamp 1698175906
transform 1 0 13048 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_237
timestamp 1698175906
transform 1 0 13944 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_241
timestamp 1698175906
transform 1 0 14168 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_260
timestamp 1698175906
transform 1 0 15232 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_292
timestamp 1698175906
transform 1 0 17024 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_308
timestamp 1698175906
transform 1 0 17920 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_312
timestamp 1698175906
transform 1 0 18144 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698175906
transform 1 0 18256 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_107
timestamp 1698175906
transform 1 0 6664 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_111
timestamp 1698175906
transform 1 0 6888 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_119
timestamp 1698175906
transform 1 0 7336 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_123
timestamp 1698175906
transform 1 0 7560 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_131
timestamp 1698175906
transform 1 0 8008 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 8456 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_150
timestamp 1698175906
transform 1 0 9072 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_160
timestamp 1698175906
transform 1 0 9632 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_201
timestamp 1698175906
transform 1 0 11928 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_235
timestamp 1698175906
transform 1 0 13832 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_237
timestamp 1698175906
transform 1 0 13944 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_267
timestamp 1698175906
transform 1 0 15624 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_271
timestamp 1698175906
transform 1 0 15848 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 16296 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 18256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 18704 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698175906
transform 1 0 2240 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698175906
transform 1 0 2464 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 4536 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_102
timestamp 1698175906
transform 1 0 6384 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698175906
transform 1 0 6496 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_118
timestamp 1698175906
transform 1 0 7280 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_134
timestamp 1698175906
transform 1 0 8176 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_138
timestamp 1698175906
transform 1 0 8400 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_140
timestamp 1698175906
transform 1 0 8512 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_168
timestamp 1698175906
transform 1 0 10080 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_172
timestamp 1698175906
transform 1 0 10304 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_190
timestamp 1698175906
transform 1 0 11312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_200
timestamp 1698175906
transform 1 0 11872 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_223
timestamp 1698175906
transform 1 0 13160 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_225
timestamp 1698175906
transform 1 0 13272 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_276
timestamp 1698175906
transform 1 0 16128 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_308
timestamp 1698175906
transform 1 0 17920 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698175906
transform 1 0 18144 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698175906
transform 1 0 18256 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 2240 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 4032 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 4480 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_88
timestamp 1698175906
transform 1 0 5600 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_93
timestamp 1698175906
transform 1 0 5880 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_112
timestamp 1698175906
transform 1 0 6944 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_128
timestamp 1698175906
transform 1 0 7840 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_136
timestamp 1698175906
transform 1 0 8288 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_148
timestamp 1698175906
transform 1 0 8960 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_175
timestamp 1698175906
transform 1 0 10472 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_203
timestamp 1698175906
transform 1 0 12040 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_207
timestamp 1698175906
transform 1 0 12264 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 12376 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_266
timestamp 1698175906
transform 1 0 15568 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_274
timestamp 1698175906
transform 1 0 16016 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 16240 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 20048 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 20160 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698175906
transform 1 0 2240 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698175906
transform 1 0 2464 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_69
timestamp 1698175906
transform 1 0 4536 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_85
timestamp 1698175906
transform 1 0 5432 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_89
timestamp 1698175906
transform 1 0 5656 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_95
timestamp 1698175906
transform 1 0 5992 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_103
timestamp 1698175906
transform 1 0 6440 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_115
timestamp 1698175906
transform 1 0 7112 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_119
timestamp 1698175906
transform 1 0 7336 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_121
timestamp 1698175906
transform 1 0 7448 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_151
timestamp 1698175906
transform 1 0 9128 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698175906
transform 1 0 10416 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698175906
transform 1 0 14280 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_256
timestamp 1698175906
transform 1 0 15008 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_288
timestamp 1698175906
transform 1 0 16800 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_304
timestamp 1698175906
transform 1 0 17696 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_312
timestamp 1698175906
transform 1 0 18144 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698175906
transform 1 0 18256 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 18648 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_74
timestamp 1698175906
transform 1 0 4816 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_113
timestamp 1698175906
transform 1 0 7000 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_117
timestamp 1698175906
transform 1 0 7224 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_121
timestamp 1698175906
transform 1 0 7448 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_128
timestamp 1698175906
transform 1 0 7840 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698175906
transform 1 0 8288 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_192
timestamp 1698175906
transform 1 0 11424 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_198
timestamp 1698175906
transform 1 0 11760 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698175906
transform 1 0 12208 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_243
timestamp 1698175906
transform 1 0 14280 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_247
timestamp 1698175906
transform 1 0 14504 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 16296 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 20048 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 20160 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 2240 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 2464 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_123
timestamp 1698175906
transform 1 0 7560 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_127
timestamp 1698175906
transform 1 0 7784 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_161
timestamp 1698175906
transform 1 0 9688 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_163
timestamp 1698175906
transform 1 0 9800 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698175906
transform 1 0 10304 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 10416 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_222
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_230
timestamp 1698175906
transform 1 0 13552 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_234
timestamp 1698175906
transform 1 0 13776 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_236
timestamp 1698175906
transform 1 0 13888 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_257
timestamp 1698175906
transform 1 0 15064 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_289
timestamp 1698175906
transform 1 0 16856 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_305
timestamp 1698175906
transform 1 0 17752 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_313
timestamp 1698175906
transform 1 0 18200 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 2240 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 4032 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 4480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_88
timestamp 1698175906
transform 1 0 5600 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_96
timestamp 1698175906
transform 1 0 6048 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_100
timestamp 1698175906
transform 1 0 6272 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698175906
transform 1 0 8400 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_193
timestamp 1698175906
transform 1 0 11480 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_197
timestamp 1698175906
transform 1 0 11704 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698175906
transform 1 0 12264 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_228
timestamp 1698175906
transform 1 0 13440 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_236
timestamp 1698175906
transform 1 0 13888 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_272
timestamp 1698175906
transform 1 0 15904 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698175906
transform 1 0 16128 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 2240 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 2464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_69
timestamp 1698175906
transform 1 0 4536 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_73
timestamp 1698175906
transform 1 0 4760 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_75
timestamp 1698175906
transform 1 0 4872 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_112
timestamp 1698175906
transform 1 0 6944 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_116
timestamp 1698175906
transform 1 0 7168 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_124
timestamp 1698175906
transform 1 0 7616 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_128
timestamp 1698175906
transform 1 0 7840 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_134
timestamp 1698175906
transform 1 0 8176 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_140
timestamp 1698175906
transform 1 0 8512 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_147
timestamp 1698175906
transform 1 0 8904 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_155
timestamp 1698175906
transform 1 0 9352 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_188
timestamp 1698175906
transform 1 0 11200 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_192
timestamp 1698175906
transform 1 0 11424 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_222
timestamp 1698175906
transform 1 0 13104 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_226
timestamp 1698175906
transform 1 0 13328 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698175906
transform 1 0 14224 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 14336 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_88
timestamp 1698175906
transform 1 0 5600 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_92
timestamp 1698175906
transform 1 0 5824 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_94
timestamp 1698175906
transform 1 0 5936 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_124
timestamp 1698175906
transform 1 0 7616 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_128
timestamp 1698175906
transform 1 0 7840 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698175906
transform 1 0 8288 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_158
timestamp 1698175906
transform 1 0 9520 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698175906
transform 1 0 12208 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_220
timestamp 1698175906
transform 1 0 12992 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_224
timestamp 1698175906
transform 1 0 13216 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_254
timestamp 1698175906
transform 1 0 14896 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_258
timestamp 1698175906
transform 1 0 15120 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_274
timestamp 1698175906
transform 1 0 16016 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698175906
transform 1 0 16240 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_136
timestamp 1698175906
transform 1 0 8288 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_140
timestamp 1698175906
transform 1 0 8512 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_148
timestamp 1698175906
transform 1 0 8960 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_159
timestamp 1698175906
transform 1 0 9576 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_167
timestamp 1698175906
transform 1 0 10024 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_169
timestamp 1698175906
transform 1 0 10136 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_185
timestamp 1698175906
transform 1 0 11032 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_187
timestamp 1698175906
transform 1 0 11144 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_190
timestamp 1698175906
transform 1 0 11312 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_222
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_226
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_233
timestamp 1698175906
transform 1 0 13720 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 14336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_252
timestamp 1698175906
transform 1 0 14784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_284
timestamp 1698175906
transform 1 0 16576 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_300
timestamp 1698175906
transform 1 0 17472 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_308
timestamp 1698175906
transform 1 0 17920 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_312
timestamp 1698175906
transform 1 0 18144 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698175906
transform 1 0 18256 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 2240 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 4032 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 4480 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_104
timestamp 1698175906
transform 1 0 6496 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_137
timestamp 1698175906
transform 1 0 8344 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 8456 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_144
timestamp 1698175906
transform 1 0 8736 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_159
timestamp 1698175906
transform 1 0 9576 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_194
timestamp 1698175906
transform 1 0 11536 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_201
timestamp 1698175906
transform 1 0 11928 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 12376 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_212
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_216
timestamp 1698175906
transform 1 0 12768 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_218
timestamp 1698175906
transform 1 0 12880 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_248
timestamp 1698175906
transform 1 0 14560 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_252
timestamp 1698175906
transform 1 0 14784 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_268
timestamp 1698175906
transform 1 0 15680 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 16128 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_123
timestamp 1698175906
transform 1 0 7560 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_127
timestamp 1698175906
transform 1 0 7784 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_163
timestamp 1698175906
transform 1 0 9800 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_167
timestamp 1698175906
transform 1 0 10024 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_179
timestamp 1698175906
transform 1 0 10696 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_209
timestamp 1698175906
transform 1 0 12376 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_213
timestamp 1698175906
transform 1 0 12600 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 18648 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_150
timestamp 1698175906
transform 1 0 9072 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_152
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_159
timestamp 1698175906
transform 1 0 9576 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_175
timestamp 1698175906
transform 1 0 10472 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_183
timestamp 1698175906
transform 1 0 10920 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_185
timestamp 1698175906
transform 1 0 11032 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_196
timestamp 1698175906
transform 1 0 11648 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_204
timestamp 1698175906
transform 1 0 12096 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698175906
transform 1 0 12320 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_123
timestamp 1698175906
transform 1 0 7560 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_131
timestamp 1698175906
transform 1 0 8008 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_159
timestamp 1698175906
transform 1 0 9576 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_158
timestamp 1698175906
transform 1 0 9520 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_162
timestamp 1698175906
transform 1 0 9744 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_189
timestamp 1698175906
transform 1 0 11256 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_205
timestamp 1698175906
transform 1 0 12152 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 14000 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 15792 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 16240 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18760 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform -1 0 2240 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform -1 0 2240 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 8120 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 2240 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 8736 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18760 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform -1 0 2240 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 9800 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 18760 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 18760 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform -1 0 2240 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 2240 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 2240 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 2240 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 18760 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 18760 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698175906
transform -1 0 12096 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13440 400 13496 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 20600 7728 21000 7784 0 FreeSans 224 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 0 8400 400 8456 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 0 11424 400 11480 0 FreeSans 224 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 0 12768 400 12824 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 8064 20600 8120 21000 0 FreeSans 224 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 0 9744 400 9800 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 9408 20600 9464 21000 0 FreeSans 224 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 20600 8064 21000 8120 0 FreeSans 224 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 0 10080 400 10136 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 9744 20600 9800 21000 0 FreeSans 224 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 20600 10080 21000 10136 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 0 8064 400 8120 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 0 9408 400 9464 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 20600 10752 21000 10808 0 FreeSans 224 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 11760 400 11816 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 10752 400 10808 0 FreeSans 224 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 11424 20600 11480 21000 0 FreeSans 224 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 20600 8400 21000 8456 0 FreeSans 224 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 12096 20600 12152 21000 0 FreeSans 224 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 20600 9072 21000 9128 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 12096 0 12152 400 0 FreeSans 224 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 14644 8708 14644 8708 0 _000_
rlabel metal2 11228 13692 11228 13692 0 _001_
rlabel metal2 13468 12908 13468 12908 0 _002_
rlabel metal2 13020 7840 13020 7840 0 _003_
rlabel metal2 10360 12852 10360 12852 0 _004_
rlabel metal2 13776 12404 13776 12404 0 _005_
rlabel metal2 14000 10276 14000 10276 0 _006_
rlabel metal2 14224 8148 14224 8148 0 _007_
rlabel metal2 14364 9520 14364 9520 0 _008_
rlabel metal3 14476 11620 14476 11620 0 _009_
rlabel metal2 6440 11676 6440 11676 0 _010_
rlabel metal2 5908 10612 5908 10612 0 _011_
rlabel metal2 8848 13468 8848 13468 0 _012_
rlabel metal2 7000 7700 7000 7700 0 _013_
rlabel metal2 5964 9352 5964 9352 0 _014_
rlabel metal2 7028 8260 7028 8260 0 _015_
rlabel metal2 8064 11060 8064 11060 0 _016_
rlabel metal2 7140 12432 7140 12432 0 _017_
rlabel metal2 8036 12628 8036 12628 0 _018_
rlabel metal2 10108 11452 10108 11452 0 _019_
rlabel metal2 5908 9772 5908 9772 0 _020_
rlabel metal2 12068 11788 12068 11788 0 _021_
rlabel metal2 9772 10164 9772 10164 0 _022_
rlabel metal2 7644 7168 7644 7168 0 _023_
rlabel metal2 7980 10752 7980 10752 0 _024_
rlabel metal2 12404 8204 12404 8204 0 _025_
rlabel metal2 11480 7308 11480 7308 0 _026_
rlabel metal2 13524 9828 13524 9828 0 _027_
rlabel metal2 15092 8904 15092 8904 0 _028_
rlabel metal2 13692 9184 13692 9184 0 _029_
rlabel metal3 12684 9212 12684 9212 0 _030_
rlabel metal2 13692 10234 13692 10234 0 _031_
rlabel metal2 11088 13972 11088 13972 0 _032_
rlabel metal2 11648 13916 11648 13916 0 _033_
rlabel metal2 11620 13748 11620 13748 0 _034_
rlabel metal2 13580 11872 13580 11872 0 _035_
rlabel metal2 13636 12768 13636 12768 0 _036_
rlabel metal2 12852 8680 12852 8680 0 _037_
rlabel metal2 12908 10920 12908 10920 0 _038_
rlabel metal2 9380 12376 9380 12376 0 _039_
rlabel metal2 10472 13804 10472 13804 0 _040_
rlabel metal2 14056 10668 14056 10668 0 _041_
rlabel metal3 14364 12684 14364 12684 0 _042_
rlabel metal2 13720 10500 13720 10500 0 _043_
rlabel metal2 13076 10780 13076 10780 0 _044_
rlabel metal2 12516 10024 12516 10024 0 _045_
rlabel metal2 13860 10248 13860 10248 0 _046_
rlabel metal2 13804 9268 13804 9268 0 _047_
rlabel metal3 14392 7980 14392 7980 0 _048_
rlabel metal2 14308 9744 14308 9744 0 _049_
rlabel metal2 13748 9604 13748 9604 0 _050_
rlabel metal2 14532 10836 14532 10836 0 _051_
rlabel metal2 14756 11088 14756 11088 0 _052_
rlabel metal2 14980 11424 14980 11424 0 _053_
rlabel metal2 6412 11424 6412 11424 0 _054_
rlabel metal2 6692 11704 6692 11704 0 _055_
rlabel metal2 6916 10808 6916 10808 0 _056_
rlabel metal2 5852 10584 5852 10584 0 _057_
rlabel metal2 9324 13244 9324 13244 0 _058_
rlabel metal2 8764 9772 8764 9772 0 _059_
rlabel metal2 8820 11676 8820 11676 0 _060_
rlabel metal3 8540 8764 8540 8764 0 _061_
rlabel metal2 7308 8372 7308 8372 0 _062_
rlabel metal2 7924 9016 7924 9016 0 _063_
rlabel metal2 7756 8568 7756 8568 0 _064_
rlabel metal2 7756 7980 7756 7980 0 _065_
rlabel metal2 7196 12656 7196 12656 0 _066_
rlabel metal2 6580 9408 6580 9408 0 _067_
rlabel metal2 7364 8428 7364 8428 0 _068_
rlabel metal2 8120 11172 8120 11172 0 _069_
rlabel metal2 8260 11480 8260 11480 0 _070_
rlabel metal3 7476 12740 7476 12740 0 _071_
rlabel metal2 7476 12628 7476 12628 0 _072_
rlabel metal2 8148 13076 8148 13076 0 _073_
rlabel metal2 8260 12768 8260 12768 0 _074_
rlabel metal2 9436 8568 9436 8568 0 _075_
rlabel metal2 6524 11228 6524 11228 0 _076_
rlabel metal3 10752 9212 10752 9212 0 _077_
rlabel metal2 10780 9324 10780 9324 0 _078_
rlabel metal2 12880 9604 12880 9604 0 _079_
rlabel metal2 12516 11200 12516 11200 0 _080_
rlabel metal2 8988 9632 8988 9632 0 _081_
rlabel metal2 10220 11648 10220 11648 0 _082_
rlabel metal2 9240 11564 9240 11564 0 _083_
rlabel metal2 10052 11312 10052 11312 0 _084_
rlabel metal2 10108 8596 10108 8596 0 _085_
rlabel metal2 10948 8932 10948 8932 0 _086_
rlabel metal2 11592 7532 11592 7532 0 _087_
rlabel metal2 10948 9436 10948 9436 0 _088_
rlabel metal2 10752 11172 10752 11172 0 _089_
rlabel metal2 11676 10388 11676 10388 0 _090_
rlabel metal3 11788 11620 11788 11620 0 _091_
rlabel metal2 10276 11480 10276 11480 0 _092_
rlabel metal2 12292 9464 12292 9464 0 _093_
rlabel metal2 10332 10164 10332 10164 0 _094_
rlabel metal2 8904 11564 8904 11564 0 _095_
rlabel metal3 9324 11620 9324 11620 0 _096_
rlabel metal2 9716 8176 9716 8176 0 _097_
rlabel metal2 7196 9800 7196 9800 0 _098_
rlabel metal2 10892 9072 10892 9072 0 _099_
rlabel metal2 6860 10024 6860 10024 0 _100_
rlabel metal2 6972 11900 6972 11900 0 _101_
rlabel metal3 6216 9940 6216 9940 0 _102_
rlabel metal2 12180 11984 12180 11984 0 _103_
rlabel metal2 14588 10192 14588 10192 0 _104_
rlabel metal2 9324 9072 9324 9072 0 _105_
rlabel metal2 8820 10976 8820 10976 0 _106_
rlabel metal3 9856 8764 9856 8764 0 _107_
rlabel metal2 11788 8624 11788 8624 0 _108_
rlabel metal2 11676 8932 11676 8932 0 _109_
rlabel metal2 11788 7728 11788 7728 0 _110_
rlabel metal2 14700 7812 14700 7812 0 _111_
rlabel metal3 1239 13468 1239 13468 0 clk
rlabel metal2 12600 10332 12600 10332 0 clknet_0_clk
rlabel metal2 8316 13496 8316 13496 0 clknet_1_0__leaf_clk
rlabel metal3 11704 13524 11704 13524 0 clknet_1_1__leaf_clk
rlabel metal2 10248 7644 10248 7644 0 dut8.count\[0\]
rlabel metal3 9016 7588 9016 7588 0 dut8.count\[1\]
rlabel metal2 9044 10500 9044 10500 0 dut8.count\[2\]
rlabel metal2 11340 8484 11340 8484 0 dut8.count\[3\]
rlabel metal3 15554 7924 15554 7924 0 net1
rlabel metal2 9716 13804 9716 13804 0 net10
rlabel metal2 15484 9800 15484 9800 0 net11
rlabel metal2 15820 11368 15820 11368 0 net12
rlabel metal2 5936 7588 5936 7588 0 net13
rlabel metal2 2156 9380 2156 9380 0 net14
rlabel metal2 18844 10948 18844 10948 0 net15
rlabel metal3 3178 11956 3178 11956 0 net16
rlabel metal2 2156 10948 2156 10948 0 net17
rlabel metal2 14644 12908 14644 12908 0 net18
rlabel metal3 11900 14028 11900 14028 0 net19
rlabel metal2 5964 8596 5964 8596 0 net2
rlabel metal2 14028 7588 14028 7588 0 net20
rlabel metal2 14196 12880 14196 12880 0 net21
rlabel metal3 12460 13580 12460 13580 0 net22
rlabel metal2 15540 8904 15540 8904 0 net23
rlabel metal2 12292 2982 12292 2982 0 net24
rlabel metal3 15960 12012 15960 12012 0 net25
rlabel metal3 11592 12460 11592 12460 0 net26
rlabel metal2 2156 11536 2156 11536 0 net3
rlabel metal2 6076 12712 6076 12712 0 net4
rlabel metal2 8148 13524 8148 13524 0 net5
rlabel metal3 3178 9996 3178 9996 0 net6
rlabel metal3 9156 19012 9156 19012 0 net7
rlabel metal2 15036 8204 15036 8204 0 net8
rlabel metal2 2100 10136 2100 10136 0 net9
rlabel metal2 20020 7924 20020 7924 0 segm[0]
rlabel metal3 679 8428 679 8428 0 segm[10]
rlabel metal3 679 11452 679 11452 0 segm[11]
rlabel metal3 679 12796 679 12796 0 segm[12]
rlabel metal2 8092 19481 8092 19481 0 segm[13]
rlabel metal3 679 9772 679 9772 0 segm[1]
rlabel metal2 9436 19845 9436 19845 0 segm[2]
rlabel metal2 19964 8232 19964 8232 0 segm[3]
rlabel metal3 679 10108 679 10108 0 segm[4]
rlabel metal2 9772 19677 9772 19677 0 segm[5]
rlabel metal2 20020 10276 20020 10276 0 segm[6]
rlabel metal3 20321 11452 20321 11452 0 segm[7]
rlabel metal3 679 8092 679 8092 0 segm[8]
rlabel metal3 679 9436 679 9436 0 segm[9]
rlabel metal2 20020 11004 20020 11004 0 sel[0]
rlabel metal3 679 11788 679 11788 0 sel[10]
rlabel metal3 679 10780 679 10780 0 sel[11]
rlabel metal2 20020 12908 20020 12908 0 sel[1]
rlabel metal2 11452 19873 11452 19873 0 sel[2]
rlabel metal2 20020 8652 20020 8652 0 sel[3]
rlabel metal2 20020 13356 20020 13356 0 sel[4]
rlabel metal2 12124 19677 12124 19677 0 sel[5]
rlabel metal3 20321 9100 20321 9100 0 sel[6]
rlabel metal2 12124 1099 12124 1099 0 sel[7]
rlabel metal2 20020 11900 20020 11900 0 sel[8]
rlabel metal2 11116 19845 11116 19845 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
