magic
tech gf180mcuD
magscale 1 10
timestamp 1699643108
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 18162 38110 18174 38162
rect 18226 38110 18238 38162
rect 22194 38110 22206 38162
rect 22258 38110 22270 38162
rect 19730 37998 19742 38050
rect 19794 37998 19806 38050
rect 23650 37998 23662 38050
rect 23714 37998 23726 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 20750 37490 20802 37502
rect 20750 37426 20802 37438
rect 19730 37214 19742 37266
rect 19794 37214 19806 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 1934 27186 1986 27198
rect 1934 27122 1986 27134
rect 4274 27022 4286 27074
rect 4338 27022 4350 27074
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 26238 26402 26290 26414
rect 26238 26338 26290 26350
rect 26014 26290 26066 26302
rect 4274 26238 4286 26290
rect 4338 26238 4350 26290
rect 17378 26238 17390 26290
rect 17442 26238 17454 26290
rect 21186 26238 21198 26290
rect 21250 26238 21262 26290
rect 26014 26226 26066 26238
rect 26350 26290 26402 26302
rect 37650 26238 37662 26290
rect 37714 26238 37726 26290
rect 26350 26226 26402 26238
rect 16942 26178 16994 26190
rect 24670 26178 24722 26190
rect 18162 26126 18174 26178
rect 18226 26126 18238 26178
rect 20290 26126 20302 26178
rect 20354 26126 20366 26178
rect 21970 26126 21982 26178
rect 22034 26126 22046 26178
rect 24098 26126 24110 26178
rect 24162 26126 24174 26178
rect 39890 26126 39902 26178
rect 39954 26126 39966 26178
rect 16942 26114 16994 26126
rect 24670 26114 24722 26126
rect 1934 26066 1986 26078
rect 1934 26002 1986 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 19966 25730 20018 25742
rect 19966 25666 20018 25678
rect 19070 25618 19122 25630
rect 2034 25566 2046 25618
rect 2098 25566 2110 25618
rect 18610 25566 18622 25618
rect 18674 25566 18686 25618
rect 19070 25554 19122 25566
rect 21982 25618 22034 25630
rect 40014 25618 40066 25630
rect 27346 25566 27358 25618
rect 27410 25566 27422 25618
rect 21982 25554 22034 25566
rect 40014 25554 40066 25566
rect 19630 25506 19682 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 14242 25454 14254 25506
rect 14306 25454 14318 25506
rect 14914 25454 14926 25506
rect 14978 25454 14990 25506
rect 15698 25454 15710 25506
rect 15762 25454 15774 25506
rect 19630 25442 19682 25454
rect 22542 25506 22594 25518
rect 22542 25442 22594 25454
rect 23214 25506 23266 25518
rect 23214 25442 23266 25454
rect 23550 25506 23602 25518
rect 24546 25454 24558 25506
rect 24610 25454 24622 25506
rect 37874 25454 37886 25506
rect 37938 25454 37950 25506
rect 23550 25442 23602 25454
rect 19854 25394 19906 25406
rect 14018 25342 14030 25394
rect 14082 25342 14094 25394
rect 14690 25342 14702 25394
rect 14754 25342 14766 25394
rect 16482 25342 16494 25394
rect 16546 25342 16558 25394
rect 19854 25330 19906 25342
rect 19966 25394 20018 25406
rect 19966 25330 20018 25342
rect 22990 25394 23042 25406
rect 22990 25330 23042 25342
rect 23438 25394 23490 25406
rect 25218 25342 25230 25394
rect 25282 25342 25294 25394
rect 23438 25330 23490 25342
rect 18958 25282 19010 25294
rect 18958 25218 19010 25230
rect 19182 25282 19234 25294
rect 19182 25218 19234 25230
rect 21870 25282 21922 25294
rect 21870 25218 21922 25230
rect 22094 25282 22146 25294
rect 22094 25218 22146 25230
rect 22654 25282 22706 25294
rect 22654 25218 22706 25230
rect 22878 25282 22930 25294
rect 22878 25218 22930 25230
rect 27806 25282 27858 25294
rect 27806 25218 27858 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 14702 24946 14754 24958
rect 14702 24882 14754 24894
rect 14926 24946 14978 24958
rect 14926 24882 14978 24894
rect 17726 24946 17778 24958
rect 17726 24882 17778 24894
rect 18622 24946 18674 24958
rect 18622 24882 18674 24894
rect 19182 24946 19234 24958
rect 23314 24894 23326 24946
rect 23378 24894 23390 24946
rect 19182 24882 19234 24894
rect 17614 24834 17666 24846
rect 17614 24770 17666 24782
rect 18398 24834 18450 24846
rect 18398 24770 18450 24782
rect 18734 24834 18786 24846
rect 18734 24770 18786 24782
rect 15038 24722 15090 24734
rect 4274 24670 4286 24722
rect 4338 24670 4350 24722
rect 11554 24670 11566 24722
rect 11618 24670 11630 24722
rect 15038 24658 15090 24670
rect 17838 24722 17890 24734
rect 17838 24658 17890 24670
rect 18286 24722 18338 24734
rect 22990 24722 23042 24734
rect 19842 24670 19854 24722
rect 19906 24670 19918 24722
rect 25218 24670 25230 24722
rect 25282 24670 25294 24722
rect 37650 24670 37662 24722
rect 37714 24670 37726 24722
rect 18286 24658 18338 24670
rect 22990 24658 23042 24670
rect 15486 24610 15538 24622
rect 23774 24610 23826 24622
rect 28590 24610 28642 24622
rect 12338 24558 12350 24610
rect 12402 24558 12414 24610
rect 14466 24558 14478 24610
rect 14530 24558 14542 24610
rect 20514 24558 20526 24610
rect 20578 24558 20590 24610
rect 22642 24558 22654 24610
rect 22706 24558 22718 24610
rect 26002 24558 26014 24610
rect 26066 24558 26078 24610
rect 28130 24558 28142 24610
rect 28194 24558 28206 24610
rect 15486 24546 15538 24558
rect 23774 24546 23826 24558
rect 28590 24546 28642 24558
rect 1934 24498 1986 24510
rect 1934 24434 1986 24446
rect 40014 24498 40066 24510
rect 40014 24434 40066 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 21422 24050 21474 24062
rect 21422 23986 21474 23998
rect 25342 24050 25394 24062
rect 25342 23986 25394 23998
rect 12574 23938 12626 23950
rect 12574 23874 12626 23886
rect 13918 23938 13970 23950
rect 13918 23874 13970 23886
rect 21982 23938 22034 23950
rect 21982 23874 22034 23886
rect 25902 23938 25954 23950
rect 25902 23874 25954 23886
rect 26238 23938 26290 23950
rect 27346 23886 27358 23938
rect 27410 23886 27422 23938
rect 26238 23874 26290 23886
rect 12910 23826 12962 23838
rect 12910 23762 12962 23774
rect 14142 23826 14194 23838
rect 14142 23762 14194 23774
rect 14366 23826 14418 23838
rect 14366 23762 14418 23774
rect 14478 23826 14530 23838
rect 25230 23826 25282 23838
rect 17378 23774 17390 23826
rect 17442 23774 17454 23826
rect 27570 23774 27582 23826
rect 27634 23774 27646 23826
rect 14478 23762 14530 23774
rect 25230 23762 25282 23774
rect 12798 23714 12850 23726
rect 12798 23650 12850 23662
rect 13582 23714 13634 23726
rect 13582 23650 13634 23662
rect 13806 23714 13858 23726
rect 13806 23650 13858 23662
rect 17726 23714 17778 23726
rect 17726 23650 17778 23662
rect 21310 23714 21362 23726
rect 21310 23650 21362 23662
rect 21534 23714 21586 23726
rect 21534 23650 21586 23662
rect 25454 23714 25506 23726
rect 25454 23650 25506 23662
rect 26126 23714 26178 23726
rect 26126 23650 26178 23662
rect 26350 23714 26402 23726
rect 26350 23650 26402 23662
rect 26574 23714 26626 23726
rect 26574 23650 26626 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 26350 23378 26402 23390
rect 26350 23314 26402 23326
rect 26574 23378 26626 23390
rect 26574 23314 26626 23326
rect 13794 23214 13806 23266
rect 13858 23214 13870 23266
rect 15038 23154 15090 23166
rect 26238 23154 26290 23166
rect 4274 23102 4286 23154
rect 4338 23102 4350 23154
rect 14466 23102 14478 23154
rect 14530 23102 14542 23154
rect 20290 23102 20302 23154
rect 20354 23102 20366 23154
rect 15038 23090 15090 23102
rect 26238 23090 26290 23102
rect 11678 23042 11730 23054
rect 20750 23042 20802 23054
rect 17378 22990 17390 23042
rect 17442 22990 17454 23042
rect 19506 22990 19518 23042
rect 19570 22990 19582 23042
rect 11678 22978 11730 22990
rect 20750 22978 20802 22990
rect 1934 22930 1986 22942
rect 1934 22866 1986 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 17950 22482 18002 22494
rect 40014 22482 40066 22494
rect 24210 22430 24222 22482
rect 24274 22430 24286 22482
rect 17950 22418 18002 22430
rect 40014 22418 40066 22430
rect 16718 22370 16770 22382
rect 16718 22306 16770 22318
rect 17166 22370 17218 22382
rect 18286 22370 18338 22382
rect 17714 22318 17726 22370
rect 17778 22318 17790 22370
rect 17166 22306 17218 22318
rect 18286 22306 18338 22318
rect 18734 22370 18786 22382
rect 21298 22318 21310 22370
rect 21362 22318 21374 22370
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 18734 22306 18786 22318
rect 17054 22258 17106 22270
rect 17054 22194 17106 22206
rect 18062 22258 18114 22270
rect 18062 22194 18114 22206
rect 18846 22258 18898 22270
rect 22082 22206 22094 22258
rect 22146 22206 22158 22258
rect 18846 22194 18898 22206
rect 14366 22146 14418 22158
rect 14366 22082 14418 22094
rect 16830 22146 16882 22158
rect 16830 22082 16882 22094
rect 18958 22146 19010 22158
rect 18958 22082 19010 22094
rect 24670 22146 24722 22158
rect 24670 22082 24722 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 16494 21810 16546 21822
rect 22878 21810 22930 21822
rect 16818 21758 16830 21810
rect 16882 21758 16894 21810
rect 16494 21746 16546 21758
rect 22878 21746 22930 21758
rect 15150 21698 15202 21710
rect 19518 21698 19570 21710
rect 12002 21646 12014 21698
rect 12066 21646 12078 21698
rect 17826 21646 17838 21698
rect 17890 21646 17902 21698
rect 18162 21646 18174 21698
rect 18226 21646 18238 21698
rect 19058 21646 19070 21698
rect 19122 21646 19134 21698
rect 15150 21634 15202 21646
rect 19518 21634 19570 21646
rect 19630 21698 19682 21710
rect 19630 21634 19682 21646
rect 22094 21698 22146 21710
rect 22094 21634 22146 21646
rect 22990 21698 23042 21710
rect 22990 21634 23042 21646
rect 23326 21698 23378 21710
rect 23326 21634 23378 21646
rect 23438 21698 23490 21710
rect 23438 21634 23490 21646
rect 27134 21698 27186 21710
rect 27134 21634 27186 21646
rect 27246 21698 27298 21710
rect 27246 21634 27298 21646
rect 27582 21698 27634 21710
rect 27582 21634 27634 21646
rect 27694 21698 27746 21710
rect 27694 21634 27746 21646
rect 14702 21586 14754 21598
rect 11330 21534 11342 21586
rect 11394 21534 11406 21586
rect 14354 21534 14366 21586
rect 14418 21583 14430 21586
rect 14578 21583 14590 21586
rect 14418 21537 14590 21583
rect 14418 21534 14430 21537
rect 14578 21534 14590 21537
rect 14642 21534 14654 21586
rect 14702 21522 14754 21534
rect 15262 21586 15314 21598
rect 15262 21522 15314 21534
rect 16158 21586 16210 21598
rect 21646 21586 21698 21598
rect 17938 21534 17950 21586
rect 18002 21534 18014 21586
rect 18834 21534 18846 21586
rect 18898 21534 18910 21586
rect 16158 21522 16210 21534
rect 21646 21522 21698 21534
rect 22318 21586 22370 21598
rect 22318 21522 22370 21534
rect 22430 21586 22482 21598
rect 22430 21522 22482 21534
rect 22654 21586 22706 21598
rect 22654 21522 22706 21534
rect 26126 21586 26178 21598
rect 26126 21522 26178 21534
rect 26350 21586 26402 21598
rect 26350 21522 26402 21534
rect 26798 21586 26850 21598
rect 26798 21522 26850 21534
rect 26910 21586 26962 21598
rect 26910 21522 26962 21534
rect 27918 21586 27970 21598
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 27918 21522 27970 21534
rect 15598 21474 15650 21486
rect 14130 21422 14142 21474
rect 14194 21422 14206 21474
rect 15598 21410 15650 21422
rect 21870 21474 21922 21486
rect 21870 21410 21922 21422
rect 25230 21474 25282 21486
rect 25230 21410 25282 21422
rect 26574 21474 26626 21486
rect 26574 21410 26626 21422
rect 40014 21474 40066 21486
rect 40014 21410 40066 21422
rect 14814 21362 14866 21374
rect 14814 21298 14866 21310
rect 19518 21362 19570 21374
rect 19518 21298 19570 21310
rect 23438 21362 23490 21374
rect 23438 21298 23490 21310
rect 25454 21362 25506 21374
rect 25454 21298 25506 21310
rect 25790 21362 25842 21374
rect 25790 21298 25842 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 20862 21026 20914 21038
rect 20862 20962 20914 20974
rect 40014 20914 40066 20926
rect 40014 20850 40066 20862
rect 14142 20802 14194 20814
rect 14142 20738 14194 20750
rect 14366 20802 14418 20814
rect 20190 20802 20242 20814
rect 19954 20750 19966 20802
rect 20018 20750 20030 20802
rect 20514 20750 20526 20802
rect 20578 20750 20590 20802
rect 21858 20750 21870 20802
rect 21922 20750 21934 20802
rect 37650 20750 37662 20802
rect 37714 20750 37726 20802
rect 14366 20738 14418 20750
rect 20190 20738 20242 20750
rect 13918 20690 13970 20702
rect 20750 20690 20802 20702
rect 15362 20638 15374 20690
rect 15426 20638 15438 20690
rect 25442 20638 25454 20690
rect 25506 20638 25518 20690
rect 13918 20626 13970 20638
rect 20750 20626 20802 20638
rect 14254 20578 14306 20590
rect 14254 20514 14306 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 14478 20130 14530 20142
rect 18174 20130 18226 20142
rect 11890 20078 11902 20130
rect 11954 20078 11966 20130
rect 16818 20078 16830 20130
rect 16882 20078 16894 20130
rect 21858 20078 21870 20130
rect 21922 20078 21934 20130
rect 26114 20078 26126 20130
rect 26178 20078 26190 20130
rect 14478 20066 14530 20078
rect 18174 20066 18226 20078
rect 17950 20018 18002 20030
rect 11218 19966 11230 20018
rect 11282 19966 11294 20018
rect 15474 19966 15486 20018
rect 15538 19966 15550 20018
rect 15698 19966 15710 20018
rect 15762 19966 15774 20018
rect 16594 19966 16606 20018
rect 16658 19966 16670 20018
rect 17602 19966 17614 20018
rect 17666 19966 17678 20018
rect 18498 19966 18510 20018
rect 18562 19966 18574 20018
rect 25442 19966 25454 20018
rect 25506 19966 25518 20018
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 17950 19954 18002 19966
rect 15934 19906 15986 19918
rect 28702 19906 28754 19918
rect 14018 19854 14030 19906
rect 14082 19854 14094 19906
rect 28242 19854 28254 19906
rect 28306 19854 28318 19906
rect 15934 19842 15986 19854
rect 28702 19842 28754 19854
rect 40014 19906 40066 19918
rect 40014 19842 40066 19854
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 14926 19458 14978 19470
rect 14926 19394 14978 19406
rect 15374 19458 15426 19470
rect 15374 19394 15426 19406
rect 17154 19294 17166 19346
rect 17218 19294 17230 19346
rect 24210 19294 24222 19346
rect 24274 19294 24286 19346
rect 28354 19294 28366 19346
rect 28418 19294 28430 19346
rect 15934 19234 15986 19246
rect 24670 19234 24722 19246
rect 16930 19182 16942 19234
rect 16994 19182 17006 19234
rect 17938 19182 17950 19234
rect 18002 19182 18014 19234
rect 19954 19182 19966 19234
rect 20018 19182 20030 19234
rect 21410 19182 21422 19234
rect 21474 19182 21486 19234
rect 25442 19182 25454 19234
rect 25506 19182 25518 19234
rect 15934 19170 15986 19182
rect 24670 19170 24722 19182
rect 14702 19122 14754 19134
rect 14702 19058 14754 19070
rect 15262 19122 15314 19134
rect 15262 19058 15314 19070
rect 17502 19122 17554 19134
rect 18162 19070 18174 19122
rect 18226 19070 18238 19122
rect 18498 19070 18510 19122
rect 18562 19070 18574 19122
rect 19618 19070 19630 19122
rect 19682 19070 19694 19122
rect 20178 19070 20190 19122
rect 20242 19070 20254 19122
rect 20626 19070 20638 19122
rect 20690 19070 20702 19122
rect 22082 19070 22094 19122
rect 22146 19070 22158 19122
rect 26226 19070 26238 19122
rect 26290 19070 26302 19122
rect 17502 19058 17554 19070
rect 14814 19010 14866 19022
rect 14814 18946 14866 18958
rect 15374 19010 15426 19022
rect 19294 19010 19346 19022
rect 16258 18958 16270 19010
rect 16322 18958 16334 19010
rect 18610 18958 18622 19010
rect 18674 18958 18686 19010
rect 15374 18946 15426 18958
rect 19294 18946 19346 18958
rect 29262 19010 29314 19022
rect 29262 18946 29314 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 14030 18674 14082 18686
rect 14030 18610 14082 18622
rect 20302 18674 20354 18686
rect 20302 18610 20354 18622
rect 20526 18674 20578 18686
rect 20526 18610 20578 18622
rect 21870 18674 21922 18686
rect 21870 18610 21922 18622
rect 26126 18674 26178 18686
rect 27122 18622 27134 18674
rect 27186 18622 27198 18674
rect 26126 18610 26178 18622
rect 16606 18562 16658 18574
rect 14354 18510 14366 18562
rect 14418 18510 14430 18562
rect 21298 18510 21310 18562
rect 21362 18510 21374 18562
rect 16606 18498 16658 18510
rect 17950 18450 18002 18462
rect 22542 18450 22594 18462
rect 14578 18398 14590 18450
rect 14642 18398 14654 18450
rect 15586 18398 15598 18450
rect 15650 18398 15662 18450
rect 15922 18398 15934 18450
rect 15986 18398 15998 18450
rect 18498 18398 18510 18450
rect 18562 18398 18574 18450
rect 18834 18398 18846 18450
rect 18898 18398 18910 18450
rect 19730 18398 19742 18450
rect 19794 18398 19806 18450
rect 20066 18398 20078 18450
rect 20130 18398 20142 18450
rect 20962 18398 20974 18450
rect 21026 18398 21038 18450
rect 17950 18386 18002 18398
rect 22542 18386 22594 18398
rect 22766 18450 22818 18462
rect 22766 18386 22818 18398
rect 23102 18450 23154 18462
rect 23102 18386 23154 18398
rect 23214 18450 23266 18462
rect 23214 18386 23266 18398
rect 25790 18450 25842 18462
rect 25790 18386 25842 18398
rect 26238 18450 26290 18462
rect 26238 18386 26290 18398
rect 26462 18450 26514 18462
rect 26462 18386 26514 18398
rect 26798 18450 26850 18462
rect 26798 18386 26850 18398
rect 20414 18338 20466 18350
rect 14914 18286 14926 18338
rect 14978 18286 14990 18338
rect 16482 18286 16494 18338
rect 16546 18286 16558 18338
rect 19170 18286 19182 18338
rect 19234 18286 19246 18338
rect 21410 18286 21422 18338
rect 21474 18286 21486 18338
rect 20414 18274 20466 18286
rect 16830 18226 16882 18238
rect 21982 18226 22034 18238
rect 18834 18174 18846 18226
rect 18898 18174 18910 18226
rect 16830 18162 16882 18174
rect 21982 18162 22034 18174
rect 22206 18226 22258 18238
rect 22206 18162 22258 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 14254 17890 14306 17902
rect 14254 17826 14306 17838
rect 14814 17890 14866 17902
rect 14814 17826 14866 17838
rect 15822 17890 15874 17902
rect 21422 17890 21474 17902
rect 17154 17838 17166 17890
rect 17218 17838 17230 17890
rect 15822 17826 15874 17838
rect 21422 17826 21474 17838
rect 21758 17890 21810 17902
rect 21758 17826 21810 17838
rect 1934 17778 1986 17790
rect 40014 17778 40066 17790
rect 15474 17726 15486 17778
rect 15538 17726 15550 17778
rect 1934 17714 1986 17726
rect 40014 17714 40066 17726
rect 15038 17666 15090 17678
rect 21982 17666 22034 17678
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 16482 17614 16494 17666
rect 16546 17614 16558 17666
rect 17154 17614 17166 17666
rect 17218 17614 17230 17666
rect 17602 17614 17614 17666
rect 17666 17614 17678 17666
rect 19506 17614 19518 17666
rect 19570 17614 19582 17666
rect 15038 17602 15090 17614
rect 21982 17602 22034 17614
rect 22430 17666 22482 17678
rect 22430 17602 22482 17614
rect 24782 17666 24834 17678
rect 24782 17602 24834 17614
rect 26014 17666 26066 17678
rect 26014 17602 26066 17614
rect 26574 17666 26626 17678
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 26574 17602 26626 17614
rect 14478 17554 14530 17566
rect 14478 17490 14530 17502
rect 14590 17554 14642 17566
rect 14590 17490 14642 17502
rect 15598 17554 15650 17566
rect 19294 17554 19346 17566
rect 16258 17502 16270 17554
rect 16322 17502 16334 17554
rect 15598 17490 15650 17502
rect 19294 17490 19346 17502
rect 19742 17554 19794 17566
rect 19742 17490 19794 17502
rect 22318 17554 22370 17566
rect 22318 17490 22370 17502
rect 25230 17554 25282 17566
rect 25230 17490 25282 17502
rect 25454 17554 25506 17566
rect 25454 17490 25506 17502
rect 25902 17554 25954 17566
rect 25902 17490 25954 17502
rect 26238 17554 26290 17566
rect 26238 17490 26290 17502
rect 19854 17442 19906 17454
rect 19854 17378 19906 17390
rect 25118 17442 25170 17454
rect 25118 17378 25170 17390
rect 25678 17442 25730 17454
rect 25678 17378 25730 17390
rect 26462 17442 26514 17454
rect 26462 17378 26514 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 14702 17106 14754 17118
rect 14702 17042 14754 17054
rect 19630 17106 19682 17118
rect 19630 17042 19682 17054
rect 19966 17106 20018 17118
rect 22082 17054 22094 17106
rect 22146 17054 22158 17106
rect 19966 17042 20018 17054
rect 15038 16994 15090 17006
rect 12786 16942 12798 16994
rect 12850 16942 12862 16994
rect 15038 16930 15090 16942
rect 15374 16994 15426 17006
rect 15374 16930 15426 16942
rect 15598 16994 15650 17006
rect 15598 16930 15650 16942
rect 15822 16994 15874 17006
rect 15822 16930 15874 16942
rect 19854 16994 19906 17006
rect 26002 16942 26014 16994
rect 26066 16942 26078 16994
rect 19854 16930 19906 16942
rect 14478 16882 14530 16894
rect 13570 16830 13582 16882
rect 13634 16830 13646 16882
rect 14478 16818 14530 16830
rect 14814 16882 14866 16894
rect 14814 16818 14866 16830
rect 19294 16882 19346 16894
rect 23998 16882 24050 16894
rect 21858 16830 21870 16882
rect 21922 16830 21934 16882
rect 19294 16818 19346 16830
rect 23998 16818 24050 16830
rect 24334 16882 24386 16894
rect 24334 16818 24386 16830
rect 24670 16882 24722 16894
rect 28590 16882 28642 16894
rect 25218 16830 25230 16882
rect 25282 16830 25294 16882
rect 37650 16830 37662 16882
rect 37714 16830 37726 16882
rect 24670 16818 24722 16830
rect 28590 16818 28642 16830
rect 14030 16770 14082 16782
rect 10658 16718 10670 16770
rect 10722 16718 10734 16770
rect 14030 16706 14082 16718
rect 15262 16770 15314 16782
rect 15262 16706 15314 16718
rect 24222 16770 24274 16782
rect 40014 16770 40066 16782
rect 28130 16718 28142 16770
rect 28194 16718 28206 16770
rect 24222 16706 24274 16718
rect 40014 16706 40066 16718
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 18386 16270 18398 16322
rect 18450 16270 18462 16322
rect 1934 16210 1986 16222
rect 1934 16146 1986 16158
rect 15710 16210 15762 16222
rect 24994 16158 25006 16210
rect 25058 16158 25070 16210
rect 27122 16158 27134 16210
rect 27186 16158 27198 16210
rect 15710 16146 15762 16158
rect 14142 16098 14194 16110
rect 4274 16046 4286 16098
rect 4338 16046 4350 16098
rect 14142 16034 14194 16046
rect 14702 16098 14754 16110
rect 14702 16034 14754 16046
rect 15598 16098 15650 16110
rect 15598 16034 15650 16046
rect 18734 16098 18786 16110
rect 18734 16034 18786 16046
rect 18958 16098 19010 16110
rect 18958 16034 19010 16046
rect 20078 16098 20130 16110
rect 20078 16034 20130 16046
rect 20302 16098 20354 16110
rect 20302 16034 20354 16046
rect 20750 16098 20802 16110
rect 27582 16098 27634 16110
rect 24210 16046 24222 16098
rect 24274 16046 24286 16098
rect 20750 16034 20802 16046
rect 27582 16034 27634 16046
rect 14366 15986 14418 15998
rect 14366 15922 14418 15934
rect 15934 15986 15986 15998
rect 15934 15922 15986 15934
rect 16158 15986 16210 15998
rect 16158 15922 16210 15934
rect 14590 15874 14642 15886
rect 14590 15810 14642 15822
rect 15150 15874 15202 15886
rect 15150 15810 15202 15822
rect 20190 15874 20242 15886
rect 20190 15810 20242 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 15710 15538 15762 15550
rect 15710 15474 15762 15486
rect 18398 15538 18450 15550
rect 18398 15474 18450 15486
rect 20302 15538 20354 15550
rect 20302 15474 20354 15486
rect 16158 15426 16210 15438
rect 16158 15362 16210 15374
rect 16382 15426 16434 15438
rect 19630 15426 19682 15438
rect 19394 15374 19406 15426
rect 19458 15374 19470 15426
rect 22978 15374 22990 15426
rect 23042 15374 23054 15426
rect 16382 15362 16434 15374
rect 19630 15362 19682 15374
rect 14702 15314 14754 15326
rect 18510 15314 18562 15326
rect 19966 15314 20018 15326
rect 24222 15314 24274 15326
rect 13906 15262 13918 15314
rect 13970 15262 13982 15314
rect 15474 15262 15486 15314
rect 15538 15262 15550 15314
rect 18274 15262 18286 15314
rect 18338 15262 18350 15314
rect 18834 15262 18846 15314
rect 18898 15262 18910 15314
rect 23650 15262 23662 15314
rect 23714 15262 23726 15314
rect 14702 15250 14754 15262
rect 18510 15250 18562 15262
rect 19966 15250 20018 15262
rect 24222 15250 24274 15262
rect 14254 15202 14306 15214
rect 19518 15202 19570 15214
rect 10994 15150 11006 15202
rect 11058 15150 11070 15202
rect 13122 15150 13134 15202
rect 13186 15150 13198 15202
rect 16034 15150 16046 15202
rect 16098 15150 16110 15202
rect 20850 15150 20862 15202
rect 20914 15150 20926 15202
rect 14254 15138 14306 15150
rect 19518 15138 19570 15150
rect 14366 15090 14418 15102
rect 14366 15026 14418 15038
rect 14590 15090 14642 15102
rect 19058 15038 19070 15090
rect 19122 15038 19134 15090
rect 14590 15026 14642 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 15262 14754 15314 14766
rect 15262 14690 15314 14702
rect 15374 14754 15426 14766
rect 15374 14690 15426 14702
rect 14242 14590 14254 14642
rect 14306 14590 14318 14642
rect 16594 14590 16606 14642
rect 16658 14590 16670 14642
rect 18722 14590 18734 14642
rect 18786 14590 18798 14642
rect 15038 14530 15090 14542
rect 15922 14478 15934 14530
rect 15986 14478 15998 14530
rect 21634 14478 21646 14530
rect 21698 14478 21710 14530
rect 22418 14478 22430 14530
rect 22482 14478 22494 14530
rect 15038 14466 15090 14478
rect 14366 14418 14418 14430
rect 14366 14354 14418 14366
rect 14590 14418 14642 14430
rect 14590 14354 14642 14366
rect 14926 14418 14978 14430
rect 14926 14354 14978 14366
rect 19182 14306 19234 14318
rect 21858 14254 21870 14306
rect 21922 14254 21934 14306
rect 22194 14254 22206 14306
rect 22258 14254 22270 14306
rect 19182 14242 19234 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 16718 13970 16770 13982
rect 16718 13906 16770 13918
rect 14130 13806 14142 13858
rect 14194 13806 14206 13858
rect 19618 13806 19630 13858
rect 19682 13806 19694 13858
rect 22206 13746 22258 13758
rect 13458 13694 13470 13746
rect 13522 13694 13534 13746
rect 18946 13694 18958 13746
rect 19010 13694 19022 13746
rect 22206 13682 22258 13694
rect 16258 13582 16270 13634
rect 16322 13582 16334 13634
rect 21746 13582 21758 13634
rect 21810 13582 21822 13634
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 40238 6018 40290 6030
rect 40238 5954 40290 5966
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 22318 5234 22370 5246
rect 22318 5170 22370 5182
rect 21298 5070 21310 5122
rect 21362 5070 21374 5122
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 21858 4286 21870 4338
rect 21922 4286 21934 4338
rect 22766 4114 22818 4126
rect 22766 4050 22818 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 16930 3502 16942 3554
rect 16994 3502 17006 3554
rect 21746 3502 21758 3554
rect 21810 3502 21822 3554
rect 18498 3390 18510 3442
rect 18562 3390 18574 3442
rect 15710 3330 15762 3342
rect 15710 3266 15762 3278
rect 22430 3330 22482 3342
rect 22430 3266 22482 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 25566 38222 25618 38274
rect 18174 38110 18226 38162
rect 22206 38110 22258 38162
rect 19742 37998 19794 38050
rect 23662 37998 23714 38050
rect 24558 37998 24610 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 20750 37438 20802 37490
rect 19742 37214 19794 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 1934 27134 1986 27186
rect 4286 27022 4338 27074
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 26238 26350 26290 26402
rect 4286 26238 4338 26290
rect 17390 26238 17442 26290
rect 21198 26238 21250 26290
rect 26014 26238 26066 26290
rect 26350 26238 26402 26290
rect 37662 26238 37714 26290
rect 16942 26126 16994 26178
rect 18174 26126 18226 26178
rect 20302 26126 20354 26178
rect 21982 26126 22034 26178
rect 24110 26126 24162 26178
rect 24670 26126 24722 26178
rect 39902 26126 39954 26178
rect 1934 26014 1986 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 19966 25678 20018 25730
rect 2046 25566 2098 25618
rect 18622 25566 18674 25618
rect 19070 25566 19122 25618
rect 21982 25566 22034 25618
rect 27358 25566 27410 25618
rect 40014 25566 40066 25618
rect 4286 25454 4338 25506
rect 14254 25454 14306 25506
rect 14926 25454 14978 25506
rect 15710 25454 15762 25506
rect 19630 25454 19682 25506
rect 22542 25454 22594 25506
rect 23214 25454 23266 25506
rect 23550 25454 23602 25506
rect 24558 25454 24610 25506
rect 37886 25454 37938 25506
rect 14030 25342 14082 25394
rect 14702 25342 14754 25394
rect 16494 25342 16546 25394
rect 19854 25342 19906 25394
rect 19966 25342 20018 25394
rect 22990 25342 23042 25394
rect 23438 25342 23490 25394
rect 25230 25342 25282 25394
rect 18958 25230 19010 25282
rect 19182 25230 19234 25282
rect 21870 25230 21922 25282
rect 22094 25230 22146 25282
rect 22654 25230 22706 25282
rect 22878 25230 22930 25282
rect 27806 25230 27858 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 14702 24894 14754 24946
rect 14926 24894 14978 24946
rect 17726 24894 17778 24946
rect 18622 24894 18674 24946
rect 19182 24894 19234 24946
rect 23326 24894 23378 24946
rect 17614 24782 17666 24834
rect 18398 24782 18450 24834
rect 18734 24782 18786 24834
rect 4286 24670 4338 24722
rect 11566 24670 11618 24722
rect 15038 24670 15090 24722
rect 17838 24670 17890 24722
rect 18286 24670 18338 24722
rect 19854 24670 19906 24722
rect 22990 24670 23042 24722
rect 25230 24670 25282 24722
rect 37662 24670 37714 24722
rect 12350 24558 12402 24610
rect 14478 24558 14530 24610
rect 15486 24558 15538 24610
rect 20526 24558 20578 24610
rect 22654 24558 22706 24610
rect 23774 24558 23826 24610
rect 26014 24558 26066 24610
rect 28142 24558 28194 24610
rect 28590 24558 28642 24610
rect 1934 24446 1986 24498
rect 40014 24446 40066 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 21422 23998 21474 24050
rect 25342 23998 25394 24050
rect 12574 23886 12626 23938
rect 13918 23886 13970 23938
rect 21982 23886 22034 23938
rect 25902 23886 25954 23938
rect 26238 23886 26290 23938
rect 27358 23886 27410 23938
rect 12910 23774 12962 23826
rect 14142 23774 14194 23826
rect 14366 23774 14418 23826
rect 14478 23774 14530 23826
rect 17390 23774 17442 23826
rect 25230 23774 25282 23826
rect 27582 23774 27634 23826
rect 12798 23662 12850 23714
rect 13582 23662 13634 23714
rect 13806 23662 13858 23714
rect 17726 23662 17778 23714
rect 21310 23662 21362 23714
rect 21534 23662 21586 23714
rect 25454 23662 25506 23714
rect 26126 23662 26178 23714
rect 26350 23662 26402 23714
rect 26574 23662 26626 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 26350 23326 26402 23378
rect 26574 23326 26626 23378
rect 13806 23214 13858 23266
rect 4286 23102 4338 23154
rect 14478 23102 14530 23154
rect 15038 23102 15090 23154
rect 20302 23102 20354 23154
rect 26238 23102 26290 23154
rect 11678 22990 11730 23042
rect 17390 22990 17442 23042
rect 19518 22990 19570 23042
rect 20750 22990 20802 23042
rect 1934 22878 1986 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 17950 22430 18002 22482
rect 24222 22430 24274 22482
rect 40014 22430 40066 22482
rect 16718 22318 16770 22370
rect 17166 22318 17218 22370
rect 17726 22318 17778 22370
rect 18286 22318 18338 22370
rect 18734 22318 18786 22370
rect 21310 22318 21362 22370
rect 37662 22318 37714 22370
rect 17054 22206 17106 22258
rect 18062 22206 18114 22258
rect 18846 22206 18898 22258
rect 22094 22206 22146 22258
rect 14366 22094 14418 22146
rect 16830 22094 16882 22146
rect 18958 22094 19010 22146
rect 24670 22094 24722 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 16494 21758 16546 21810
rect 16830 21758 16882 21810
rect 22878 21758 22930 21810
rect 12014 21646 12066 21698
rect 15150 21646 15202 21698
rect 17838 21646 17890 21698
rect 18174 21646 18226 21698
rect 19070 21646 19122 21698
rect 19518 21646 19570 21698
rect 19630 21646 19682 21698
rect 22094 21646 22146 21698
rect 22990 21646 23042 21698
rect 23326 21646 23378 21698
rect 23438 21646 23490 21698
rect 27134 21646 27186 21698
rect 27246 21646 27298 21698
rect 27582 21646 27634 21698
rect 27694 21646 27746 21698
rect 11342 21534 11394 21586
rect 14366 21534 14418 21586
rect 14590 21534 14642 21586
rect 14702 21534 14754 21586
rect 15262 21534 15314 21586
rect 16158 21534 16210 21586
rect 17950 21534 18002 21586
rect 18846 21534 18898 21586
rect 21646 21534 21698 21586
rect 22318 21534 22370 21586
rect 22430 21534 22482 21586
rect 22654 21534 22706 21586
rect 26126 21534 26178 21586
rect 26350 21534 26402 21586
rect 26798 21534 26850 21586
rect 26910 21534 26962 21586
rect 27918 21534 27970 21586
rect 37662 21534 37714 21586
rect 14142 21422 14194 21474
rect 15598 21422 15650 21474
rect 21870 21422 21922 21474
rect 25230 21422 25282 21474
rect 26574 21422 26626 21474
rect 40014 21422 40066 21474
rect 14814 21310 14866 21362
rect 19518 21310 19570 21362
rect 23438 21310 23490 21362
rect 25454 21310 25506 21362
rect 25790 21310 25842 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 20862 20974 20914 21026
rect 40014 20862 40066 20914
rect 14142 20750 14194 20802
rect 14366 20750 14418 20802
rect 19966 20750 20018 20802
rect 20190 20750 20242 20802
rect 20526 20750 20578 20802
rect 21870 20750 21922 20802
rect 37662 20750 37714 20802
rect 13918 20638 13970 20690
rect 15374 20638 15426 20690
rect 20750 20638 20802 20690
rect 25454 20638 25506 20690
rect 14254 20526 14306 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 11902 20078 11954 20130
rect 14478 20078 14530 20130
rect 16830 20078 16882 20130
rect 18174 20078 18226 20130
rect 21870 20078 21922 20130
rect 26126 20078 26178 20130
rect 11230 19966 11282 20018
rect 15486 19966 15538 20018
rect 15710 19966 15762 20018
rect 16606 19966 16658 20018
rect 17614 19966 17666 20018
rect 17950 19966 18002 20018
rect 18510 19966 18562 20018
rect 25454 19966 25506 20018
rect 37662 19966 37714 20018
rect 14030 19854 14082 19906
rect 15934 19854 15986 19906
rect 28254 19854 28306 19906
rect 28702 19854 28754 19906
rect 40014 19854 40066 19906
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 14926 19406 14978 19458
rect 15374 19406 15426 19458
rect 17166 19294 17218 19346
rect 24222 19294 24274 19346
rect 28366 19294 28418 19346
rect 15934 19182 15986 19234
rect 16942 19182 16994 19234
rect 17950 19182 18002 19234
rect 19966 19182 20018 19234
rect 21422 19182 21474 19234
rect 24670 19182 24722 19234
rect 25454 19182 25506 19234
rect 14702 19070 14754 19122
rect 15262 19070 15314 19122
rect 17502 19070 17554 19122
rect 18174 19070 18226 19122
rect 18510 19070 18562 19122
rect 19630 19070 19682 19122
rect 20190 19070 20242 19122
rect 20638 19070 20690 19122
rect 22094 19070 22146 19122
rect 26238 19070 26290 19122
rect 14814 18958 14866 19010
rect 15374 18958 15426 19010
rect 16270 18958 16322 19010
rect 18622 18958 18674 19010
rect 19294 18958 19346 19010
rect 29262 18958 29314 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 14030 18622 14082 18674
rect 20302 18622 20354 18674
rect 20526 18622 20578 18674
rect 21870 18622 21922 18674
rect 26126 18622 26178 18674
rect 27134 18622 27186 18674
rect 14366 18510 14418 18562
rect 16606 18510 16658 18562
rect 21310 18510 21362 18562
rect 14590 18398 14642 18450
rect 15598 18398 15650 18450
rect 15934 18398 15986 18450
rect 17950 18398 18002 18450
rect 18510 18398 18562 18450
rect 18846 18398 18898 18450
rect 19742 18398 19794 18450
rect 20078 18398 20130 18450
rect 20974 18398 21026 18450
rect 22542 18398 22594 18450
rect 22766 18398 22818 18450
rect 23102 18398 23154 18450
rect 23214 18398 23266 18450
rect 25790 18398 25842 18450
rect 26238 18398 26290 18450
rect 26462 18398 26514 18450
rect 26798 18398 26850 18450
rect 14926 18286 14978 18338
rect 16494 18286 16546 18338
rect 19182 18286 19234 18338
rect 20414 18286 20466 18338
rect 21422 18286 21474 18338
rect 16830 18174 16882 18226
rect 18846 18174 18898 18226
rect 21982 18174 22034 18226
rect 22206 18174 22258 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 14254 17838 14306 17890
rect 14814 17838 14866 17890
rect 15822 17838 15874 17890
rect 17166 17838 17218 17890
rect 21422 17838 21474 17890
rect 21758 17838 21810 17890
rect 1934 17726 1986 17778
rect 15486 17726 15538 17778
rect 40014 17726 40066 17778
rect 4286 17614 4338 17666
rect 15038 17614 15090 17666
rect 16494 17614 16546 17666
rect 17166 17614 17218 17666
rect 17614 17614 17666 17666
rect 19518 17614 19570 17666
rect 21982 17614 22034 17666
rect 22430 17614 22482 17666
rect 24782 17614 24834 17666
rect 26014 17614 26066 17666
rect 26574 17614 26626 17666
rect 37662 17614 37714 17666
rect 14478 17502 14530 17554
rect 14590 17502 14642 17554
rect 15598 17502 15650 17554
rect 16270 17502 16322 17554
rect 19294 17502 19346 17554
rect 19742 17502 19794 17554
rect 22318 17502 22370 17554
rect 25230 17502 25282 17554
rect 25454 17502 25506 17554
rect 25902 17502 25954 17554
rect 26238 17502 26290 17554
rect 19854 17390 19906 17442
rect 25118 17390 25170 17442
rect 25678 17390 25730 17442
rect 26462 17390 26514 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 14702 17054 14754 17106
rect 19630 17054 19682 17106
rect 19966 17054 20018 17106
rect 22094 17054 22146 17106
rect 12798 16942 12850 16994
rect 15038 16942 15090 16994
rect 15374 16942 15426 16994
rect 15598 16942 15650 16994
rect 15822 16942 15874 16994
rect 19854 16942 19906 16994
rect 26014 16942 26066 16994
rect 13582 16830 13634 16882
rect 14478 16830 14530 16882
rect 14814 16830 14866 16882
rect 19294 16830 19346 16882
rect 21870 16830 21922 16882
rect 23998 16830 24050 16882
rect 24334 16830 24386 16882
rect 24670 16830 24722 16882
rect 25230 16830 25282 16882
rect 28590 16830 28642 16882
rect 37662 16830 37714 16882
rect 10670 16718 10722 16770
rect 14030 16718 14082 16770
rect 15262 16718 15314 16770
rect 24222 16718 24274 16770
rect 28142 16718 28194 16770
rect 40014 16718 40066 16770
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 18398 16270 18450 16322
rect 1934 16158 1986 16210
rect 15710 16158 15762 16210
rect 25006 16158 25058 16210
rect 27134 16158 27186 16210
rect 4286 16046 4338 16098
rect 14142 16046 14194 16098
rect 14702 16046 14754 16098
rect 15598 16046 15650 16098
rect 18734 16046 18786 16098
rect 18958 16046 19010 16098
rect 20078 16046 20130 16098
rect 20302 16046 20354 16098
rect 20750 16046 20802 16098
rect 24222 16046 24274 16098
rect 27582 16046 27634 16098
rect 14366 15934 14418 15986
rect 15934 15934 15986 15986
rect 16158 15934 16210 15986
rect 14590 15822 14642 15874
rect 15150 15822 15202 15874
rect 20190 15822 20242 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 15710 15486 15762 15538
rect 18398 15486 18450 15538
rect 20302 15486 20354 15538
rect 16158 15374 16210 15426
rect 16382 15374 16434 15426
rect 19406 15374 19458 15426
rect 19630 15374 19682 15426
rect 22990 15374 23042 15426
rect 13918 15262 13970 15314
rect 14702 15262 14754 15314
rect 15486 15262 15538 15314
rect 18286 15262 18338 15314
rect 18510 15262 18562 15314
rect 18846 15262 18898 15314
rect 19966 15262 20018 15314
rect 23662 15262 23714 15314
rect 24222 15262 24274 15314
rect 11006 15150 11058 15202
rect 13134 15150 13186 15202
rect 14254 15150 14306 15202
rect 16046 15150 16098 15202
rect 19518 15150 19570 15202
rect 20862 15150 20914 15202
rect 14366 15038 14418 15090
rect 14590 15038 14642 15090
rect 19070 15038 19122 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 15262 14702 15314 14754
rect 15374 14702 15426 14754
rect 14254 14590 14306 14642
rect 16606 14590 16658 14642
rect 18734 14590 18786 14642
rect 15038 14478 15090 14530
rect 15934 14478 15986 14530
rect 21646 14478 21698 14530
rect 22430 14478 22482 14530
rect 14366 14366 14418 14418
rect 14590 14366 14642 14418
rect 14926 14366 14978 14418
rect 19182 14254 19234 14306
rect 21870 14254 21922 14306
rect 22206 14254 22258 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 16718 13918 16770 13970
rect 14142 13806 14194 13858
rect 19630 13806 19682 13858
rect 13470 13694 13522 13746
rect 18958 13694 19010 13746
rect 22206 13694 22258 13746
rect 16270 13582 16322 13634
rect 21758 13582 21810 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 40238 5966 40290 6018
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 22318 5182 22370 5234
rect 21310 5070 21362 5122
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 21870 4286 21922 4338
rect 22766 4062 22818 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 16942 3502 16994 3554
rect 21758 3502 21810 3554
rect 18510 3390 18562 3442
rect 15710 3278 15762 3330
rect 22430 3278 22482 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 18144 41200 18256 42000
rect 19488 41200 19600 42000
rect 22176 41200 22288 42000
rect 23520 41200 23632 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 18172 38162 18228 41200
rect 18172 38110 18174 38162
rect 18226 38110 18228 38162
rect 18172 38098 18228 38110
rect 19516 37492 19572 41200
rect 22204 38162 22260 41200
rect 23548 38276 23604 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 23548 38210 23604 38220
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 22204 38110 22206 38162
rect 22258 38110 22260 38162
rect 22204 38098 22260 38110
rect 19740 38052 19796 38062
rect 19628 38050 19796 38052
rect 19628 37998 19742 38050
rect 19794 37998 19796 38050
rect 19628 37996 19796 37998
rect 19628 37492 19684 37996
rect 19740 37986 19796 37996
rect 23660 38050 23716 38062
rect 23660 37998 23662 38050
rect 23714 37998 23716 38050
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20748 37492 20804 37502
rect 19628 37436 19908 37492
rect 19516 37426 19572 37436
rect 19740 37268 19796 37278
rect 18844 37266 19796 37268
rect 18844 37214 19742 37266
rect 19794 37214 19796 37266
rect 18844 37212 19796 37214
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 1932 27186 1988 27198
rect 1932 27134 1934 27186
rect 1986 27134 1988 27186
rect 1932 26292 1988 27134
rect 4284 27076 4340 27086
rect 4284 26982 4340 27020
rect 14028 27076 14084 27086
rect 1932 26226 1988 26236
rect 4284 26292 4340 26302
rect 4284 26198 4340 26236
rect 1932 26066 1988 26078
rect 1932 26014 1934 26066
rect 1986 26014 1988 26066
rect 1932 25620 1988 26014
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 1932 25554 1988 25564
rect 2044 25618 2100 25630
rect 2044 25566 2046 25618
rect 2098 25566 2100 25618
rect 2044 24948 2100 25566
rect 2044 24882 2100 24892
rect 4284 25506 4340 25518
rect 4284 25454 4286 25506
rect 4338 25454 4340 25506
rect 4284 24948 4340 25454
rect 14028 25394 14084 27020
rect 18844 26852 18900 37212
rect 19740 37202 19796 37212
rect 19852 36260 19908 37436
rect 20748 37398 20804 37436
rect 18844 26786 18900 26796
rect 18956 36204 19908 36260
rect 18956 26628 19012 36204
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20188 26852 20244 26862
rect 18620 26572 19012 26628
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 14700 26292 14756 26302
rect 14028 25342 14030 25394
rect 14082 25342 14084 25394
rect 14028 25330 14084 25342
rect 14252 25506 14308 25518
rect 14252 25454 14254 25506
rect 14306 25454 14308 25506
rect 4284 24882 4340 24892
rect 11564 24948 11620 24958
rect 14252 24948 14308 25454
rect 14700 25394 14756 26236
rect 17388 26290 17444 26302
rect 17388 26238 17390 26290
rect 17442 26238 17444 26290
rect 16940 26180 16996 26190
rect 17388 26180 17444 26238
rect 16940 26178 17444 26180
rect 16940 26126 16942 26178
rect 16994 26126 17444 26178
rect 16940 26124 17444 26126
rect 18172 26180 18228 26190
rect 14700 25342 14702 25394
rect 14754 25342 14756 25394
rect 14700 25330 14756 25342
rect 14924 25506 14980 25518
rect 14924 25454 14926 25506
rect 14978 25454 14980 25506
rect 14700 24948 14756 24958
rect 11620 24892 11732 24948
rect 11564 24882 11620 24892
rect 4284 24724 4340 24734
rect 11564 24724 11620 24734
rect 4284 24630 4340 24668
rect 11340 24722 11620 24724
rect 11340 24670 11566 24722
rect 11618 24670 11620 24722
rect 11340 24668 11620 24670
rect 1932 24500 1988 24510
rect 1932 24406 1988 24444
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4172 23604 4228 23614
rect 1932 22932 1988 22942
rect 1932 22838 1988 22876
rect 4172 19348 4228 23548
rect 4284 23156 4340 23166
rect 4284 23062 4340 23100
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 11340 21586 11396 24668
rect 11564 24658 11620 24668
rect 11676 23042 11732 24892
rect 14252 24882 14308 24892
rect 14364 24946 14756 24948
rect 14364 24894 14702 24946
rect 14754 24894 14756 24946
rect 14364 24892 14756 24894
rect 14364 24724 14420 24892
rect 14700 24882 14756 24892
rect 14924 24948 14980 25454
rect 14924 24854 14980 24892
rect 15708 25508 15764 25518
rect 13916 24668 14420 24724
rect 14476 24724 14532 24734
rect 12348 24612 12404 24622
rect 12348 24610 12628 24612
rect 12348 24558 12350 24610
rect 12402 24558 12628 24610
rect 12348 24556 12628 24558
rect 12348 24546 12404 24556
rect 12572 23938 12628 24556
rect 12572 23886 12574 23938
rect 12626 23886 12628 23938
rect 12572 23874 12628 23886
rect 13916 23938 13972 24668
rect 14476 24612 14532 24668
rect 13916 23886 13918 23938
rect 13970 23886 13972 23938
rect 13916 23874 13972 23886
rect 14364 24610 14532 24612
rect 14364 24558 14478 24610
rect 14530 24558 14532 24610
rect 14364 24556 14532 24558
rect 12908 23828 12964 23838
rect 12908 23734 12964 23772
rect 14140 23828 14196 23838
rect 14140 23734 14196 23772
rect 14364 23826 14420 24556
rect 14476 24546 14532 24556
rect 15036 24722 15092 24734
rect 15036 24670 15038 24722
rect 15090 24670 15092 24722
rect 14364 23774 14366 23826
rect 14418 23774 14420 23826
rect 14364 23762 14420 23774
rect 14476 23828 14532 23838
rect 14476 23734 14532 23772
rect 15036 23828 15092 24670
rect 15036 23762 15092 23772
rect 15484 24612 15540 24622
rect 15708 24612 15764 25452
rect 16940 25508 16996 26124
rect 18172 26086 18228 26124
rect 16492 25394 16548 25406
rect 16492 25342 16494 25394
rect 16546 25342 16548 25394
rect 16492 24948 16548 25342
rect 16940 25060 16996 25452
rect 16940 24994 16996 25004
rect 18620 25618 18676 26572
rect 18620 25566 18622 25618
rect 18674 25566 18676 25618
rect 16492 24882 16548 24892
rect 17724 24948 17780 24958
rect 17724 24854 17780 24892
rect 18620 24946 18676 25566
rect 19068 26180 19124 26190
rect 20188 26180 20244 26796
rect 21196 26290 21252 26302
rect 21196 26238 21198 26290
rect 21250 26238 21252 26290
rect 20300 26180 20356 26190
rect 19068 25618 19124 26124
rect 20076 26178 20356 26180
rect 20076 26126 20302 26178
rect 20354 26126 20356 26178
rect 20076 26124 20356 26126
rect 19964 25732 20020 25742
rect 19068 25566 19070 25618
rect 19122 25566 19124 25618
rect 19068 25554 19124 25566
rect 19628 25730 20020 25732
rect 19628 25678 19966 25730
rect 20018 25678 20020 25730
rect 19628 25676 20020 25678
rect 19628 25506 19684 25676
rect 19964 25666 20020 25676
rect 19628 25454 19630 25506
rect 19682 25454 19684 25506
rect 19628 25442 19684 25454
rect 19852 25394 19908 25406
rect 19852 25342 19854 25394
rect 19906 25342 19908 25394
rect 18956 25284 19012 25294
rect 19180 25284 19236 25294
rect 19852 25284 19908 25342
rect 19964 25396 20020 25406
rect 20076 25396 20132 26124
rect 20300 26114 20356 26124
rect 19964 25394 20132 25396
rect 19964 25342 19966 25394
rect 20018 25342 20132 25394
rect 19964 25340 20132 25342
rect 19964 25330 20020 25340
rect 18956 25190 19012 25228
rect 19068 25282 19236 25284
rect 19068 25230 19182 25282
rect 19234 25230 19236 25282
rect 19068 25228 19236 25230
rect 18620 24894 18622 24946
rect 18674 24894 18676 24946
rect 18620 24882 18676 24894
rect 18732 24948 18788 24958
rect 17612 24836 17668 24846
rect 17612 24742 17668 24780
rect 18396 24834 18452 24846
rect 18396 24782 18398 24834
rect 18450 24782 18452 24834
rect 15484 24610 15764 24612
rect 15484 24558 15486 24610
rect 15538 24558 15764 24610
rect 15484 24556 15764 24558
rect 17836 24722 17892 24734
rect 17836 24670 17838 24722
rect 17890 24670 17892 24722
rect 11676 22990 11678 23042
rect 11730 22990 11732 23042
rect 11676 22978 11732 22990
rect 12796 23714 12852 23726
rect 12796 23662 12798 23714
rect 12850 23662 12852 23714
rect 12012 22148 12068 22158
rect 12012 21698 12068 22092
rect 12012 21646 12014 21698
rect 12066 21646 12068 21698
rect 12012 21634 12068 21646
rect 11340 21534 11342 21586
rect 11394 21534 11396 21586
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 11340 20132 11396 21534
rect 11228 20076 11340 20132
rect 11228 20018 11284 20076
rect 11340 20066 11396 20076
rect 11900 20580 11956 20590
rect 11900 20130 11956 20524
rect 11900 20078 11902 20130
rect 11954 20078 11956 20130
rect 11900 20066 11956 20078
rect 11228 19966 11230 20018
rect 11282 19966 11284 20018
rect 11228 19954 11284 19966
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4172 19282 4228 19292
rect 12796 18228 12852 23662
rect 13580 23716 13636 23726
rect 13804 23716 13860 23726
rect 13580 23714 13748 23716
rect 13580 23662 13582 23714
rect 13634 23662 13748 23714
rect 13580 23660 13748 23662
rect 13580 23650 13636 23660
rect 13692 23268 13748 23660
rect 13804 23714 13972 23716
rect 13804 23662 13806 23714
rect 13858 23662 13972 23714
rect 13804 23660 13972 23662
rect 13804 23650 13860 23660
rect 13804 23268 13860 23278
rect 13692 23266 13860 23268
rect 13692 23214 13806 23266
rect 13858 23214 13860 23266
rect 13692 23212 13860 23214
rect 13804 23202 13860 23212
rect 13916 20692 13972 23660
rect 14476 23156 14532 23166
rect 15036 23156 15092 23166
rect 15484 23156 15540 24556
rect 17388 23828 17444 23838
rect 17388 23734 17444 23772
rect 17724 23716 17780 23726
rect 17724 23622 17780 23660
rect 14476 23154 15540 23156
rect 14476 23102 14478 23154
rect 14530 23102 15038 23154
rect 15090 23102 15540 23154
rect 14476 23100 15540 23102
rect 17388 23156 17444 23166
rect 14140 22596 14196 22606
rect 13692 20690 13972 20692
rect 13692 20638 13918 20690
rect 13970 20638 13972 20690
rect 13692 20636 13972 20638
rect 13692 19572 13748 20636
rect 13916 20626 13972 20636
rect 14028 22540 14140 22596
rect 14028 21252 14084 22540
rect 14140 22530 14196 22540
rect 14364 22148 14420 22158
rect 14476 22148 14532 23100
rect 15036 23090 15092 23100
rect 17388 23042 17444 23100
rect 17388 22990 17390 23042
rect 17442 22990 17444 23042
rect 17388 22978 17444 22990
rect 16716 22596 16772 22606
rect 16716 22370 16772 22540
rect 16716 22318 16718 22370
rect 16770 22318 16772 22370
rect 16716 22306 16772 22318
rect 17164 22372 17220 22382
rect 17724 22372 17780 22382
rect 17164 22370 17780 22372
rect 17164 22318 17166 22370
rect 17218 22318 17726 22370
rect 17778 22318 17780 22370
rect 17164 22316 17780 22318
rect 17052 22258 17108 22270
rect 17052 22206 17054 22258
rect 17106 22206 17108 22258
rect 14364 22146 14532 22148
rect 14364 22094 14366 22146
rect 14418 22094 14532 22146
rect 14364 22092 14532 22094
rect 14364 22082 14420 22092
rect 14364 21588 14420 21598
rect 14140 21586 14420 21588
rect 14140 21534 14366 21586
rect 14418 21534 14420 21586
rect 14140 21532 14420 21534
rect 14140 21474 14196 21532
rect 14364 21522 14420 21532
rect 14140 21422 14142 21474
rect 14194 21422 14196 21474
rect 14140 21410 14196 21422
rect 14028 21196 14420 21252
rect 14028 20188 14084 21196
rect 14140 20804 14196 20814
rect 14140 20710 14196 20748
rect 14364 20802 14420 21196
rect 14364 20750 14366 20802
rect 14418 20750 14420 20802
rect 14364 20738 14420 20750
rect 14476 20692 14532 22092
rect 16828 22148 16884 22158
rect 16828 22054 16884 22092
rect 16492 21812 16548 21822
rect 15148 21810 16548 21812
rect 15148 21758 16494 21810
rect 16546 21758 16548 21810
rect 15148 21756 16548 21758
rect 15148 21698 15204 21756
rect 15148 21646 15150 21698
rect 15202 21646 15204 21698
rect 15148 21634 15204 21646
rect 14588 21588 14644 21598
rect 14700 21588 14756 21598
rect 14588 21586 14756 21588
rect 14588 21534 14590 21586
rect 14642 21534 14702 21586
rect 14754 21534 14756 21586
rect 14588 21532 14756 21534
rect 14588 21522 14644 21532
rect 14252 20580 14308 20590
rect 14252 20486 14308 20524
rect 13692 19506 13748 19516
rect 13916 20132 14084 20188
rect 14140 20132 14196 20142
rect 14476 20132 14532 20636
rect 12796 18162 12852 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 13916 17892 13972 20132
rect 14196 20130 14532 20132
rect 14196 20078 14478 20130
rect 14530 20078 14532 20130
rect 14196 20076 14532 20078
rect 14028 19906 14084 19918
rect 14028 19854 14030 19906
rect 14082 19854 14084 19906
rect 14028 19460 14084 19854
rect 14028 19394 14084 19404
rect 14028 18676 14084 18686
rect 14028 18582 14084 18620
rect 13916 17826 13972 17836
rect 1932 17778 1988 17790
rect 1932 17726 1934 17778
rect 1986 17726 1988 17778
rect 1932 16884 1988 17726
rect 4284 17668 4340 17678
rect 4284 17574 4340 17612
rect 10668 17668 10724 17678
rect 1932 16818 1988 16828
rect 10668 16996 10724 17612
rect 10668 16770 10724 16940
rect 12796 17220 12852 17230
rect 12796 16994 12852 17164
rect 12796 16942 12798 16994
rect 12850 16942 12852 16994
rect 12796 16930 12852 16942
rect 10668 16718 10670 16770
rect 10722 16718 10724 16770
rect 10668 16706 10724 16718
rect 13580 16882 13636 16894
rect 13580 16830 13582 16882
rect 13634 16830 13636 16882
rect 13580 16772 13636 16830
rect 14028 16772 14084 16782
rect 14140 16772 14196 20076
rect 14476 20038 14532 20076
rect 14588 19572 14644 19582
rect 14364 18562 14420 18574
rect 14364 18510 14366 18562
rect 14418 18510 14420 18562
rect 14252 18228 14308 18238
rect 14252 17890 14308 18172
rect 14252 17838 14254 17890
rect 14306 17838 14308 17890
rect 14252 17826 14308 17838
rect 14364 17444 14420 18510
rect 14588 18450 14644 19516
rect 14700 19236 14756 21532
rect 15260 21588 15316 21598
rect 15260 21494 15316 21532
rect 15596 21474 15652 21486
rect 15596 21422 15598 21474
rect 15650 21422 15652 21474
rect 14812 21362 14868 21374
rect 14812 21310 14814 21362
rect 14866 21310 14868 21362
rect 14812 20020 14868 21310
rect 15596 20804 15652 21422
rect 15372 20692 15428 20702
rect 15372 20598 15428 20636
rect 14812 19954 14868 19964
rect 15484 20020 15540 20030
rect 15484 19926 15540 19964
rect 15372 19572 15428 19582
rect 14924 19460 14980 19470
rect 14924 19366 14980 19404
rect 15372 19458 15428 19516
rect 15372 19406 15374 19458
rect 15426 19406 15428 19458
rect 15372 19394 15428 19406
rect 14700 19122 14756 19180
rect 14700 19070 14702 19122
rect 14754 19070 14756 19122
rect 14700 19058 14756 19070
rect 15260 19122 15316 19134
rect 15260 19070 15262 19122
rect 15314 19070 15316 19122
rect 14812 19010 14868 19022
rect 14812 18958 14814 19010
rect 14866 18958 14868 19010
rect 14812 18900 14868 18958
rect 15260 18900 15316 19070
rect 14812 18844 15316 18900
rect 15372 19010 15428 19022
rect 15372 18958 15374 19010
rect 15426 18958 15428 19010
rect 14812 18676 14868 18844
rect 14812 18610 14868 18620
rect 14588 18398 14590 18450
rect 14642 18398 14644 18450
rect 14588 18386 14644 18398
rect 14924 18338 14980 18350
rect 14924 18286 14926 18338
rect 14978 18286 14980 18338
rect 14812 17892 14868 17902
rect 14812 17798 14868 17836
rect 14364 17378 14420 17388
rect 14476 17554 14532 17566
rect 14476 17502 14478 17554
rect 14530 17502 14532 17554
rect 14476 17108 14532 17502
rect 13580 16770 14196 16772
rect 13580 16718 14030 16770
rect 14082 16718 14196 16770
rect 13580 16716 14196 16718
rect 14252 17052 14532 17108
rect 14588 17554 14644 17566
rect 14588 17502 14590 17554
rect 14642 17502 14644 17554
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 1932 16210 1988 16222
rect 1932 16158 1934 16210
rect 1986 16158 1988 16210
rect 1932 15540 1988 16158
rect 4284 16100 4340 16110
rect 4284 16006 4340 16044
rect 11004 16100 11060 16110
rect 1932 15474 1988 15484
rect 11004 15202 11060 16044
rect 13468 15316 13524 15326
rect 11004 15150 11006 15202
rect 11058 15150 11060 15202
rect 11004 15138 11060 15150
rect 13132 15204 13188 15214
rect 13132 15110 13188 15148
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 13468 13746 13524 15260
rect 13916 15316 13972 15326
rect 14028 15316 14084 16716
rect 14140 16100 14196 16110
rect 14140 16006 14196 16044
rect 14252 15988 14308 17052
rect 14476 16882 14532 16894
rect 14476 16830 14478 16882
rect 14530 16830 14532 16882
rect 14476 16772 14532 16830
rect 14476 16706 14532 16716
rect 14588 16100 14644 17502
rect 14812 17220 14868 17230
rect 14700 17108 14756 17118
rect 14812 17108 14868 17164
rect 14700 17106 14868 17108
rect 14700 17054 14702 17106
rect 14754 17054 14868 17106
rect 14700 17052 14868 17054
rect 14700 17042 14756 17052
rect 14812 16882 14868 16894
rect 14812 16830 14814 16882
rect 14866 16830 14868 16882
rect 14812 16212 14868 16830
rect 14812 16146 14868 16156
rect 14476 16044 14644 16100
rect 14700 16100 14756 16110
rect 14364 15988 14420 15998
rect 14252 15986 14420 15988
rect 14252 15934 14366 15986
rect 14418 15934 14420 15986
rect 14252 15932 14420 15934
rect 14364 15428 14420 15932
rect 14364 15362 14420 15372
rect 13972 15260 14084 15316
rect 13916 15222 13972 15260
rect 14252 15204 14308 15214
rect 14476 15204 14532 16044
rect 14700 16006 14756 16044
rect 14588 15874 14644 15886
rect 14588 15822 14590 15874
rect 14642 15822 14644 15874
rect 14588 15316 14644 15822
rect 14700 15316 14756 15326
rect 14588 15314 14756 15316
rect 14588 15262 14702 15314
rect 14754 15262 14756 15314
rect 14588 15260 14756 15262
rect 14700 15250 14756 15260
rect 14476 15148 14644 15204
rect 14252 15110 14308 15148
rect 14364 15092 14420 15102
rect 14252 14642 14308 14654
rect 14252 14590 14254 14642
rect 14306 14590 14308 14642
rect 14140 13860 14196 13870
rect 14252 13860 14308 14590
rect 14364 14418 14420 15036
rect 14588 15090 14644 15148
rect 14588 15038 14590 15090
rect 14642 15038 14644 15090
rect 14588 15026 14644 15038
rect 14924 15092 14980 18286
rect 15372 18004 15428 18958
rect 15596 18900 15652 20748
rect 15708 20018 15764 21756
rect 16492 21746 16548 21756
rect 16828 21812 16884 21822
rect 16828 21718 16884 21756
rect 16156 21588 16212 21598
rect 16156 21494 16212 21532
rect 17052 21364 17108 22206
rect 17052 21298 17108 21308
rect 16828 20132 16884 20142
rect 16828 20038 16884 20076
rect 15708 19966 15710 20018
rect 15762 19966 15764 20018
rect 15708 19460 15764 19966
rect 16604 20020 16660 20030
rect 16604 19926 16660 19964
rect 15932 19908 15988 19918
rect 15708 19394 15764 19404
rect 15820 19906 15988 19908
rect 15820 19854 15934 19906
rect 15986 19854 15988 19906
rect 15820 19852 15988 19854
rect 15596 18834 15652 18844
rect 15820 19124 15876 19852
rect 15932 19842 15988 19852
rect 17164 19346 17220 22316
rect 17724 22306 17780 22316
rect 17836 22148 17892 24670
rect 18284 24724 18340 24734
rect 18396 24724 18452 24782
rect 18284 24722 18452 24724
rect 18284 24670 18286 24722
rect 18338 24670 18452 24722
rect 18284 24668 18452 24670
rect 18732 24834 18788 24892
rect 18732 24782 18734 24834
rect 18786 24782 18788 24834
rect 18284 24658 18340 24668
rect 18620 23940 18676 23950
rect 18396 23716 18452 23726
rect 17948 23044 18004 23054
rect 17948 22482 18004 22988
rect 17948 22430 17950 22482
rect 18002 22430 18004 22482
rect 17948 22418 18004 22430
rect 18284 22370 18340 22382
rect 18284 22318 18286 22370
rect 18338 22318 18340 22370
rect 18060 22260 18116 22270
rect 18060 22166 18116 22204
rect 17612 22092 17892 22148
rect 18172 22148 18228 22158
rect 17612 21364 17668 22092
rect 18172 21924 18228 22092
rect 17612 21298 17668 21308
rect 17724 21868 18228 21924
rect 17612 20020 17668 20030
rect 17612 19926 17668 19964
rect 17164 19294 17166 19346
rect 17218 19294 17220 19346
rect 15932 19236 15988 19246
rect 15932 19142 15988 19180
rect 16940 19234 16996 19246
rect 16940 19182 16942 19234
rect 16994 19182 16996 19234
rect 15372 17938 15428 17948
rect 15596 18452 15652 18462
rect 15820 18452 15876 19068
rect 16940 19124 16996 19182
rect 16940 19058 16996 19068
rect 16268 19010 16324 19022
rect 16268 18958 16270 19010
rect 16322 18958 16324 19010
rect 16268 18564 16324 18958
rect 16604 18564 16660 18574
rect 16268 18562 16660 18564
rect 16268 18510 16606 18562
rect 16658 18510 16660 18562
rect 16268 18508 16660 18510
rect 15596 18450 15876 18452
rect 15596 18398 15598 18450
rect 15650 18398 15876 18450
rect 15596 18396 15876 18398
rect 15932 18450 15988 18462
rect 15932 18398 15934 18450
rect 15986 18398 15988 18450
rect 15484 17780 15540 17790
rect 15260 17778 15540 17780
rect 15260 17726 15486 17778
rect 15538 17726 15540 17778
rect 15260 17724 15540 17726
rect 15036 17666 15092 17678
rect 15036 17614 15038 17666
rect 15090 17614 15092 17666
rect 15036 17332 15092 17614
rect 15036 17266 15092 17276
rect 15260 17108 15316 17724
rect 15484 17714 15540 17724
rect 15596 17554 15652 18396
rect 15932 18340 15988 18398
rect 16604 18452 16660 18508
rect 16604 18386 16660 18396
rect 16492 18340 16548 18350
rect 15932 18338 16548 18340
rect 15932 18286 16494 18338
rect 16546 18286 16548 18338
rect 15932 18284 16548 18286
rect 15596 17502 15598 17554
rect 15650 17502 15652 17554
rect 15596 17490 15652 17502
rect 15708 18228 15764 18238
rect 15036 17052 15316 17108
rect 15484 17444 15540 17454
rect 15036 16994 15092 17052
rect 15036 16942 15038 16994
rect 15090 16942 15092 16994
rect 15036 16930 15092 16942
rect 15372 16996 15428 17006
rect 15372 16902 15428 16940
rect 15260 16772 15316 16782
rect 15484 16772 15540 17388
rect 15596 17332 15652 17342
rect 15596 16996 15652 17276
rect 15708 16996 15764 18172
rect 15820 17892 15876 17902
rect 15932 17892 15988 18284
rect 16492 18274 16548 18284
rect 16828 18226 16884 18238
rect 16828 18174 16830 18226
rect 16882 18174 16884 18226
rect 16492 18004 16548 18014
rect 15820 17890 15988 17892
rect 15820 17838 15822 17890
rect 15874 17838 15988 17890
rect 15820 17836 15988 17838
rect 16268 17892 16324 17902
rect 15820 17826 15876 17836
rect 16268 17554 16324 17836
rect 16268 17502 16270 17554
rect 16322 17502 16324 17554
rect 16268 17490 16324 17502
rect 16492 17668 16548 17948
rect 16828 18004 16884 18174
rect 16828 17938 16884 17948
rect 17164 17890 17220 19294
rect 17164 17838 17166 17890
rect 17218 17838 17220 17890
rect 17164 17826 17220 17838
rect 17500 19122 17556 19134
rect 17500 19070 17502 19122
rect 17554 19070 17556 19122
rect 15820 16996 15876 17006
rect 15708 16994 15876 16996
rect 15708 16942 15822 16994
rect 15874 16942 15876 16994
rect 15708 16940 15876 16942
rect 15596 16902 15652 16940
rect 15820 16930 15876 16940
rect 15596 16772 15652 16782
rect 15484 16716 15596 16772
rect 15260 16678 15316 16716
rect 15260 16100 15316 16110
rect 15148 15874 15204 15886
rect 15148 15822 15150 15874
rect 15202 15822 15204 15874
rect 15148 15316 15204 15822
rect 15036 15092 15092 15102
rect 14924 15036 15036 15092
rect 15036 15026 15092 15036
rect 15036 14530 15092 14542
rect 15036 14478 15038 14530
rect 15090 14478 15092 14530
rect 14364 14366 14366 14418
rect 14418 14366 14420 14418
rect 14364 14354 14420 14366
rect 14588 14420 14644 14430
rect 14924 14420 14980 14430
rect 14588 14418 14980 14420
rect 14588 14366 14590 14418
rect 14642 14366 14926 14418
rect 14978 14366 14980 14418
rect 14588 14364 14980 14366
rect 14588 14354 14644 14364
rect 14924 14354 14980 14364
rect 14140 13858 14308 13860
rect 14140 13806 14142 13858
rect 14194 13806 14308 13858
rect 14140 13804 14308 13806
rect 14140 13794 14196 13804
rect 13468 13694 13470 13746
rect 13522 13694 13524 13746
rect 13468 13682 13524 13694
rect 15036 13524 15092 14478
rect 15148 14308 15204 15260
rect 15260 14754 15316 16044
rect 15596 16100 15652 16716
rect 16492 16324 16548 17612
rect 17164 17668 17220 17678
rect 17164 17574 17220 17612
rect 17500 17108 17556 19070
rect 17612 18452 17668 18462
rect 17612 17666 17668 18396
rect 17612 17614 17614 17666
rect 17666 17614 17668 17666
rect 17612 17602 17668 17614
rect 17500 17042 17556 17052
rect 17724 16996 17780 21868
rect 17836 21700 17892 21710
rect 17836 20132 17892 21644
rect 18172 21698 18228 21868
rect 18284 21812 18340 22318
rect 18284 21746 18340 21756
rect 18172 21646 18174 21698
rect 18226 21646 18228 21698
rect 18172 21634 18228 21646
rect 17836 19796 17892 20076
rect 17948 21588 18004 21598
rect 17948 20018 18004 21532
rect 18396 20356 18452 23660
rect 18172 20300 18452 20356
rect 18508 21812 18564 21822
rect 18172 20130 18228 20300
rect 18508 20188 18564 21756
rect 18172 20078 18174 20130
rect 18226 20078 18228 20130
rect 18172 20066 18228 20078
rect 18284 20132 18564 20188
rect 18620 20188 18676 23884
rect 18732 23828 18788 24782
rect 19068 23940 19124 25228
rect 19180 25218 19236 25228
rect 19628 25228 19908 25284
rect 19180 25060 19236 25070
rect 19180 24946 19236 25004
rect 19180 24894 19182 24946
rect 19234 24894 19236 24946
rect 19180 24882 19236 24894
rect 19628 24948 19684 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19628 24882 19684 24892
rect 19852 24724 19908 24734
rect 20300 24724 20356 24734
rect 19852 24722 20300 24724
rect 19852 24670 19854 24722
rect 19906 24670 20300 24722
rect 19852 24668 20300 24670
rect 19852 24658 19908 24668
rect 19180 23940 19236 23950
rect 19068 23884 19180 23940
rect 19180 23874 19236 23884
rect 18732 23762 18788 23772
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 18732 23156 18788 23166
rect 18732 22370 18788 23100
rect 20300 23154 20356 24668
rect 21196 24724 21252 26238
rect 21980 26178 22036 26190
rect 21980 26126 21982 26178
rect 22034 26126 22036 26178
rect 21980 25618 22036 26126
rect 21980 25566 21982 25618
rect 22034 25566 22036 25618
rect 21980 25554 22036 25566
rect 22540 25564 23156 25620
rect 22540 25506 22596 25564
rect 22540 25454 22542 25506
rect 22594 25454 22596 25506
rect 22540 25442 22596 25454
rect 23100 25508 23156 25564
rect 23212 25508 23268 25518
rect 23100 25506 23268 25508
rect 23100 25454 23214 25506
rect 23266 25454 23268 25506
rect 23100 25452 23268 25454
rect 23212 25442 23268 25452
rect 23548 25508 23604 25518
rect 22988 25394 23044 25406
rect 22988 25342 22990 25394
rect 23042 25342 23044 25394
rect 21196 24658 21252 24668
rect 21644 25284 21700 25294
rect 20524 24612 20580 24622
rect 20524 24610 21140 24612
rect 20524 24558 20526 24610
rect 20578 24558 21140 24610
rect 20524 24556 21140 24558
rect 20524 24546 20580 24556
rect 21084 24164 21140 24556
rect 21084 24108 21476 24164
rect 21420 24050 21476 24108
rect 21420 23998 21422 24050
rect 21474 23998 21476 24050
rect 21420 23986 21476 23998
rect 21532 23940 21588 23950
rect 21308 23716 21364 23726
rect 21308 23714 21476 23716
rect 21308 23662 21310 23714
rect 21362 23662 21476 23714
rect 21308 23660 21476 23662
rect 21308 23650 21364 23660
rect 20300 23102 20302 23154
rect 20354 23102 20356 23154
rect 19516 23044 19572 23054
rect 20300 23044 20356 23102
rect 20748 23044 20804 23054
rect 20300 23042 20804 23044
rect 20300 22990 20750 23042
rect 20802 22990 20804 23042
rect 20300 22988 20804 22990
rect 19516 22950 19572 22988
rect 18732 22318 18734 22370
rect 18786 22318 18788 22370
rect 18732 22306 18788 22318
rect 20748 22372 20804 22988
rect 21308 22372 21364 22382
rect 20748 22370 21364 22372
rect 20748 22318 21310 22370
rect 21362 22318 21364 22370
rect 20748 22316 21364 22318
rect 18844 22260 18900 22270
rect 18844 22166 18900 22204
rect 18956 22148 19012 22158
rect 18956 22146 19124 22148
rect 18956 22094 18958 22146
rect 19010 22094 19124 22146
rect 18956 22092 19124 22094
rect 18956 22082 19012 22092
rect 19068 21700 19124 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19628 21812 19684 21822
rect 19516 21700 19572 21710
rect 19068 21698 19572 21700
rect 19068 21646 19070 21698
rect 19122 21646 19518 21698
rect 19570 21646 19572 21698
rect 19068 21644 19572 21646
rect 19068 21634 19124 21644
rect 18844 21588 18900 21598
rect 18844 21494 18900 21532
rect 19404 20188 19460 21644
rect 19516 21634 19572 21644
rect 19628 21698 19684 21756
rect 19628 21646 19630 21698
rect 19682 21646 19684 21698
rect 19628 21634 19684 21646
rect 20188 21812 20244 21822
rect 19516 21364 19572 21374
rect 19516 21270 19572 21308
rect 19964 20804 20020 20814
rect 19964 20710 20020 20748
rect 20188 20802 20244 21756
rect 20188 20750 20190 20802
rect 20242 20750 20244 20802
rect 20188 20738 20244 20750
rect 20524 21588 20580 21598
rect 20748 21588 20804 21598
rect 20524 20802 20580 21532
rect 20524 20750 20526 20802
rect 20578 20750 20580 20802
rect 20524 20738 20580 20750
rect 20636 21532 20748 21588
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 18620 20132 18788 20188
rect 19404 20132 19572 20188
rect 17948 19966 17950 20018
rect 18002 19966 18004 20018
rect 17948 19954 18004 19966
rect 17836 19740 18116 19796
rect 17836 19348 17892 19358
rect 17836 18452 17892 19292
rect 17948 19234 18004 19246
rect 17948 19182 17950 19234
rect 18002 19182 18004 19234
rect 17948 18676 18004 19182
rect 18060 19124 18116 19740
rect 18060 19058 18116 19068
rect 18172 19124 18228 19134
rect 18284 19124 18340 20132
rect 18508 20018 18564 20030
rect 18508 19966 18510 20018
rect 18562 19966 18564 20018
rect 18508 19348 18564 19966
rect 18508 19282 18564 19292
rect 18172 19122 18340 19124
rect 18172 19070 18174 19122
rect 18226 19070 18340 19122
rect 18172 19068 18340 19070
rect 18508 19124 18564 19134
rect 18172 19058 18228 19068
rect 18508 19030 18564 19068
rect 18620 19010 18676 19022
rect 18620 18958 18622 19010
rect 18674 18958 18676 19010
rect 18508 18900 18564 18910
rect 17948 18620 18340 18676
rect 17948 18452 18004 18462
rect 17836 18450 18004 18452
rect 17836 18398 17950 18450
rect 18002 18398 18004 18450
rect 17836 18396 18004 18398
rect 17948 18386 18004 18396
rect 17724 16930 17780 16940
rect 15708 16212 15764 16222
rect 15708 16118 15764 16156
rect 15596 16006 15652 16044
rect 15484 15988 15540 15998
rect 15260 14702 15262 14754
rect 15314 14702 15316 14754
rect 15260 14690 15316 14702
rect 15372 15932 15484 15988
rect 15372 14754 15428 15932
rect 15484 15922 15540 15932
rect 15932 15986 15988 15998
rect 15932 15934 15934 15986
rect 15986 15934 15988 15986
rect 15932 15652 15988 15934
rect 16156 15988 16212 15998
rect 16156 15894 16212 15932
rect 15708 15596 16324 15652
rect 15708 15538 15764 15596
rect 15708 15486 15710 15538
rect 15762 15486 15764 15538
rect 15708 15474 15764 15486
rect 16156 15428 16212 15438
rect 16156 15334 16212 15372
rect 15484 15314 15540 15326
rect 15484 15262 15486 15314
rect 15538 15262 15540 15314
rect 15484 15204 15540 15262
rect 16044 15204 16100 15214
rect 15484 15202 16100 15204
rect 15484 15150 16046 15202
rect 16098 15150 16100 15202
rect 15484 15148 16100 15150
rect 16044 15138 16100 15148
rect 15372 14702 15374 14754
rect 15426 14702 15428 14754
rect 15372 14690 15428 14702
rect 16268 14644 16324 15596
rect 16380 15428 16436 15438
rect 16492 15428 16548 16268
rect 18284 15540 18340 18620
rect 18508 18450 18564 18844
rect 18508 18398 18510 18450
rect 18562 18398 18564 18450
rect 18508 18386 18564 18398
rect 18508 18228 18564 18238
rect 18620 18228 18676 18958
rect 18564 18172 18676 18228
rect 18508 18162 18564 18172
rect 18620 18004 18676 18014
rect 18732 18004 18788 20132
rect 19292 19012 19348 19022
rect 18844 19010 19348 19012
rect 18844 18958 19294 19010
rect 19346 18958 19348 19010
rect 18844 18956 19348 18958
rect 18844 18452 18900 18956
rect 19292 18946 19348 18956
rect 19516 18452 19572 20132
rect 19964 19234 20020 19246
rect 19964 19182 19966 19234
rect 20018 19182 20020 19234
rect 19628 19124 19684 19134
rect 19628 19030 19684 19068
rect 19964 19012 20020 19182
rect 19964 18946 20020 18956
rect 20188 19124 20244 19134
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19740 18452 19796 18462
rect 19516 18450 19796 18452
rect 19516 18398 19742 18450
rect 19794 18398 19796 18450
rect 19516 18396 19796 18398
rect 18844 18386 18900 18396
rect 19180 18338 19236 18350
rect 19180 18286 19182 18338
rect 19234 18286 19236 18338
rect 18676 17948 18788 18004
rect 18844 18226 18900 18238
rect 18844 18174 18846 18226
rect 18898 18174 18900 18226
rect 18620 17938 18676 17948
rect 18396 16324 18452 16334
rect 18396 16230 18452 16268
rect 18732 16098 18788 16110
rect 18732 16046 18734 16098
rect 18786 16046 18788 16098
rect 18396 15540 18452 15550
rect 18284 15538 18452 15540
rect 18284 15486 18398 15538
rect 18450 15486 18452 15538
rect 18284 15484 18452 15486
rect 16380 15426 16548 15428
rect 16380 15374 16382 15426
rect 16434 15374 16548 15426
rect 16380 15372 16548 15374
rect 18396 15428 18452 15484
rect 16380 15362 16436 15372
rect 18396 15362 18452 15372
rect 18284 15314 18340 15326
rect 18284 15262 18286 15314
rect 18338 15262 18340 15314
rect 18284 15204 18340 15262
rect 18508 15316 18564 15326
rect 18732 15316 18788 16046
rect 18564 15260 18788 15316
rect 18508 15222 18564 15260
rect 18284 15138 18340 15148
rect 16604 14644 16660 14654
rect 16268 14642 16660 14644
rect 16268 14590 16606 14642
rect 16658 14590 16660 14642
rect 16268 14588 16660 14590
rect 16604 14578 16660 14588
rect 18732 14642 18788 15260
rect 18844 15988 18900 18174
rect 19180 18004 19236 18286
rect 19180 17938 19236 17948
rect 19516 18228 19572 18238
rect 19516 17666 19572 18172
rect 19516 17614 19518 17666
rect 19570 17614 19572 17666
rect 19516 17602 19572 17614
rect 19628 17892 19684 17902
rect 19292 17556 19348 17566
rect 19292 17462 19348 17500
rect 19628 17106 19684 17836
rect 19740 17554 19796 18396
rect 19740 17502 19742 17554
rect 19794 17502 19796 17554
rect 19740 17490 19796 17502
rect 20076 18450 20132 18462
rect 20076 18398 20078 18450
rect 20130 18398 20132 18450
rect 20076 17556 20132 18398
rect 20188 17780 20244 19068
rect 20636 19122 20692 21532
rect 20748 21522 20804 21532
rect 20860 21028 20916 21038
rect 20860 20934 20916 20972
rect 20748 20692 20804 20702
rect 20748 20598 20804 20636
rect 21308 20188 21364 22316
rect 21420 22148 21476 23660
rect 21420 22082 21476 22092
rect 21532 23714 21588 23884
rect 21532 23662 21534 23714
rect 21586 23662 21588 23714
rect 21308 20132 21476 20188
rect 21420 19236 21476 20132
rect 21420 19142 21476 19180
rect 20636 19070 20638 19122
rect 20690 19070 20692 19122
rect 20300 19012 20356 19022
rect 20300 18674 20356 18956
rect 20300 18622 20302 18674
rect 20354 18622 20356 18674
rect 20300 18610 20356 18622
rect 20524 18676 20580 18686
rect 20524 18582 20580 18620
rect 20412 18340 20468 18350
rect 20412 18246 20468 18284
rect 20636 18228 20692 19070
rect 21532 18676 21588 23662
rect 21644 21588 21700 25228
rect 21868 25282 21924 25294
rect 21868 25230 21870 25282
rect 21922 25230 21924 25282
rect 21868 24724 21924 25230
rect 22092 25284 22148 25294
rect 22652 25284 22708 25294
rect 22876 25284 22932 25294
rect 22092 25190 22148 25228
rect 22204 25282 22708 25284
rect 22204 25230 22654 25282
rect 22706 25230 22708 25282
rect 22204 25228 22708 25230
rect 21868 23940 21924 24668
rect 21868 23874 21924 23884
rect 21980 23940 22036 23950
rect 22204 23940 22260 25228
rect 22652 25218 22708 25228
rect 22764 25228 22876 25284
rect 22652 24612 22708 24622
rect 22764 24612 22820 25228
rect 22876 25190 22932 25228
rect 22988 25172 23044 25342
rect 23436 25396 23492 25406
rect 23436 25302 23492 25340
rect 23548 25172 23604 25452
rect 23660 25284 23716 37998
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 24556 31948 24612 37998
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 24108 31892 24612 31948
rect 24108 26178 24164 31892
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 26236 26402 26292 26414
rect 26236 26350 26238 26402
rect 26290 26350 26292 26402
rect 26012 26292 26068 26302
rect 25900 26290 26068 26292
rect 25900 26238 26014 26290
rect 26066 26238 26068 26290
rect 25900 26236 26068 26238
rect 24668 26180 24724 26190
rect 24108 26126 24110 26178
rect 24162 26126 24164 26178
rect 24108 25396 24164 26126
rect 24108 25330 24164 25340
rect 24556 26178 24724 26180
rect 24556 26126 24670 26178
rect 24722 26126 24724 26178
rect 24556 26124 24724 26126
rect 24556 25506 24612 26124
rect 24668 26114 24724 26124
rect 24556 25454 24558 25506
rect 24610 25454 24612 25506
rect 23660 25218 23716 25228
rect 22988 25116 23604 25172
rect 23324 24946 23380 25116
rect 23324 24894 23326 24946
rect 23378 24894 23380 24946
rect 23324 24882 23380 24894
rect 22652 24610 22820 24612
rect 22652 24558 22654 24610
rect 22706 24558 22820 24610
rect 22652 24556 22820 24558
rect 22988 24722 23044 24734
rect 22988 24670 22990 24722
rect 23042 24670 23044 24722
rect 22652 24546 22708 24556
rect 21980 23938 22260 23940
rect 21980 23886 21982 23938
rect 22034 23886 22260 23938
rect 21980 23884 22260 23886
rect 21980 23874 22036 23884
rect 22988 23716 23044 24670
rect 23772 24612 23828 24622
rect 23772 24518 23828 24556
rect 24556 24612 24612 25454
rect 25228 25396 25284 25406
rect 25228 25394 25396 25396
rect 25228 25342 25230 25394
rect 25282 25342 25396 25394
rect 25228 25340 25396 25342
rect 25228 25330 25284 25340
rect 25228 24724 25284 24734
rect 24556 24546 24612 24556
rect 25116 24722 25284 24724
rect 25116 24670 25230 24722
rect 25282 24670 25284 24722
rect 25116 24668 25284 24670
rect 25116 24612 25172 24668
rect 25228 24658 25284 24668
rect 22092 22258 22148 22270
rect 22092 22206 22094 22258
rect 22146 22206 22148 22258
rect 22092 21698 22148 22206
rect 22876 21812 22932 21822
rect 22876 21718 22932 21756
rect 22092 21646 22094 21698
rect 22146 21646 22148 21698
rect 22092 21634 22148 21646
rect 22988 21700 23044 23660
rect 24220 22484 24276 22494
rect 24220 21924 24276 22428
rect 24668 22148 24724 22158
rect 25116 22148 25172 24556
rect 25340 24050 25396 25340
rect 25340 23998 25342 24050
rect 25394 23998 25396 24050
rect 25340 23986 25396 23998
rect 25900 23938 25956 26236
rect 26012 26226 26068 26236
rect 26236 25620 26292 26350
rect 26236 25554 26292 25564
rect 26348 26290 26404 26302
rect 26348 26238 26350 26290
rect 26402 26238 26404 26290
rect 26348 25508 26404 26238
rect 37660 26290 37716 26302
rect 37660 26238 37662 26290
rect 37714 26238 37716 26290
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 37660 25732 37716 26238
rect 37660 25666 37716 25676
rect 39900 26178 39956 26190
rect 39900 26126 39902 26178
rect 39954 26126 39956 26178
rect 27356 25620 27412 25630
rect 27356 25526 27412 25564
rect 39900 25620 39956 26126
rect 39900 25554 39956 25564
rect 40012 25618 40068 25630
rect 40012 25566 40014 25618
rect 40066 25566 40068 25618
rect 26348 25060 26404 25452
rect 37884 25506 37940 25518
rect 37884 25454 37886 25506
rect 37938 25454 37940 25506
rect 27804 25282 27860 25294
rect 27804 25230 27806 25282
rect 27858 25230 27860 25282
rect 26348 25004 26740 25060
rect 26012 24610 26068 24622
rect 26012 24558 26014 24610
rect 26066 24558 26068 24610
rect 26012 24052 26068 24558
rect 26012 23996 26292 24052
rect 25900 23886 25902 23938
rect 25954 23886 25956 23938
rect 25900 23874 25956 23886
rect 26236 23938 26292 23996
rect 26236 23886 26238 23938
rect 26290 23886 26292 23938
rect 26236 23874 26292 23886
rect 25228 23828 25284 23838
rect 25228 23734 25284 23772
rect 25452 23714 25508 23726
rect 25452 23662 25454 23714
rect 25506 23662 25508 23714
rect 25452 23492 25508 23662
rect 25452 23426 25508 23436
rect 26124 23714 26180 23726
rect 26124 23662 26126 23714
rect 26178 23662 26180 23714
rect 26124 22596 26180 23662
rect 26348 23714 26404 23726
rect 26348 23662 26350 23714
rect 26402 23662 26404 23714
rect 26348 23604 26404 23662
rect 26348 23538 26404 23548
rect 26460 23716 26516 23726
rect 26348 23380 26404 23390
rect 26460 23380 26516 23660
rect 26348 23378 26516 23380
rect 26348 23326 26350 23378
rect 26402 23326 26516 23378
rect 26348 23324 26516 23326
rect 26572 23714 26628 23726
rect 26572 23662 26574 23714
rect 26626 23662 26628 23714
rect 26572 23378 26628 23662
rect 26572 23326 26574 23378
rect 26626 23326 26628 23378
rect 26348 23314 26404 23324
rect 26572 23314 26628 23326
rect 26236 23156 26292 23166
rect 26684 23156 26740 25004
rect 27804 24612 27860 25230
rect 37660 24722 37716 24734
rect 37660 24670 37662 24722
rect 37714 24670 37716 24722
rect 27804 24546 27860 24556
rect 28140 24610 28196 24622
rect 28140 24558 28142 24610
rect 28194 24558 28196 24610
rect 27356 23938 27412 23950
rect 27356 23886 27358 23938
rect 27410 23886 27412 23938
rect 27356 23716 27412 23886
rect 27580 23940 27636 23950
rect 27580 23826 27636 23884
rect 27580 23774 27582 23826
rect 27634 23774 27636 23826
rect 27580 23762 27636 23774
rect 27356 23650 27412 23660
rect 28140 23716 28196 24558
rect 28588 24612 28644 24622
rect 28588 24518 28644 24556
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 28140 23650 28196 23660
rect 37660 23716 37716 24670
rect 37884 23940 37940 25454
rect 40012 24948 40068 25566
rect 40012 24882 40068 24892
rect 40012 24498 40068 24510
rect 40012 24446 40014 24498
rect 40066 24446 40068 24498
rect 40012 24276 40068 24446
rect 40012 24210 40068 24220
rect 37884 23874 37940 23884
rect 37660 23650 37716 23660
rect 26236 23154 26740 23156
rect 26236 23102 26238 23154
rect 26290 23102 26740 23154
rect 26236 23100 26740 23102
rect 27244 23492 27300 23502
rect 26236 23090 26292 23100
rect 26124 22530 26180 22540
rect 25340 22148 25396 22158
rect 25116 22092 25340 22148
rect 24668 22054 24724 22092
rect 24220 21858 24276 21868
rect 23324 21700 23380 21710
rect 22988 21698 23380 21700
rect 22988 21646 22990 21698
rect 23042 21646 23326 21698
rect 23378 21646 23380 21698
rect 22988 21644 23380 21646
rect 22988 21634 23044 21644
rect 23324 21634 23380 21644
rect 23436 21700 23492 21710
rect 23436 21606 23492 21644
rect 24220 21700 24276 21710
rect 21644 21494 21700 21532
rect 22316 21586 22372 21598
rect 22316 21534 22318 21586
rect 22370 21534 22372 21586
rect 21868 21476 21924 21486
rect 21868 21382 21924 21420
rect 21868 20804 21924 20814
rect 21868 20130 21924 20748
rect 21868 20078 21870 20130
rect 21922 20078 21924 20130
rect 21868 20066 21924 20078
rect 22316 20692 22372 21534
rect 22428 21588 22484 21598
rect 22652 21588 22708 21598
rect 22428 21586 22708 21588
rect 22428 21534 22430 21586
rect 22482 21534 22654 21586
rect 22706 21534 22708 21586
rect 22428 21532 22708 21534
rect 22428 21522 22484 21532
rect 22652 21522 22708 21532
rect 23436 21364 23492 21374
rect 22092 19124 22148 19134
rect 21308 18562 21364 18574
rect 21308 18510 21310 18562
rect 21362 18510 21364 18562
rect 20636 18162 20692 18172
rect 20972 18450 21028 18462
rect 20972 18398 20974 18450
rect 21026 18398 21028 18450
rect 20972 18116 21028 18398
rect 21308 18452 21364 18510
rect 21308 18386 21364 18396
rect 21420 18340 21476 18350
rect 21532 18340 21588 18620
rect 21868 19122 22148 19124
rect 21868 19070 22094 19122
rect 22146 19070 22148 19122
rect 21868 19068 22148 19070
rect 21868 18674 21924 19068
rect 22092 19058 22148 19068
rect 21868 18622 21870 18674
rect 21922 18622 21924 18674
rect 21868 18610 21924 18622
rect 21420 18338 21588 18340
rect 21420 18286 21422 18338
rect 21474 18286 21588 18338
rect 21420 18284 21588 18286
rect 21420 18274 21476 18284
rect 21980 18228 22036 18238
rect 21980 18134 22036 18172
rect 22204 18228 22260 18238
rect 22204 18134 22260 18172
rect 21084 18116 21140 18126
rect 20972 18060 21084 18116
rect 21084 18050 21140 18060
rect 21420 18004 21476 18014
rect 20188 17714 20244 17724
rect 20300 17892 20356 17902
rect 19852 17444 19908 17482
rect 20076 17444 20132 17500
rect 20076 17388 20244 17444
rect 19852 17378 19908 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 17054 19630 17106
rect 19682 17054 19684 17106
rect 19628 17042 19684 17054
rect 19964 17108 20020 17118
rect 20188 17108 20244 17388
rect 19964 17106 20244 17108
rect 19964 17054 19966 17106
rect 20018 17054 20244 17106
rect 19964 17052 20244 17054
rect 19852 16996 19908 17006
rect 19852 16902 19908 16940
rect 19292 16884 19348 16894
rect 19292 16790 19348 16828
rect 19964 16324 20020 17052
rect 19628 16268 20020 16324
rect 20076 16884 20132 16894
rect 18844 15314 18900 15932
rect 18844 15262 18846 15314
rect 18898 15262 18900 15314
rect 18844 15250 18900 15262
rect 18956 16098 19012 16110
rect 18956 16046 18958 16098
rect 19010 16046 19012 16098
rect 18956 15204 19012 16046
rect 19404 15876 19460 15886
rect 19404 15426 19460 15820
rect 19404 15374 19406 15426
rect 19458 15374 19460 15426
rect 19404 15362 19460 15374
rect 19628 15426 19684 16268
rect 20076 16098 20132 16828
rect 20076 16046 20078 16098
rect 20130 16046 20132 16098
rect 20076 16034 20132 16046
rect 20300 16098 20356 17836
rect 21420 17890 21476 17948
rect 21420 17838 21422 17890
rect 21474 17838 21476 17890
rect 21420 17826 21476 17838
rect 21756 17892 21812 17902
rect 21756 17798 21812 17836
rect 21980 17668 22036 17678
rect 22036 17612 22148 17668
rect 21980 17574 22036 17612
rect 22092 17106 22148 17612
rect 22092 17054 22094 17106
rect 22146 17054 22148 17106
rect 22092 17042 22148 17054
rect 22316 17556 22372 20636
rect 22764 21362 23492 21364
rect 22764 21310 23438 21362
rect 23490 21310 23492 21362
rect 22764 21308 23492 21310
rect 22540 18452 22596 18462
rect 22428 17668 22484 17678
rect 22540 17668 22596 18396
rect 22764 18450 22820 21308
rect 23436 21298 23492 21308
rect 23212 21140 23268 21150
rect 22764 18398 22766 18450
rect 22818 18398 22820 18450
rect 22764 18386 22820 18398
rect 23100 18450 23156 18462
rect 23100 18398 23102 18450
rect 23154 18398 23156 18450
rect 23100 17892 23156 18398
rect 23212 18450 23268 21084
rect 24220 19348 24276 21644
rect 25228 21476 25284 21486
rect 25228 21382 25284 21420
rect 25340 20692 25396 22092
rect 27132 21700 27188 21710
rect 27132 21606 27188 21644
rect 27244 21700 27300 23436
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 37660 22372 37716 22382
rect 37660 22278 37716 22316
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 27580 21700 27636 21710
rect 27244 21698 27636 21700
rect 27244 21646 27246 21698
rect 27298 21646 27582 21698
rect 27634 21646 27636 21698
rect 27244 21644 27636 21646
rect 26124 21588 26180 21598
rect 26012 21586 26180 21588
rect 26012 21534 26126 21586
rect 26178 21534 26180 21586
rect 26012 21532 26180 21534
rect 25452 21362 25508 21374
rect 25452 21310 25454 21362
rect 25506 21310 25508 21362
rect 25452 21028 25508 21310
rect 25452 20962 25508 20972
rect 25788 21362 25844 21374
rect 25788 21310 25790 21362
rect 25842 21310 25844 21362
rect 25452 20692 25508 20702
rect 25340 20690 25508 20692
rect 25340 20638 25454 20690
rect 25506 20638 25508 20690
rect 25340 20636 25508 20638
rect 24220 19254 24276 19292
rect 25452 20018 25508 20636
rect 25452 19966 25454 20018
rect 25506 19966 25508 20018
rect 24668 19236 24724 19246
rect 24668 19142 24724 19180
rect 25340 19236 25396 19246
rect 25452 19236 25508 19966
rect 25396 19234 25508 19236
rect 25396 19182 25454 19234
rect 25506 19182 25508 19234
rect 25396 19180 25508 19182
rect 23212 18398 23214 18450
rect 23266 18398 23268 18450
rect 23212 18228 23268 18398
rect 23212 18162 23268 18172
rect 24780 18340 24836 18350
rect 23100 17826 23156 17836
rect 22484 17612 22596 17668
rect 24780 17666 24836 18284
rect 24780 17614 24782 17666
rect 24834 17614 24836 17666
rect 22428 17574 22484 17612
rect 24780 17602 24836 17614
rect 22316 16996 22372 17500
rect 22316 16930 22372 16940
rect 22988 17556 23044 17566
rect 21868 16882 21924 16894
rect 21868 16830 21870 16882
rect 21922 16830 21924 16882
rect 20300 16046 20302 16098
rect 20354 16046 20356 16098
rect 20188 15876 20244 15886
rect 20188 15782 20244 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20300 15538 20356 16046
rect 20300 15486 20302 15538
rect 20354 15486 20356 15538
rect 20300 15474 20356 15486
rect 20748 16098 20804 16110
rect 20748 16046 20750 16098
rect 20802 16046 20804 16098
rect 19628 15374 19630 15426
rect 19682 15374 19684 15426
rect 19628 15362 19684 15374
rect 19964 15316 20020 15326
rect 19964 15222 20020 15260
rect 18956 15138 19012 15148
rect 19516 15202 19572 15214
rect 19516 15150 19518 15202
rect 19570 15150 19572 15202
rect 19068 15092 19124 15102
rect 19068 14998 19124 15036
rect 18732 14590 18734 14642
rect 18786 14590 18788 14642
rect 18732 14578 18788 14590
rect 15148 14242 15204 14252
rect 15932 14530 15988 14542
rect 15932 14478 15934 14530
rect 15986 14478 15988 14530
rect 15932 14308 15988 14478
rect 15932 14242 15988 14252
rect 16716 14308 16772 14318
rect 16716 13970 16772 14252
rect 19180 14308 19236 14318
rect 19180 14214 19236 14252
rect 16716 13918 16718 13970
rect 16770 13918 16772 13970
rect 16716 13906 16772 13918
rect 19516 13860 19572 15150
rect 20748 14532 20804 16046
rect 20860 15204 20916 15214
rect 20860 15110 20916 15148
rect 21868 15204 21924 16830
rect 22988 15426 23044 17500
rect 25228 17556 25284 17566
rect 25228 17462 25284 17500
rect 23996 17444 24052 17454
rect 23996 16882 24052 17388
rect 24220 17444 24276 17454
rect 24220 16996 24276 17388
rect 25116 17442 25172 17454
rect 25116 17390 25118 17442
rect 25170 17390 25172 17442
rect 25116 16996 25172 17390
rect 24220 16940 24388 16996
rect 23996 16830 23998 16882
rect 24050 16830 24052 16882
rect 23996 16818 24052 16830
rect 24332 16882 24388 16940
rect 25116 16930 25172 16940
rect 24332 16830 24334 16882
rect 24386 16830 24388 16882
rect 24332 16818 24388 16830
rect 24668 16884 24724 16894
rect 24668 16790 24724 16828
rect 25228 16884 25284 16894
rect 25340 16884 25396 19180
rect 25452 19170 25508 19180
rect 25788 18450 25844 21310
rect 25788 18398 25790 18450
rect 25842 18398 25844 18450
rect 25788 18386 25844 18398
rect 26012 18004 26068 21532
rect 26124 21522 26180 21532
rect 26348 21586 26404 21598
rect 26348 21534 26350 21586
rect 26402 21534 26404 21586
rect 26348 21028 26404 21534
rect 26796 21588 26852 21598
rect 26796 21494 26852 21532
rect 26908 21586 26964 21598
rect 26908 21534 26910 21586
rect 26962 21534 26964 21586
rect 26348 20962 26404 20972
rect 26572 21474 26628 21486
rect 26572 21422 26574 21474
rect 26626 21422 26628 21474
rect 26572 20188 26628 21422
rect 26124 20132 26628 20188
rect 26124 20130 26180 20132
rect 26124 20078 26126 20130
rect 26178 20078 26180 20130
rect 26124 20066 26180 20078
rect 26908 19348 26964 21534
rect 26348 19292 26964 19348
rect 26236 19122 26292 19134
rect 26236 19070 26238 19122
rect 26290 19070 26292 19122
rect 26124 18676 26180 18686
rect 26236 18676 26292 19070
rect 26124 18674 26292 18676
rect 26124 18622 26126 18674
rect 26178 18622 26292 18674
rect 26124 18620 26292 18622
rect 26124 18610 26180 18620
rect 26236 18452 26292 18462
rect 26348 18452 26404 19292
rect 27132 18676 27188 18686
rect 27244 18676 27300 21644
rect 27580 21634 27636 21644
rect 27692 21698 27748 21710
rect 27692 21646 27694 21698
rect 27746 21646 27748 21698
rect 27692 20244 27748 21646
rect 28364 21700 28420 21710
rect 27916 21588 27972 21598
rect 27916 21494 27972 21532
rect 27692 20178 27748 20188
rect 28252 20244 28308 20254
rect 28252 19906 28308 20188
rect 28252 19854 28254 19906
rect 28306 19854 28308 19906
rect 28252 19842 28308 19854
rect 28364 19346 28420 21644
rect 37660 21588 37716 21598
rect 37660 21494 37716 21532
rect 40012 21588 40068 21598
rect 40012 21474 40068 21532
rect 40012 21422 40014 21474
rect 40066 21422 40068 21474
rect 40012 21410 40068 21422
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 40012 20916 40068 20926
rect 40012 20822 40068 20860
rect 37660 20802 37716 20814
rect 37660 20750 37662 20802
rect 37714 20750 37716 20802
rect 37660 20244 37716 20750
rect 37660 20178 37716 20188
rect 40012 20132 40068 20142
rect 37660 20018 37716 20030
rect 37660 19966 37662 20018
rect 37714 19966 37716 20018
rect 28700 19908 28756 19918
rect 28364 19294 28366 19346
rect 28418 19294 28420 19346
rect 28364 19282 28420 19294
rect 28588 19906 28756 19908
rect 28588 19854 28702 19906
rect 28754 19854 28756 19906
rect 28588 19852 28756 19854
rect 27132 18674 27300 18676
rect 27132 18622 27134 18674
rect 27186 18622 27300 18674
rect 27132 18620 27300 18622
rect 28588 19012 28644 19852
rect 28700 19842 28756 19852
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 37660 19348 37716 19966
rect 40012 19906 40068 20076
rect 40012 19854 40014 19906
rect 40066 19854 40068 19906
rect 40012 19842 40068 19854
rect 37660 19282 37716 19292
rect 27132 18610 27188 18620
rect 26236 18450 26404 18452
rect 26236 18398 26238 18450
rect 26290 18398 26404 18450
rect 26236 18396 26404 18398
rect 26460 18450 26516 18462
rect 26460 18398 26462 18450
rect 26514 18398 26516 18450
rect 26236 18386 26292 18396
rect 26460 18004 26516 18398
rect 26012 17948 26516 18004
rect 26796 18450 26852 18462
rect 26796 18398 26798 18450
rect 26850 18398 26852 18450
rect 26012 17780 26068 17790
rect 25900 17668 25956 17678
rect 25452 17554 25508 17566
rect 25452 17502 25454 17554
rect 25506 17502 25508 17554
rect 25452 17108 25508 17502
rect 25900 17554 25956 17612
rect 26012 17666 26068 17724
rect 26012 17614 26014 17666
rect 26066 17614 26068 17666
rect 26012 17602 26068 17614
rect 25900 17502 25902 17554
rect 25954 17502 25956 17554
rect 25900 17490 25956 17502
rect 26236 17556 26292 17566
rect 26236 17462 26292 17500
rect 25676 17444 25732 17454
rect 25676 17350 25732 17388
rect 25452 17042 25508 17052
rect 26348 17108 26404 17948
rect 26796 17780 26852 18398
rect 26572 17724 26796 17780
rect 26572 17666 26628 17724
rect 26796 17714 26852 17724
rect 26572 17614 26574 17666
rect 26626 17614 26628 17666
rect 26572 17602 26628 17614
rect 27132 17668 27188 17678
rect 26348 17042 26404 17052
rect 26460 17442 26516 17454
rect 26460 17390 26462 17442
rect 26514 17390 26516 17442
rect 26012 16996 26068 17006
rect 26012 16902 26068 16940
rect 25228 16882 25396 16884
rect 25228 16830 25230 16882
rect 25282 16830 25396 16882
rect 25228 16828 25396 16830
rect 26460 16884 26516 17390
rect 24220 16770 24276 16782
rect 24220 16718 24222 16770
rect 24274 16718 24276 16770
rect 24220 16324 24276 16718
rect 24220 16268 25060 16324
rect 25004 16210 25060 16268
rect 25004 16158 25006 16210
rect 25058 16158 25060 16210
rect 25004 16146 25060 16158
rect 22988 15374 22990 15426
rect 23042 15374 23044 15426
rect 22988 15362 23044 15374
rect 24220 16100 24276 16110
rect 21868 15138 21924 15148
rect 23660 15316 23716 15326
rect 24220 15316 24276 16044
rect 25228 16100 25284 16828
rect 26460 16818 26516 16828
rect 27132 16210 27188 17612
rect 28140 16884 28196 16894
rect 28588 16884 28644 18956
rect 29260 19012 29316 19022
rect 29260 18918 29316 18956
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 37660 17668 37716 17678
rect 37660 17574 37716 17612
rect 40012 17556 40068 17726
rect 40012 17490 40068 17500
rect 28140 16770 28196 16828
rect 28140 16718 28142 16770
rect 28194 16718 28196 16770
rect 28140 16706 28196 16718
rect 28476 16882 28644 16884
rect 28476 16830 28590 16882
rect 28642 16830 28644 16882
rect 28476 16828 28644 16830
rect 27132 16158 27134 16210
rect 27186 16158 27188 16210
rect 27132 16146 27188 16158
rect 25228 16034 25284 16044
rect 27580 16100 27636 16110
rect 27580 16006 27636 16044
rect 28364 16100 28420 16110
rect 28476 16100 28532 16828
rect 28588 16818 28644 16828
rect 37660 16884 37716 16894
rect 37660 16790 37716 16828
rect 40012 16884 40068 16894
rect 40012 16770 40068 16828
rect 40012 16718 40014 16770
rect 40066 16718 40068 16770
rect 40012 16706 40068 16718
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 28420 16044 28532 16100
rect 28364 16034 28420 16044
rect 23660 15314 24276 15316
rect 23660 15262 23662 15314
rect 23714 15262 24222 15314
rect 24274 15262 24276 15314
rect 23660 15260 24276 15262
rect 20748 14466 20804 14476
rect 21644 14532 21700 14542
rect 21756 14532 21812 14542
rect 21644 14530 21756 14532
rect 21644 14478 21646 14530
rect 21698 14478 21756 14530
rect 21644 14476 21756 14478
rect 21644 14466 21700 14476
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19628 13860 19684 13870
rect 19516 13858 19684 13860
rect 19516 13806 19630 13858
rect 19682 13806 19684 13858
rect 19516 13804 19684 13806
rect 19628 13794 19684 13804
rect 18956 13748 19012 13758
rect 18956 13654 19012 13692
rect 15036 13458 15092 13468
rect 16268 13634 16324 13646
rect 16268 13582 16270 13634
rect 16322 13582 16324 13634
rect 16268 13524 16324 13582
rect 21756 13634 21812 14476
rect 22428 14532 22484 14542
rect 22428 14438 22484 14476
rect 21756 13582 21758 13634
rect 21810 13582 21812 13634
rect 16268 13458 16324 13468
rect 16940 13524 16996 13534
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 16940 3554 16996 13468
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 21756 8428 21812 13582
rect 21308 8372 21812 8428
rect 21868 14306 21924 14318
rect 22204 14308 22260 14318
rect 21868 14254 21870 14306
rect 21922 14254 21924 14306
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20860 5236 20916 5246
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 16940 3502 16942 3554
rect 16994 3502 16996 3554
rect 16940 3490 16996 3502
rect 16156 3444 16212 3454
rect 15708 3332 15764 3342
rect 15484 3330 15764 3332
rect 15484 3278 15710 3330
rect 15762 3278 15764 3330
rect 15484 3276 15764 3278
rect 15484 800 15540 3276
rect 15708 3266 15764 3276
rect 16156 800 16212 3388
rect 18508 3444 18564 3454
rect 18508 3350 18564 3388
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20860 800 20916 5180
rect 21308 5122 21364 8372
rect 21308 5070 21310 5122
rect 21362 5070 21364 5122
rect 21308 5058 21364 5070
rect 21868 4338 21924 14254
rect 21868 4286 21870 4338
rect 21922 4286 21924 4338
rect 21868 4274 21924 4286
rect 21980 14306 22260 14308
rect 21980 14254 22206 14306
rect 22258 14254 22260 14306
rect 21980 14252 22260 14254
rect 21532 4116 21588 4126
rect 21980 4116 22036 14252
rect 22204 14242 22260 14252
rect 22204 13748 22260 13758
rect 22204 13654 22260 13692
rect 23660 13748 23716 15260
rect 24220 15250 24276 15260
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 23660 13682 23716 13692
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 40236 6018 40292 6030
rect 40236 5966 40238 6018
rect 40290 5966 40292 6018
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 40236 5460 40292 5966
rect 40236 5394 40292 5404
rect 22316 5236 22372 5246
rect 22316 5142 22372 5180
rect 21532 800 21588 4060
rect 21756 4060 22036 4116
rect 22764 4116 22820 4126
rect 21756 3554 21812 4060
rect 22764 4022 22820 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 21756 3502 21758 3554
rect 21810 3502 21812 3554
rect 21756 3490 21812 3502
rect 22428 3332 22484 3342
rect 22204 3330 22484 3332
rect 22204 3278 22430 3330
rect 22482 3278 22484 3330
rect 22204 3276 22484 3278
rect 22204 800 22260 3276
rect 22428 3266 22484 3276
rect 15456 0 15568 800
rect 16128 0 16240 800
rect 20832 0 20944 800
rect 21504 0 21616 800
rect 22176 0 22288 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 23548 38220 23604 38276
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 19516 37436 19572 37492
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4284 27074 4340 27076
rect 4284 27022 4286 27074
rect 4286 27022 4338 27074
rect 4338 27022 4340 27074
rect 4284 27020 4340 27022
rect 14028 27020 14084 27076
rect 1932 26236 1988 26292
rect 4284 26290 4340 26292
rect 4284 26238 4286 26290
rect 4286 26238 4338 26290
rect 4338 26238 4340 26290
rect 4284 26236 4340 26238
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 1932 25564 1988 25620
rect 2044 24892 2100 24948
rect 20748 37490 20804 37492
rect 20748 37438 20750 37490
rect 20750 37438 20802 37490
rect 20802 37438 20804 37490
rect 20748 37436 20804 37438
rect 18844 26796 18900 26852
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 20188 26796 20244 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 14700 26236 14756 26292
rect 4284 24892 4340 24948
rect 18172 26178 18228 26180
rect 18172 26126 18174 26178
rect 18174 26126 18226 26178
rect 18226 26126 18228 26178
rect 18172 26124 18228 26126
rect 11564 24892 11620 24948
rect 4284 24722 4340 24724
rect 4284 24670 4286 24722
rect 4286 24670 4338 24722
rect 4338 24670 4340 24722
rect 4284 24668 4340 24670
rect 1932 24498 1988 24500
rect 1932 24446 1934 24498
rect 1934 24446 1986 24498
rect 1986 24446 1988 24498
rect 1932 24444 1988 24446
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4172 23548 4228 23604
rect 1932 22930 1988 22932
rect 1932 22878 1934 22930
rect 1934 22878 1986 22930
rect 1986 22878 1988 22930
rect 1932 22876 1988 22878
rect 4284 23154 4340 23156
rect 4284 23102 4286 23154
rect 4286 23102 4338 23154
rect 4338 23102 4340 23154
rect 4284 23100 4340 23102
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 14252 24892 14308 24948
rect 14924 24946 14980 24948
rect 14924 24894 14926 24946
rect 14926 24894 14978 24946
rect 14978 24894 14980 24946
rect 14924 24892 14980 24894
rect 15708 25506 15764 25508
rect 15708 25454 15710 25506
rect 15710 25454 15762 25506
rect 15762 25454 15764 25506
rect 15708 25452 15764 25454
rect 14476 24668 14532 24724
rect 12908 23826 12964 23828
rect 12908 23774 12910 23826
rect 12910 23774 12962 23826
rect 12962 23774 12964 23826
rect 12908 23772 12964 23774
rect 14140 23826 14196 23828
rect 14140 23774 14142 23826
rect 14142 23774 14194 23826
rect 14194 23774 14196 23826
rect 14140 23772 14196 23774
rect 14476 23826 14532 23828
rect 14476 23774 14478 23826
rect 14478 23774 14530 23826
rect 14530 23774 14532 23826
rect 14476 23772 14532 23774
rect 15036 23772 15092 23828
rect 16940 25452 16996 25508
rect 16940 25004 16996 25060
rect 16492 24892 16548 24948
rect 17724 24946 17780 24948
rect 17724 24894 17726 24946
rect 17726 24894 17778 24946
rect 17778 24894 17780 24946
rect 17724 24892 17780 24894
rect 19068 26124 19124 26180
rect 18956 25282 19012 25284
rect 18956 25230 18958 25282
rect 18958 25230 19010 25282
rect 19010 25230 19012 25282
rect 18956 25228 19012 25230
rect 18732 24892 18788 24948
rect 17612 24834 17668 24836
rect 17612 24782 17614 24834
rect 17614 24782 17666 24834
rect 17666 24782 17668 24834
rect 17612 24780 17668 24782
rect 12012 22092 12068 22148
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 11340 20076 11396 20132
rect 11900 20524 11956 20580
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4172 19292 4228 19348
rect 17388 23826 17444 23828
rect 17388 23774 17390 23826
rect 17390 23774 17442 23826
rect 17442 23774 17444 23826
rect 17388 23772 17444 23774
rect 17724 23714 17780 23716
rect 17724 23662 17726 23714
rect 17726 23662 17778 23714
rect 17778 23662 17780 23714
rect 17724 23660 17780 23662
rect 17388 23100 17444 23156
rect 14140 22540 14196 22596
rect 16716 22540 16772 22596
rect 14140 20802 14196 20804
rect 14140 20750 14142 20802
rect 14142 20750 14194 20802
rect 14194 20750 14196 20802
rect 14140 20748 14196 20750
rect 16828 22146 16884 22148
rect 16828 22094 16830 22146
rect 16830 22094 16882 22146
rect 16882 22094 16884 22146
rect 16828 22092 16884 22094
rect 14476 20636 14532 20692
rect 14252 20578 14308 20580
rect 14252 20526 14254 20578
rect 14254 20526 14306 20578
rect 14306 20526 14308 20578
rect 14252 20524 14308 20526
rect 13692 19516 13748 19572
rect 12796 18172 12852 18228
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 14140 20076 14196 20132
rect 14028 19404 14084 19460
rect 14028 18674 14084 18676
rect 14028 18622 14030 18674
rect 14030 18622 14082 18674
rect 14082 18622 14084 18674
rect 14028 18620 14084 18622
rect 13916 17836 13972 17892
rect 4284 17666 4340 17668
rect 4284 17614 4286 17666
rect 4286 17614 4338 17666
rect 4338 17614 4340 17666
rect 4284 17612 4340 17614
rect 10668 17612 10724 17668
rect 1932 16828 1988 16884
rect 10668 16940 10724 16996
rect 12796 17164 12852 17220
rect 14588 19516 14644 19572
rect 14252 18172 14308 18228
rect 15260 21586 15316 21588
rect 15260 21534 15262 21586
rect 15262 21534 15314 21586
rect 15314 21534 15316 21586
rect 15260 21532 15316 21534
rect 15596 20748 15652 20804
rect 15372 20690 15428 20692
rect 15372 20638 15374 20690
rect 15374 20638 15426 20690
rect 15426 20638 15428 20690
rect 15372 20636 15428 20638
rect 14812 19964 14868 20020
rect 15484 20018 15540 20020
rect 15484 19966 15486 20018
rect 15486 19966 15538 20018
rect 15538 19966 15540 20018
rect 15484 19964 15540 19966
rect 15372 19516 15428 19572
rect 14924 19458 14980 19460
rect 14924 19406 14926 19458
rect 14926 19406 14978 19458
rect 14978 19406 14980 19458
rect 14924 19404 14980 19406
rect 14700 19180 14756 19236
rect 14812 18620 14868 18676
rect 14812 17890 14868 17892
rect 14812 17838 14814 17890
rect 14814 17838 14866 17890
rect 14866 17838 14868 17890
rect 14812 17836 14868 17838
rect 14364 17388 14420 17444
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4284 16098 4340 16100
rect 4284 16046 4286 16098
rect 4286 16046 4338 16098
rect 4338 16046 4340 16098
rect 4284 16044 4340 16046
rect 11004 16044 11060 16100
rect 1932 15484 1988 15540
rect 13468 15260 13524 15316
rect 13132 15202 13188 15204
rect 13132 15150 13134 15202
rect 13134 15150 13186 15202
rect 13186 15150 13188 15202
rect 13132 15148 13188 15150
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 14140 16098 14196 16100
rect 14140 16046 14142 16098
rect 14142 16046 14194 16098
rect 14194 16046 14196 16098
rect 14140 16044 14196 16046
rect 14476 16716 14532 16772
rect 14812 17164 14868 17220
rect 14812 16156 14868 16212
rect 14700 16098 14756 16100
rect 14700 16046 14702 16098
rect 14702 16046 14754 16098
rect 14754 16046 14756 16098
rect 14700 16044 14756 16046
rect 14364 15372 14420 15428
rect 13916 15314 13972 15316
rect 13916 15262 13918 15314
rect 13918 15262 13970 15314
rect 13970 15262 13972 15314
rect 13916 15260 13972 15262
rect 14252 15202 14308 15204
rect 14252 15150 14254 15202
rect 14254 15150 14306 15202
rect 14306 15150 14308 15202
rect 14252 15148 14308 15150
rect 14364 15090 14420 15092
rect 14364 15038 14366 15090
rect 14366 15038 14418 15090
rect 14418 15038 14420 15090
rect 14364 15036 14420 15038
rect 16828 21810 16884 21812
rect 16828 21758 16830 21810
rect 16830 21758 16882 21810
rect 16882 21758 16884 21810
rect 16828 21756 16884 21758
rect 16156 21586 16212 21588
rect 16156 21534 16158 21586
rect 16158 21534 16210 21586
rect 16210 21534 16212 21586
rect 16156 21532 16212 21534
rect 17052 21308 17108 21364
rect 16828 20130 16884 20132
rect 16828 20078 16830 20130
rect 16830 20078 16882 20130
rect 16882 20078 16884 20130
rect 16828 20076 16884 20078
rect 16604 20018 16660 20020
rect 16604 19966 16606 20018
rect 16606 19966 16658 20018
rect 16658 19966 16660 20018
rect 16604 19964 16660 19966
rect 15708 19404 15764 19460
rect 15596 18844 15652 18900
rect 18620 23884 18676 23940
rect 18396 23660 18452 23716
rect 17948 22988 18004 23044
rect 18060 22258 18116 22260
rect 18060 22206 18062 22258
rect 18062 22206 18114 22258
rect 18114 22206 18116 22258
rect 18060 22204 18116 22206
rect 18172 22092 18228 22148
rect 17612 21308 17668 21364
rect 17612 20018 17668 20020
rect 17612 19966 17614 20018
rect 17614 19966 17666 20018
rect 17666 19966 17668 20018
rect 17612 19964 17668 19966
rect 15932 19234 15988 19236
rect 15932 19182 15934 19234
rect 15934 19182 15986 19234
rect 15986 19182 15988 19234
rect 15932 19180 15988 19182
rect 15820 19068 15876 19124
rect 15372 17948 15428 18004
rect 16940 19068 16996 19124
rect 15036 17276 15092 17332
rect 16604 18396 16660 18452
rect 15708 18172 15764 18228
rect 15484 17388 15540 17444
rect 15372 16994 15428 16996
rect 15372 16942 15374 16994
rect 15374 16942 15426 16994
rect 15426 16942 15428 16994
rect 15372 16940 15428 16942
rect 15260 16770 15316 16772
rect 15260 16718 15262 16770
rect 15262 16718 15314 16770
rect 15314 16718 15316 16770
rect 15260 16716 15316 16718
rect 15596 17276 15652 17332
rect 15596 16994 15652 16996
rect 15596 16942 15598 16994
rect 15598 16942 15650 16994
rect 15650 16942 15652 16994
rect 15596 16940 15652 16942
rect 16492 17948 16548 18004
rect 16268 17836 16324 17892
rect 16828 17948 16884 18004
rect 16492 17666 16548 17668
rect 16492 17614 16494 17666
rect 16494 17614 16546 17666
rect 16546 17614 16548 17666
rect 16492 17612 16548 17614
rect 15596 16716 15652 16772
rect 15260 16044 15316 16100
rect 15148 15260 15204 15316
rect 15036 15036 15092 15092
rect 17164 17666 17220 17668
rect 17164 17614 17166 17666
rect 17166 17614 17218 17666
rect 17218 17614 17220 17666
rect 17164 17612 17220 17614
rect 17612 18396 17668 18452
rect 17500 17052 17556 17108
rect 17836 21698 17892 21700
rect 17836 21646 17838 21698
rect 17838 21646 17890 21698
rect 17890 21646 17892 21698
rect 17836 21644 17892 21646
rect 18284 21756 18340 21812
rect 17836 20076 17892 20132
rect 17948 21586 18004 21588
rect 17948 21534 17950 21586
rect 17950 21534 18002 21586
rect 18002 21534 18004 21586
rect 17948 21532 18004 21534
rect 18508 21756 18564 21812
rect 19180 25004 19236 25060
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19628 24892 19684 24948
rect 20300 24668 20356 24724
rect 19180 23884 19236 23940
rect 18732 23772 18788 23828
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 18732 23100 18788 23156
rect 23548 25506 23604 25508
rect 23548 25454 23550 25506
rect 23550 25454 23602 25506
rect 23602 25454 23604 25506
rect 23548 25452 23604 25454
rect 21196 24668 21252 24724
rect 21644 25228 21700 25284
rect 21532 23884 21588 23940
rect 19516 23042 19572 23044
rect 19516 22990 19518 23042
rect 19518 22990 19570 23042
rect 19570 22990 19572 23042
rect 19516 22988 19572 22990
rect 18844 22258 18900 22260
rect 18844 22206 18846 22258
rect 18846 22206 18898 22258
rect 18898 22206 18900 22258
rect 18844 22204 18900 22206
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19628 21756 19684 21812
rect 18844 21586 18900 21588
rect 18844 21534 18846 21586
rect 18846 21534 18898 21586
rect 18898 21534 18900 21586
rect 18844 21532 18900 21534
rect 20188 21756 20244 21812
rect 19516 21362 19572 21364
rect 19516 21310 19518 21362
rect 19518 21310 19570 21362
rect 19570 21310 19572 21362
rect 19516 21308 19572 21310
rect 19964 20802 20020 20804
rect 19964 20750 19966 20802
rect 19966 20750 20018 20802
rect 20018 20750 20020 20802
rect 19964 20748 20020 20750
rect 20524 21532 20580 21588
rect 20748 21532 20804 21588
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 17836 19292 17892 19348
rect 18060 19068 18116 19124
rect 18508 19292 18564 19348
rect 18508 19122 18564 19124
rect 18508 19070 18510 19122
rect 18510 19070 18562 19122
rect 18562 19070 18564 19122
rect 18508 19068 18564 19070
rect 18508 18844 18564 18900
rect 17724 16940 17780 16996
rect 16492 16268 16548 16324
rect 15708 16210 15764 16212
rect 15708 16158 15710 16210
rect 15710 16158 15762 16210
rect 15762 16158 15764 16210
rect 15708 16156 15764 16158
rect 15596 16098 15652 16100
rect 15596 16046 15598 16098
rect 15598 16046 15650 16098
rect 15650 16046 15652 16098
rect 15596 16044 15652 16046
rect 15484 15932 15540 15988
rect 16156 15986 16212 15988
rect 16156 15934 16158 15986
rect 16158 15934 16210 15986
rect 16210 15934 16212 15986
rect 16156 15932 16212 15934
rect 16156 15426 16212 15428
rect 16156 15374 16158 15426
rect 16158 15374 16210 15426
rect 16210 15374 16212 15426
rect 16156 15372 16212 15374
rect 18508 18172 18564 18228
rect 18844 18450 18900 18452
rect 18844 18398 18846 18450
rect 18846 18398 18898 18450
rect 18898 18398 18900 18450
rect 18844 18396 18900 18398
rect 19628 19122 19684 19124
rect 19628 19070 19630 19122
rect 19630 19070 19682 19122
rect 19682 19070 19684 19122
rect 19628 19068 19684 19070
rect 19964 18956 20020 19012
rect 20188 19122 20244 19124
rect 20188 19070 20190 19122
rect 20190 19070 20242 19122
rect 20242 19070 20244 19122
rect 20188 19068 20244 19070
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 18620 17948 18676 18004
rect 18396 16322 18452 16324
rect 18396 16270 18398 16322
rect 18398 16270 18450 16322
rect 18450 16270 18452 16322
rect 18396 16268 18452 16270
rect 18396 15372 18452 15428
rect 18508 15314 18564 15316
rect 18508 15262 18510 15314
rect 18510 15262 18562 15314
rect 18562 15262 18564 15314
rect 18508 15260 18564 15262
rect 18284 15148 18340 15204
rect 19180 17948 19236 18004
rect 19516 18172 19572 18228
rect 19628 17836 19684 17892
rect 19292 17554 19348 17556
rect 19292 17502 19294 17554
rect 19294 17502 19346 17554
rect 19346 17502 19348 17554
rect 19292 17500 19348 17502
rect 20860 21026 20916 21028
rect 20860 20974 20862 21026
rect 20862 20974 20914 21026
rect 20914 20974 20916 21026
rect 20860 20972 20916 20974
rect 20748 20690 20804 20692
rect 20748 20638 20750 20690
rect 20750 20638 20802 20690
rect 20802 20638 20804 20690
rect 20748 20636 20804 20638
rect 21420 22092 21476 22148
rect 21420 19234 21476 19236
rect 21420 19182 21422 19234
rect 21422 19182 21474 19234
rect 21474 19182 21476 19234
rect 21420 19180 21476 19182
rect 20300 18956 20356 19012
rect 20524 18674 20580 18676
rect 20524 18622 20526 18674
rect 20526 18622 20578 18674
rect 20578 18622 20580 18674
rect 20524 18620 20580 18622
rect 20412 18338 20468 18340
rect 20412 18286 20414 18338
rect 20414 18286 20466 18338
rect 20466 18286 20468 18338
rect 20412 18284 20468 18286
rect 22092 25282 22148 25284
rect 22092 25230 22094 25282
rect 22094 25230 22146 25282
rect 22146 25230 22148 25282
rect 22092 25228 22148 25230
rect 21868 24668 21924 24724
rect 21868 23884 21924 23940
rect 22876 25282 22932 25284
rect 22876 25230 22878 25282
rect 22878 25230 22930 25282
rect 22930 25230 22932 25282
rect 22876 25228 22932 25230
rect 23436 25394 23492 25396
rect 23436 25342 23438 25394
rect 23438 25342 23490 25394
rect 23490 25342 23492 25394
rect 23436 25340 23492 25342
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 24108 25340 24164 25396
rect 23660 25228 23716 25284
rect 23772 24610 23828 24612
rect 23772 24558 23774 24610
rect 23774 24558 23826 24610
rect 23826 24558 23828 24610
rect 23772 24556 23828 24558
rect 24556 24556 24612 24612
rect 25116 24556 25172 24612
rect 22988 23660 23044 23716
rect 22876 21810 22932 21812
rect 22876 21758 22878 21810
rect 22878 21758 22930 21810
rect 22930 21758 22932 21810
rect 22876 21756 22932 21758
rect 24220 22482 24276 22484
rect 24220 22430 24222 22482
rect 24222 22430 24274 22482
rect 24274 22430 24276 22482
rect 24220 22428 24276 22430
rect 24668 22146 24724 22148
rect 24668 22094 24670 22146
rect 24670 22094 24722 22146
rect 24722 22094 24724 22146
rect 24668 22092 24724 22094
rect 26236 25564 26292 25620
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 37660 25676 37716 25732
rect 27356 25618 27412 25620
rect 27356 25566 27358 25618
rect 27358 25566 27410 25618
rect 27410 25566 27412 25618
rect 27356 25564 27412 25566
rect 39900 25564 39956 25620
rect 26348 25452 26404 25508
rect 25228 23826 25284 23828
rect 25228 23774 25230 23826
rect 25230 23774 25282 23826
rect 25282 23774 25284 23826
rect 25228 23772 25284 23774
rect 25452 23436 25508 23492
rect 26348 23548 26404 23604
rect 26460 23660 26516 23716
rect 27804 24556 27860 24612
rect 27580 23884 27636 23940
rect 27356 23660 27412 23716
rect 28588 24610 28644 24612
rect 28588 24558 28590 24610
rect 28590 24558 28642 24610
rect 28642 24558 28644 24610
rect 28588 24556 28644 24558
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 28140 23660 28196 23716
rect 40012 24892 40068 24948
rect 40012 24220 40068 24276
rect 37884 23884 37940 23940
rect 37660 23660 37716 23716
rect 27244 23436 27300 23492
rect 26124 22540 26180 22596
rect 25340 22092 25396 22148
rect 24220 21868 24276 21924
rect 23436 21698 23492 21700
rect 23436 21646 23438 21698
rect 23438 21646 23490 21698
rect 23490 21646 23492 21698
rect 23436 21644 23492 21646
rect 24220 21644 24276 21700
rect 21644 21586 21700 21588
rect 21644 21534 21646 21586
rect 21646 21534 21698 21586
rect 21698 21534 21700 21586
rect 21644 21532 21700 21534
rect 21868 21474 21924 21476
rect 21868 21422 21870 21474
rect 21870 21422 21922 21474
rect 21922 21422 21924 21474
rect 21868 21420 21924 21422
rect 21868 20802 21924 20804
rect 21868 20750 21870 20802
rect 21870 20750 21922 20802
rect 21922 20750 21924 20802
rect 21868 20748 21924 20750
rect 22316 20636 22372 20692
rect 21532 18620 21588 18676
rect 20636 18172 20692 18228
rect 21308 18396 21364 18452
rect 21980 18226 22036 18228
rect 21980 18174 21982 18226
rect 21982 18174 22034 18226
rect 22034 18174 22036 18226
rect 21980 18172 22036 18174
rect 22204 18226 22260 18228
rect 22204 18174 22206 18226
rect 22206 18174 22258 18226
rect 22258 18174 22260 18226
rect 22204 18172 22260 18174
rect 21084 18060 21140 18116
rect 21420 17948 21476 18004
rect 20188 17724 20244 17780
rect 20300 17836 20356 17892
rect 20076 17500 20132 17556
rect 19852 17442 19908 17444
rect 19852 17390 19854 17442
rect 19854 17390 19906 17442
rect 19906 17390 19908 17442
rect 19852 17388 19908 17390
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19852 16994 19908 16996
rect 19852 16942 19854 16994
rect 19854 16942 19906 16994
rect 19906 16942 19908 16994
rect 19852 16940 19908 16942
rect 19292 16882 19348 16884
rect 19292 16830 19294 16882
rect 19294 16830 19346 16882
rect 19346 16830 19348 16882
rect 19292 16828 19348 16830
rect 20076 16828 20132 16884
rect 18844 15932 18900 15988
rect 19404 15820 19460 15876
rect 21756 17890 21812 17892
rect 21756 17838 21758 17890
rect 21758 17838 21810 17890
rect 21810 17838 21812 17890
rect 21756 17836 21812 17838
rect 21980 17666 22036 17668
rect 21980 17614 21982 17666
rect 21982 17614 22034 17666
rect 22034 17614 22036 17666
rect 21980 17612 22036 17614
rect 22540 18450 22596 18452
rect 22540 18398 22542 18450
rect 22542 18398 22594 18450
rect 22594 18398 22596 18450
rect 22540 18396 22596 18398
rect 23212 21084 23268 21140
rect 25228 21474 25284 21476
rect 25228 21422 25230 21474
rect 25230 21422 25282 21474
rect 25282 21422 25284 21474
rect 25228 21420 25284 21422
rect 27132 21698 27188 21700
rect 27132 21646 27134 21698
rect 27134 21646 27186 21698
rect 27186 21646 27188 21698
rect 27132 21644 27188 21646
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 37660 22370 37716 22372
rect 37660 22318 37662 22370
rect 37662 22318 37714 22370
rect 37714 22318 37716 22370
rect 37660 22316 37716 22318
rect 40012 22204 40068 22260
rect 25452 20972 25508 21028
rect 24220 19346 24276 19348
rect 24220 19294 24222 19346
rect 24222 19294 24274 19346
rect 24274 19294 24276 19346
rect 24220 19292 24276 19294
rect 24668 19234 24724 19236
rect 24668 19182 24670 19234
rect 24670 19182 24722 19234
rect 24722 19182 24724 19234
rect 24668 19180 24724 19182
rect 25340 19180 25396 19236
rect 23212 18172 23268 18228
rect 24780 18284 24836 18340
rect 23100 17836 23156 17892
rect 22428 17666 22484 17668
rect 22428 17614 22430 17666
rect 22430 17614 22482 17666
rect 22482 17614 22484 17666
rect 22428 17612 22484 17614
rect 22316 17554 22372 17556
rect 22316 17502 22318 17554
rect 22318 17502 22370 17554
rect 22370 17502 22372 17554
rect 22316 17500 22372 17502
rect 22316 16940 22372 16996
rect 22988 17500 23044 17556
rect 20188 15874 20244 15876
rect 20188 15822 20190 15874
rect 20190 15822 20242 15874
rect 20242 15822 20244 15874
rect 20188 15820 20244 15822
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19964 15314 20020 15316
rect 19964 15262 19966 15314
rect 19966 15262 20018 15314
rect 20018 15262 20020 15314
rect 19964 15260 20020 15262
rect 18956 15148 19012 15204
rect 19068 15090 19124 15092
rect 19068 15038 19070 15090
rect 19070 15038 19122 15090
rect 19122 15038 19124 15090
rect 19068 15036 19124 15038
rect 15148 14252 15204 14308
rect 15932 14252 15988 14308
rect 16716 14252 16772 14308
rect 19180 14306 19236 14308
rect 19180 14254 19182 14306
rect 19182 14254 19234 14306
rect 19234 14254 19236 14306
rect 19180 14252 19236 14254
rect 20860 15202 20916 15204
rect 20860 15150 20862 15202
rect 20862 15150 20914 15202
rect 20914 15150 20916 15202
rect 20860 15148 20916 15150
rect 25228 17554 25284 17556
rect 25228 17502 25230 17554
rect 25230 17502 25282 17554
rect 25282 17502 25284 17554
rect 25228 17500 25284 17502
rect 23996 17388 24052 17444
rect 24220 17388 24276 17444
rect 25116 16940 25172 16996
rect 24668 16882 24724 16884
rect 24668 16830 24670 16882
rect 24670 16830 24722 16882
rect 24722 16830 24724 16882
rect 24668 16828 24724 16830
rect 26796 21586 26852 21588
rect 26796 21534 26798 21586
rect 26798 21534 26850 21586
rect 26850 21534 26852 21586
rect 26796 21532 26852 21534
rect 26348 20972 26404 21028
rect 28364 21644 28420 21700
rect 27916 21586 27972 21588
rect 27916 21534 27918 21586
rect 27918 21534 27970 21586
rect 27970 21534 27972 21586
rect 27916 21532 27972 21534
rect 27692 20188 27748 20244
rect 28252 20188 28308 20244
rect 37660 21586 37716 21588
rect 37660 21534 37662 21586
rect 37662 21534 37714 21586
rect 37714 21534 37716 21586
rect 37660 21532 37716 21534
rect 40012 21532 40068 21588
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 40012 20914 40068 20916
rect 40012 20862 40014 20914
rect 40014 20862 40066 20914
rect 40066 20862 40068 20914
rect 40012 20860 40068 20862
rect 37660 20188 37716 20244
rect 40012 20076 40068 20132
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 37660 19292 37716 19348
rect 28588 18956 28644 19012
rect 26012 17724 26068 17780
rect 25900 17612 25956 17668
rect 26236 17554 26292 17556
rect 26236 17502 26238 17554
rect 26238 17502 26290 17554
rect 26290 17502 26292 17554
rect 26236 17500 26292 17502
rect 25676 17442 25732 17444
rect 25676 17390 25678 17442
rect 25678 17390 25730 17442
rect 25730 17390 25732 17442
rect 25676 17388 25732 17390
rect 25452 17052 25508 17108
rect 26796 17724 26852 17780
rect 27132 17612 27188 17668
rect 26348 17052 26404 17108
rect 26012 16994 26068 16996
rect 26012 16942 26014 16994
rect 26014 16942 26066 16994
rect 26066 16942 26068 16994
rect 26012 16940 26068 16942
rect 26460 16828 26516 16884
rect 24220 16098 24276 16100
rect 24220 16046 24222 16098
rect 24222 16046 24274 16098
rect 24274 16046 24276 16098
rect 24220 16044 24276 16046
rect 21868 15148 21924 15204
rect 29260 19010 29316 19012
rect 29260 18958 29262 19010
rect 29262 18958 29314 19010
rect 29314 18958 29316 19010
rect 29260 18956 29316 18958
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 37660 17666 37716 17668
rect 37660 17614 37662 17666
rect 37662 17614 37714 17666
rect 37714 17614 37716 17666
rect 37660 17612 37716 17614
rect 40012 17500 40068 17556
rect 28140 16828 28196 16884
rect 25228 16044 25284 16100
rect 27580 16098 27636 16100
rect 27580 16046 27582 16098
rect 27582 16046 27634 16098
rect 27634 16046 27636 16098
rect 27580 16044 27636 16046
rect 37660 16882 37716 16884
rect 37660 16830 37662 16882
rect 37662 16830 37714 16882
rect 37714 16830 37716 16882
rect 37660 16828 37716 16830
rect 40012 16828 40068 16884
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 28364 16044 28420 16100
rect 20748 14476 20804 14532
rect 21756 14476 21812 14532
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 18956 13746 19012 13748
rect 18956 13694 18958 13746
rect 18958 13694 19010 13746
rect 19010 13694 19012 13746
rect 18956 13692 19012 13694
rect 15036 13468 15092 13524
rect 22428 14530 22484 14532
rect 22428 14478 22430 14530
rect 22430 14478 22482 14530
rect 22482 14478 22484 14530
rect 22428 14476 22484 14478
rect 16268 13468 16324 13524
rect 16940 13468 16996 13524
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 20860 5180 20916 5236
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 16156 3388 16212 3444
rect 18508 3442 18564 3444
rect 18508 3390 18510 3442
rect 18510 3390 18562 3442
rect 18562 3390 18564 3442
rect 18508 3388 18564 3390
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 22204 13746 22260 13748
rect 22204 13694 22206 13746
rect 22206 13694 22258 13746
rect 22258 13694 22260 13746
rect 22204 13692 22260 13694
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 23660 13692 23716 13748
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 40236 5404 40292 5460
rect 22316 5234 22372 5236
rect 22316 5182 22318 5234
rect 22318 5182 22370 5234
rect 22370 5182 22372 5234
rect 22316 5180 22372 5182
rect 21532 4060 21588 4116
rect 22764 4114 22820 4116
rect 22764 4062 22766 4114
rect 22766 4062 22818 4114
rect 22818 4062 22820 4114
rect 22764 4060 22820 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 23538 38220 23548 38276
rect 23604 38220 25564 38276
rect 25620 38220 25630 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 19506 37436 19516 37492
rect 19572 37436 20748 37492
rect 20804 37436 20814 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 4274 27020 4284 27076
rect 4340 27020 14028 27076
rect 14084 27020 14094 27076
rect 18834 26796 18844 26852
rect 18900 26796 20188 26852
rect 20244 26796 20254 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 0 26292 800 26320
rect 0 26236 1932 26292
rect 1988 26236 1998 26292
rect 4274 26236 4284 26292
rect 4340 26236 14700 26292
rect 14756 26236 14766 26292
rect 0 26208 800 26236
rect 18162 26124 18172 26180
rect 18228 26124 19068 26180
rect 19124 26124 19134 26180
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 31892 25676 37660 25732
rect 37716 25676 37726 25732
rect 0 25620 800 25648
rect 31892 25620 31948 25676
rect 41200 25620 42000 25648
rect 0 25564 1932 25620
rect 1988 25564 1998 25620
rect 26226 25564 26236 25620
rect 26292 25564 27356 25620
rect 27412 25564 31948 25620
rect 39890 25564 39900 25620
rect 39956 25564 42000 25620
rect 0 25536 800 25564
rect 41200 25536 42000 25564
rect 15698 25452 15708 25508
rect 15764 25452 16940 25508
rect 16996 25452 17006 25508
rect 23538 25452 23548 25508
rect 23604 25452 26348 25508
rect 26404 25452 26414 25508
rect 23426 25340 23436 25396
rect 23492 25340 24108 25396
rect 24164 25340 24174 25396
rect 18946 25228 18956 25284
rect 19012 25228 21644 25284
rect 21700 25228 22092 25284
rect 22148 25228 22158 25284
rect 22866 25228 22876 25284
rect 22932 25228 23660 25284
rect 23716 25228 23726 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 16930 25004 16940 25060
rect 16996 25004 19180 25060
rect 19236 25004 19246 25060
rect 0 24948 800 24976
rect 41200 24948 42000 24976
rect 0 24892 2044 24948
rect 2100 24892 2110 24948
rect 4274 24892 4284 24948
rect 4340 24892 11564 24948
rect 11620 24892 14252 24948
rect 14308 24892 14924 24948
rect 14980 24892 14990 24948
rect 16482 24892 16492 24948
rect 16548 24892 17724 24948
rect 17780 24892 17790 24948
rect 18722 24892 18732 24948
rect 18788 24892 19628 24948
rect 19684 24892 19694 24948
rect 40002 24892 40012 24948
rect 40068 24892 42000 24948
rect 0 24864 800 24892
rect 41200 24864 42000 24892
rect 17602 24780 17612 24836
rect 17668 24780 21924 24836
rect 21868 24724 21924 24780
rect 4274 24668 4284 24724
rect 4340 24668 14476 24724
rect 14532 24668 14542 24724
rect 20290 24668 20300 24724
rect 20356 24668 21196 24724
rect 21252 24668 21262 24724
rect 21858 24668 21868 24724
rect 21924 24668 21934 24724
rect 23762 24556 23772 24612
rect 23828 24556 24556 24612
rect 24612 24556 25116 24612
rect 25172 24556 27804 24612
rect 27860 24556 28588 24612
rect 28644 24556 28654 24612
rect 1922 24444 1932 24500
rect 1988 24444 1998 24500
rect 0 24276 800 24304
rect 1932 24276 1988 24444
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 41200 24276 42000 24304
rect 0 24220 1988 24276
rect 40002 24220 40012 24276
rect 40068 24220 42000 24276
rect 0 24192 800 24220
rect 41200 24192 42000 24220
rect 18610 23884 18620 23940
rect 18676 23884 19180 23940
rect 19236 23884 20188 23940
rect 21522 23884 21532 23940
rect 21588 23884 21868 23940
rect 21924 23884 21934 23940
rect 27570 23884 27580 23940
rect 27636 23884 37884 23940
rect 37940 23884 37950 23940
rect 20132 23828 20188 23884
rect 12898 23772 12908 23828
rect 12964 23772 14140 23828
rect 14196 23772 14206 23828
rect 14466 23772 14476 23828
rect 14532 23772 15036 23828
rect 15092 23772 17388 23828
rect 17444 23772 18732 23828
rect 18788 23772 18798 23828
rect 20132 23772 25228 23828
rect 25284 23772 25294 23828
rect 17714 23660 17724 23716
rect 17780 23660 18396 23716
rect 18452 23660 22988 23716
rect 23044 23660 23054 23716
rect 26450 23660 26460 23716
rect 26516 23660 27356 23716
rect 27412 23660 28140 23716
rect 28196 23660 37660 23716
rect 37716 23660 37726 23716
rect 0 23604 800 23632
rect 0 23548 4172 23604
rect 4228 23548 4238 23604
rect 26338 23548 26348 23604
rect 26404 23548 26414 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 26348 23492 26404 23548
rect 25442 23436 25452 23492
rect 25508 23436 27244 23492
rect 27300 23436 27310 23492
rect 4274 23100 4284 23156
rect 4340 23100 17388 23156
rect 17444 23100 18732 23156
rect 18788 23100 18798 23156
rect 17938 22988 17948 23044
rect 18004 22988 19516 23044
rect 19572 22988 19582 23044
rect 0 22932 800 22960
rect 0 22876 1932 22932
rect 1988 22876 1998 22932
rect 0 22848 800 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 14130 22540 14140 22596
rect 14196 22540 16716 22596
rect 16772 22540 26124 22596
rect 26180 22540 26190 22596
rect 24210 22428 24220 22484
rect 24276 22428 31948 22484
rect 31892 22372 31948 22428
rect 31892 22316 37660 22372
rect 37716 22316 37726 22372
rect 41200 22260 42000 22288
rect 18050 22204 18060 22260
rect 18116 22204 18844 22260
rect 18900 22204 18910 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 41200 22176 42000 22204
rect 12002 22092 12012 22148
rect 12068 22092 16828 22148
rect 16884 22092 16894 22148
rect 18162 22092 18172 22148
rect 18228 22092 21420 22148
rect 21476 22092 21486 22148
rect 24658 22092 24668 22148
rect 24724 22092 25340 22148
rect 25396 22092 25406 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 24210 21868 24220 21924
rect 24276 21868 24286 21924
rect 24220 21812 24276 21868
rect 16818 21756 16828 21812
rect 16884 21756 18284 21812
rect 18340 21756 18508 21812
rect 18564 21756 19628 21812
rect 19684 21756 20188 21812
rect 20244 21756 20254 21812
rect 22866 21756 22876 21812
rect 22932 21756 24276 21812
rect 17826 21644 17836 21700
rect 17892 21644 18564 21700
rect 23426 21644 23436 21700
rect 23492 21644 24220 21700
rect 24276 21644 24286 21700
rect 27122 21644 27132 21700
rect 27188 21644 28364 21700
rect 28420 21644 31948 21700
rect 18508 21588 18564 21644
rect 31892 21588 31948 21644
rect 41200 21588 42000 21616
rect 15250 21532 15260 21588
rect 15316 21532 16156 21588
rect 16212 21532 17948 21588
rect 18004 21532 18014 21588
rect 18508 21532 18844 21588
rect 18900 21532 20524 21588
rect 20580 21532 20590 21588
rect 20738 21532 20748 21588
rect 20804 21532 21644 21588
rect 21700 21532 21710 21588
rect 26786 21532 26796 21588
rect 26852 21532 27916 21588
rect 27972 21532 27982 21588
rect 31892 21532 37660 21588
rect 37716 21532 37726 21588
rect 40002 21532 40012 21588
rect 40068 21532 42000 21588
rect 41200 21504 42000 21532
rect 21858 21420 21868 21476
rect 21924 21420 25228 21476
rect 25284 21420 25294 21476
rect 17042 21308 17052 21364
rect 17108 21308 17612 21364
rect 17668 21308 19516 21364
rect 19572 21308 19582 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 23212 21140 23268 21420
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 23202 21084 23212 21140
rect 23268 21084 23278 21140
rect 20850 20972 20860 21028
rect 20916 20972 25452 21028
rect 25508 20972 26348 21028
rect 26404 20972 26414 21028
rect 41200 20916 42000 20944
rect 40002 20860 40012 20916
rect 40068 20860 42000 20916
rect 41200 20832 42000 20860
rect 14130 20748 14140 20804
rect 14196 20748 15596 20804
rect 15652 20748 15662 20804
rect 19954 20748 19964 20804
rect 20020 20748 21868 20804
rect 21924 20748 21934 20804
rect 14466 20636 14476 20692
rect 14532 20636 15372 20692
rect 15428 20636 15438 20692
rect 20738 20636 20748 20692
rect 20804 20636 22316 20692
rect 22372 20636 22382 20692
rect 11890 20524 11900 20580
rect 11956 20524 14252 20580
rect 14308 20524 14318 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 41200 20244 42000 20272
rect 27682 20188 27692 20244
rect 27748 20188 28252 20244
rect 28308 20188 37660 20244
rect 37716 20188 37726 20244
rect 40012 20188 42000 20244
rect 40012 20132 40068 20188
rect 41200 20160 42000 20188
rect 11330 20076 11340 20132
rect 11396 20076 14140 20132
rect 14196 20076 14206 20132
rect 16818 20076 16828 20132
rect 16884 20076 17836 20132
rect 17892 20076 17902 20132
rect 40002 20076 40012 20132
rect 40068 20076 40078 20132
rect 14802 19964 14812 20020
rect 14868 19964 15484 20020
rect 15540 19964 16604 20020
rect 16660 19964 17612 20020
rect 17668 19964 17678 20020
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 13682 19516 13692 19572
rect 13748 19516 14588 19572
rect 14644 19516 15372 19572
rect 15428 19516 15438 19572
rect 14018 19404 14028 19460
rect 14084 19404 14924 19460
rect 14980 19404 15708 19460
rect 15764 19404 15774 19460
rect 4162 19292 4172 19348
rect 4228 19292 17836 19348
rect 17892 19292 18508 19348
rect 18564 19292 18574 19348
rect 24210 19292 24220 19348
rect 24276 19292 37660 19348
rect 37716 19292 37726 19348
rect 14690 19180 14700 19236
rect 14756 19180 15932 19236
rect 15988 19180 15998 19236
rect 21410 19180 21420 19236
rect 21476 19180 24668 19236
rect 24724 19180 25340 19236
rect 25396 19180 25406 19236
rect 15810 19068 15820 19124
rect 15876 19068 16940 19124
rect 16996 19068 17006 19124
rect 18050 19068 18060 19124
rect 18116 19068 18508 19124
rect 18564 19068 18574 19124
rect 19618 19068 19628 19124
rect 19684 19068 20188 19124
rect 20244 19068 20254 19124
rect 18508 18956 19964 19012
rect 20020 18956 20300 19012
rect 20356 18956 20366 19012
rect 28578 18956 28588 19012
rect 28644 18956 29260 19012
rect 29316 18956 29326 19012
rect 18508 18900 18564 18956
rect 15586 18844 15596 18900
rect 15652 18844 18508 18900
rect 18564 18844 18574 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 14018 18620 14028 18676
rect 14084 18620 14812 18676
rect 14868 18620 14878 18676
rect 20514 18620 20524 18676
rect 20580 18620 21532 18676
rect 21588 18620 21598 18676
rect 16594 18396 16604 18452
rect 16660 18396 17612 18452
rect 17668 18396 18844 18452
rect 18900 18396 18910 18452
rect 21298 18396 21308 18452
rect 21364 18396 22540 18452
rect 22596 18396 22606 18452
rect 20402 18284 20412 18340
rect 20468 18284 24780 18340
rect 24836 18284 24846 18340
rect 12786 18172 12796 18228
rect 12852 18172 14252 18228
rect 14308 18172 15708 18228
rect 15764 18172 18508 18228
rect 18564 18172 19516 18228
rect 19572 18172 19582 18228
rect 20626 18172 20636 18228
rect 20692 18172 21980 18228
rect 22036 18172 22046 18228
rect 22194 18172 22204 18228
rect 22260 18172 23212 18228
rect 23268 18172 23278 18228
rect 22204 18116 22260 18172
rect 21074 18060 21084 18116
rect 21140 18060 22260 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 15362 17948 15372 18004
rect 15428 17948 16492 18004
rect 16548 17948 16558 18004
rect 16818 17948 16828 18004
rect 16884 17948 18620 18004
rect 18676 17948 19180 18004
rect 19236 17948 21420 18004
rect 21476 17948 21486 18004
rect 13906 17836 13916 17892
rect 13972 17836 14812 17892
rect 14868 17836 16268 17892
rect 16324 17836 16334 17892
rect 19618 17836 19628 17892
rect 19684 17836 20300 17892
rect 20356 17836 21756 17892
rect 21812 17836 23100 17892
rect 23156 17836 23166 17892
rect 20178 17724 20188 17780
rect 20244 17724 26012 17780
rect 26068 17724 26796 17780
rect 26852 17724 26862 17780
rect 4274 17612 4284 17668
rect 4340 17612 10668 17668
rect 10724 17612 10734 17668
rect 16482 17612 16492 17668
rect 16548 17612 17164 17668
rect 17220 17612 17230 17668
rect 21970 17612 21980 17668
rect 22036 17612 22428 17668
rect 22484 17612 22494 17668
rect 25890 17612 25900 17668
rect 25956 17612 27132 17668
rect 27188 17612 37660 17668
rect 37716 17612 37726 17668
rect 41200 17556 42000 17584
rect 19282 17500 19292 17556
rect 19348 17500 20076 17556
rect 20132 17500 20142 17556
rect 22306 17500 22316 17556
rect 22372 17500 22988 17556
rect 23044 17500 23054 17556
rect 25218 17500 25228 17556
rect 25284 17500 26236 17556
rect 26292 17500 26302 17556
rect 40002 17500 40012 17556
rect 40068 17500 42000 17556
rect 41200 17472 42000 17500
rect 14354 17388 14364 17444
rect 14420 17388 15484 17444
rect 15540 17388 15550 17444
rect 19842 17388 19852 17444
rect 19908 17388 23996 17444
rect 24052 17388 24062 17444
rect 24210 17388 24220 17444
rect 24276 17388 25676 17444
rect 25732 17388 25742 17444
rect 15026 17276 15036 17332
rect 15092 17276 15596 17332
rect 15652 17276 15662 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 12786 17164 12796 17220
rect 12852 17164 14812 17220
rect 14868 17164 14878 17220
rect 17490 17052 17500 17108
rect 17556 17052 25452 17108
rect 25508 17052 26348 17108
rect 26404 17052 26414 17108
rect 24444 16996 24500 17052
rect 10658 16940 10668 16996
rect 10724 16940 15372 16996
rect 15428 16940 15438 16996
rect 15586 16940 15596 16996
rect 15652 16940 17724 16996
rect 17780 16940 19572 16996
rect 19842 16940 19852 16996
rect 19908 16940 22316 16996
rect 22372 16940 22382 16996
rect 24444 16940 24724 16996
rect 25106 16940 25116 16996
rect 25172 16940 26012 16996
rect 26068 16940 26078 16996
rect 0 16884 800 16912
rect 19516 16884 19572 16940
rect 24668 16884 24724 16940
rect 41200 16884 42000 16912
rect 0 16828 1932 16884
rect 1988 16828 1998 16884
rect 15596 16828 19292 16884
rect 19348 16828 19358 16884
rect 19516 16828 20076 16884
rect 20132 16828 20142 16884
rect 24658 16828 24668 16884
rect 24724 16828 24734 16884
rect 26450 16828 26460 16884
rect 26516 16828 28140 16884
rect 28196 16828 37660 16884
rect 37716 16828 37726 16884
rect 40002 16828 40012 16884
rect 40068 16828 42000 16884
rect 0 16800 800 16828
rect 15596 16772 15652 16828
rect 41200 16800 42000 16828
rect 14466 16716 14476 16772
rect 14532 16716 15260 16772
rect 15316 16716 15326 16772
rect 15586 16716 15596 16772
rect 15652 16716 15662 16772
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 16482 16268 16492 16324
rect 16548 16268 18396 16324
rect 18452 16268 18462 16324
rect 14802 16156 14812 16212
rect 14868 16156 15708 16212
rect 15764 16156 15774 16212
rect 4274 16044 4284 16100
rect 4340 16044 11004 16100
rect 11060 16044 14140 16100
rect 14196 16044 14206 16100
rect 14690 16044 14700 16100
rect 14756 16044 15260 16100
rect 15316 16044 15596 16100
rect 15652 16044 15662 16100
rect 24210 16044 24220 16100
rect 24276 16044 25228 16100
rect 25284 16044 27580 16100
rect 27636 16044 28364 16100
rect 28420 16044 28430 16100
rect 15474 15932 15484 15988
rect 15540 15932 16156 15988
rect 16212 15932 18844 15988
rect 18900 15932 18910 15988
rect 19394 15820 19404 15876
rect 19460 15820 20188 15876
rect 20244 15820 20254 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 0 15540 800 15568
rect 0 15484 1932 15540
rect 1988 15484 1998 15540
rect 0 15456 800 15484
rect 14354 15372 14364 15428
rect 14420 15372 16156 15428
rect 16212 15372 18396 15428
rect 18452 15372 18462 15428
rect 13458 15260 13468 15316
rect 13524 15260 13916 15316
rect 13972 15260 15148 15316
rect 15204 15260 15214 15316
rect 18498 15260 18508 15316
rect 18564 15260 19964 15316
rect 20020 15260 20030 15316
rect 13122 15148 13132 15204
rect 13188 15148 14252 15204
rect 14308 15148 14318 15204
rect 18274 15148 18284 15204
rect 18340 15148 18956 15204
rect 19012 15148 20860 15204
rect 20916 15148 21868 15204
rect 21924 15148 21934 15204
rect 14354 15036 14364 15092
rect 14420 15036 15036 15092
rect 15092 15036 19068 15092
rect 19124 15036 19134 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 20738 14476 20748 14532
rect 20804 14476 21756 14532
rect 21812 14476 22428 14532
rect 22484 14476 22494 14532
rect 15138 14252 15148 14308
rect 15204 14252 15932 14308
rect 15988 14252 16716 14308
rect 16772 14252 19180 14308
rect 19236 14252 19246 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 18946 13692 18956 13748
rect 19012 13692 22204 13748
rect 22260 13692 23660 13748
rect 23716 13692 23726 13748
rect 15026 13468 15036 13524
rect 15092 13468 16268 13524
rect 16324 13468 16940 13524
rect 16996 13468 17006 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 41200 5460 42000 5488
rect 40226 5404 40236 5460
rect 40292 5404 42000 5460
rect 41200 5376 42000 5404
rect 20850 5180 20860 5236
rect 20916 5180 22316 5236
rect 22372 5180 22382 5236
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 21522 4060 21532 4116
rect 21588 4060 22764 4116
rect 22820 4060 22830 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 16146 3388 16156 3444
rect 16212 3388 18508 3444
rect 18564 3388 18574 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _084_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21616 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _085_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19824 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _086_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22176 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _087_
timestamp 1698175906
transform 1 0 15792 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _088_
timestamp 1698175906
transform 1 0 19152 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _089_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15008 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _090_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16352 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _091_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _092_
timestamp 1698175906
transform 1 0 14560 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _093_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _094_
timestamp 1698175906
transform -1 0 17920 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _095_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19712 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _096_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18816 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _097_
timestamp 1698175906
transform 1 0 26656 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _098_
timestamp 1698175906
transform -1 0 27440 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _099_
timestamp 1698175906
transform 1 0 22960 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _100_
timestamp 1698175906
transform -1 0 22624 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _101_
timestamp 1698175906
transform 1 0 16352 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _102_
timestamp 1698175906
transform 1 0 16352 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _104_
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14784 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19152 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _107_
timestamp 1698175906
transform -1 0 18032 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _108_
timestamp 1698175906
transform 1 0 16576 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25760 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1698175906
transform 1 0 18592 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _111_
timestamp 1698175906
transform -1 0 19824 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _112_
timestamp 1698175906
transform -1 0 21728 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _113_
timestamp 1698175906
transform -1 0 18928 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _114_
timestamp 1698175906
transform 1 0 17472 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform 1 0 22848 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _116_
timestamp 1698175906
transform -1 0 23744 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _117_
timestamp 1698175906
transform 1 0 21728 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _118_
timestamp 1698175906
transform -1 0 18704 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _119_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16576 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _120_
timestamp 1698175906
transform 1 0 15232 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform -1 0 16800 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _122_
timestamp 1698175906
transform -1 0 15120 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _123_
timestamp 1698175906
transform 1 0 15120 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _124_
timestamp 1698175906
transform -1 0 14560 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _125_
timestamp 1698175906
transform 1 0 16576 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19152 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _127_
timestamp 1698175906
transform -1 0 14672 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _128_
timestamp 1698175906
transform -1 0 13104 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _129_
timestamp 1698175906
transform -1 0 15232 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _130_
timestamp 1698175906
transform -1 0 14112 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _131_
timestamp 1698175906
transform 1 0 17360 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _132_
timestamp 1698175906
transform 1 0 19936 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _133_
timestamp 1698175906
transform 1 0 13888 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _134_
timestamp 1698175906
transform 1 0 19264 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _135_
timestamp 1698175906
transform -1 0 17024 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _136_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14560 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19600 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19824 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _139_
timestamp 1698175906
transform -1 0 23184 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _140_
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _141_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14112 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _142_
timestamp 1698175906
transform -1 0 14896 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _143_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15008 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _144_
timestamp 1698175906
transform -1 0 26544 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _145_
timestamp 1698175906
transform 1 0 25088 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _146_
timestamp 1698175906
transform -1 0 15680 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _147_
timestamp 1698175906
transform -1 0 14784 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _148_
timestamp 1698175906
transform 1 0 15456 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _149_
timestamp 1698175906
transform -1 0 16016 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _150_
timestamp 1698175906
transform -1 0 16016 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _151_
timestamp 1698175906
transform 1 0 14336 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _152_
timestamp 1698175906
transform -1 0 19152 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _153_
timestamp 1698175906
transform -1 0 18256 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _154_
timestamp 1698175906
transform 1 0 23184 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _155_
timestamp 1698175906
transform -1 0 22960 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _156_
timestamp 1698175906
transform -1 0 23184 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _157_
timestamp 1698175906
transform -1 0 22624 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698175906
transform 1 0 27440 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _159_
timestamp 1698175906
transform -1 0 26880 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform 1 0 26096 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _161_
timestamp 1698175906
transform 1 0 25984 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _162_
timestamp 1698175906
transform -1 0 26208 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _163_
timestamp 1698175906
transform 1 0 19152 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _164_
timestamp 1698175906
transform 1 0 23968 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _165_
timestamp 1698175906
transform -1 0 26768 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _166_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20720 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _167_
timestamp 1698175906
transform 1 0 24752 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _168_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _169_
timestamp 1698175906
transform 1 0 25312 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _170_
timestamp 1698175906
transform 1 0 15568 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _171_
timestamp 1698175906
transform 1 0 21056 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _172_
timestamp 1698175906
transform -1 0 23968 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _173_
timestamp 1698175906
transform 1 0 15680 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _174_
timestamp 1698175906
transform 1 0 10976 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _175_
timestamp 1698175906
transform 1 0 11088 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _176_
timestamp 1698175906
transform 1 0 11424 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _177_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14784 0 -1 23520
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _178_
timestamp 1698175906
transform 1 0 18704 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _179_
timestamp 1698175906
transform 1 0 19600 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _180_
timestamp 1698175906
transform -1 0 14112 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _181_
timestamp 1698175906
transform 1 0 24304 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _182_
timestamp 1698175906
transform 1 0 13216 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _183_
timestamp 1698175906
transform -1 0 13776 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _184_
timestamp 1698175906
transform -1 0 20496 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _185_
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _186_
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _187_
timestamp 1698175906
transform 1 0 25200 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _188_
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _189_
timestamp 1698175906
transform 1 0 24080 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _190_
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _193_
timestamp 1698175906
transform -1 0 14560 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _194_
timestamp 1698175906
transform 1 0 21392 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _195_
timestamp 1698175906
transform 1 0 27104 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _196_
timestamp 1698175906
transform -1 0 22736 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _197_
timestamp 1698175906
transform -1 0 15232 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__168__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__CLK
timestamp 1698175906
transform 1 0 29232 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__170__CLK
timestamp 1698175906
transform 1 0 19152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__CLK
timestamp 1698175906
transform -1 0 24752 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__CLK
timestamp 1698175906
transform 1 0 24192 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__173__CLK
timestamp 1698175906
transform 1 0 19152 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__CLK
timestamp 1698175906
transform 1 0 14448 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__CLK
timestamp 1698175906
transform 1 0 14336 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__CLK
timestamp 1698175906
transform 1 0 15456 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__CLK
timestamp 1698175906
transform 1 0 15008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__CLK
timestamp 1698175906
transform 1 0 22176 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__CLK
timestamp 1698175906
transform 1 0 23744 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__CLK
timestamp 1698175906
transform 1 0 15120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__CLK
timestamp 1698175906
transform 1 0 27776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__CLK
timestamp 1698175906
transform 1 0 16688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__CLK
timestamp 1698175906
transform 1 0 14000 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__CLK
timestamp 1698175906
transform 1 0 20720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__CLK
timestamp 1698175906
transform 1 0 24640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__CLK
timestamp 1698175906
transform 1 0 24640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__CLK
timestamp 1698175906
transform 1 0 28672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__CLK
timestamp 1698175906
transform 1 0 28560 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__CLK
timestamp 1698175906
transform 1 0 27552 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__CLK
timestamp 1698175906
transform 1 0 28560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 18032 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18368 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 20160 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 21728 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_104 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_120 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14784 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_124 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_126 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15456 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_131
timestamp 1698175906
transform 1 0 16016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_135
timestamp 1698175906
transform 1 0 16464 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_164
timestamp 1698175906
transform 1 0 19712 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_168
timestamp 1698175906
transform 1 0 20160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_174
timestamp 1698175906
transform 1 0 20832 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_178
timestamp 1698175906
transform 1 0 21280 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_180
timestamp 1698175906
transform 1 0 21504 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_203
timestamp 1698175906
transform 1 0 24080 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_235 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27664 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_243
timestamp 1698175906
transform 1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_314
timestamp 1698175906
transform 1 0 36512 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_330
timestamp 1698175906
transform 1 0 38304 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_338
timestamp 1698175906
transform 1 0 39200 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_342
timestamp 1698175906
transform 1 0 39648 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_344
timestamp 1698175906
transform 1 0 39872 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_104
timestamp 1698175906
transform 1 0 12992 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_135
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698175906
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_150
timestamp 1698175906
transform 1 0 18144 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_154
timestamp 1698175906
transform 1 0 18592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_184
timestamp 1698175906
transform 1 0 21952 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_188
timestamp 1698175906
transform 1 0 22400 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_204
timestamp 1698175906
transform 1 0 24192 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698175906
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_111
timestamp 1698175906
transform 1 0 13776 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_113
timestamp 1698175906
transform 1 0 14000 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_157
timestamp 1698175906
transform 1 0 18928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_161
timestamp 1698175906
transform 1 0 19376 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_169
timestamp 1698175906
transform 1 0 20272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698175906
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_191
timestamp 1698175906
transform 1 0 22736 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_223
timestamp 1698175906
transform 1 0 26320 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_239
timestamp 1698175906
transform 1 0 28112 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698175906
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_80
timestamp 1698175906
transform 1 0 10304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_84
timestamp 1698175906
transform 1 0 10752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_122
timestamp 1698175906
transform 1 0 15008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_144
timestamp 1698175906
transform 1 0 17472 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_171
timestamp 1698175906
transform 1 0 20496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_202
timestamp 1698175906
transform 1 0 23968 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698175906
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_28
timestamp 1698175906
transform 1 0 4480 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698175906
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_111
timestamp 1698175906
transform 1 0 13776 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_121
timestamp 1698175906
transform 1 0 14896 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_125
timestamp 1698175906
transform 1 0 15344 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_134
timestamp 1698175906
transform 1 0 16352 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_150
timestamp 1698175906
transform 1 0 18144 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_159
timestamp 1698175906
transform 1 0 19152 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_163
timestamp 1698175906
transform 1 0 19600 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_165
timestamp 1698175906
transform 1 0 19824 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_193
timestamp 1698175906
transform 1 0 22960 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_201
timestamp 1698175906
transform 1 0 23856 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_232
timestamp 1698175906
transform 1 0 27328 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_236
timestamp 1698175906
transform 1 0 27776 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_80
timestamp 1698175906
transform 1 0 10304 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_111
timestamp 1698175906
transform 1 0 13776 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_115
timestamp 1698175906
transform 1 0 14224 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_131
timestamp 1698175906
transform 1 0 16016 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_158
timestamp 1698175906
transform 1 0 19040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_167
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_175
timestamp 1698175906
transform 1 0 20944 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_179
timestamp 1698175906
transform 1 0 21392 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_187
timestamp 1698175906
transform 1 0 22288 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_195
timestamp 1698175906
transform 1 0 23184 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_199
timestamp 1698175906
transform 1 0 23632 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_201
timestamp 1698175906
transform 1 0 23856 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_241
timestamp 1698175906
transform 1 0 28336 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_245
timestamp 1698175906
transform 1 0 28784 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698175906
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 36512 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 37408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_111
timestamp 1698175906
transform 1 0 13776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_113
timestamp 1698175906
transform 1 0 14000 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_131
timestamp 1698175906
transform 1 0 16016 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_138
timestamp 1698175906
transform 1 0 16800 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_149
timestamp 1698175906
transform 1 0 18032 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_157
timestamp 1698175906
transform 1 0 18928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_166
timestamp 1698175906
transform 1 0 19936 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_190
timestamp 1698175906
transform 1 0 22624 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_206
timestamp 1698175906
transform 1 0 24416 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_208
timestamp 1698175906
transform 1 0 24640 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_227
timestamp 1698175906
transform 1 0 26768 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698175906
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_104
timestamp 1698175906
transform 1 0 12992 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_133
timestamp 1698175906
transform 1 0 16240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_146
timestamp 1698175906
transform 1 0 17696 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_197
timestamp 1698175906
transform 1 0 23408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_205
timestamp 1698175906
transform 1 0 24304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_216
timestamp 1698175906
transform 1 0 25536 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_232
timestamp 1698175906
transform 1 0 27328 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_264
timestamp 1698175906
transform 1 0 30912 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 40320 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_115
timestamp 1698175906
transform 1 0 14224 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_128
timestamp 1698175906
transform 1 0 15680 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_135
timestamp 1698175906
transform 1 0 16464 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698175906
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_206
timestamp 1698175906
transform 1 0 24416 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_210
timestamp 1698175906
transform 1 0 24864 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698175906
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_251
timestamp 1698175906
transform 1 0 29456 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_80
timestamp 1698175906
transform 1 0 10304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_84
timestamp 1698175906
transform 1 0 10752 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_115
timestamp 1698175906
transform 1 0 14224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_119
timestamp 1698175906
transform 1 0 14672 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_132
timestamp 1698175906
transform 1 0 16128 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_202
timestamp 1698175906
transform 1 0 23968 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_242
timestamp 1698175906
transform 1 0 28448 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_246
timestamp 1698175906
transform 1 0 28896 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_109
timestamp 1698175906
transform 1 0 13552 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_181
timestamp 1698175906
transform 1 0 21616 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_232
timestamp 1698175906
transform 1 0 27328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_240
timestamp 1698175906
transform 1 0 28224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_80
timestamp 1698175906
transform 1 0 10304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_84
timestamp 1698175906
transform 1 0 10752 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_86
timestamp 1698175906
transform 1 0 10976 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_116
timestamp 1698175906
transform 1 0 14336 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_152
timestamp 1698175906
transform 1 0 18368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_165
timestamp 1698175906
transform 1 0 19824 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_173
timestamp 1698175906
transform 1 0 20720 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_177
timestamp 1698175906
transform 1 0 21168 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_200
timestamp 1698175906
transform 1 0 23744 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698175906
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_238
timestamp 1698175906
transform 1 0 28000 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_270
timestamp 1698175906
transform 1 0 31584 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_115
timestamp 1698175906
transform 1 0 14224 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_118
timestamp 1698175906
transform 1 0 14560 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_134
timestamp 1698175906
transform 1 0 16352 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_144
timestamp 1698175906
transform 1 0 17472 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_159
timestamp 1698175906
transform 1 0 19152 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_206
timestamp 1698175906
transform 1 0 24416 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_210
timestamp 1698175906
transform 1 0 24864 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_242
timestamp 1698175906
transform 1 0 28448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 4480 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_88
timestamp 1698175906
transform 1 0 11200 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_120
timestamp 1698175906
transform 1 0 14784 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_124
timestamp 1698175906
transform 1 0 15232 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_171
timestamp 1698175906
transform 1 0 20496 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_175
timestamp 1698175906
transform 1 0 20944 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698175906
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_220
timestamp 1698175906
transform 1 0 25984 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_226
timestamp 1698175906
transform 1 0 26656 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_258
timestamp 1698175906
transform 1 0 30240 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_274
timestamp 1698175906
transform 1 0 32032 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698175906
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 40320 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_69
timestamp 1698175906
transform 1 0 9072 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_85
timestamp 1698175906
transform 1 0 10864 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_93
timestamp 1698175906
transform 1 0 11760 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_97
timestamp 1698175906
transform 1 0 12208 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_99
timestamp 1698175906
transform 1 0 12432 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_119
timestamp 1698175906
transform 1 0 14672 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_135
timestamp 1698175906
transform 1 0 16464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_139
timestamp 1698175906
transform 1 0 16912 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_141
timestamp 1698175906
transform 1 0 17136 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_148
timestamp 1698175906
transform 1 0 17920 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_164
timestamp 1698175906
transform 1 0 19712 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698175906
transform 1 0 20608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_185
timestamp 1698175906
transform 1 0 22064 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_201
timestamp 1698175906
transform 1 0 23856 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_209
timestamp 1698175906
transform 1 0 24752 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_211
timestamp 1698175906
transform 1 0 24976 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_228
timestamp 1698175906
transform 1 0 26880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_236
timestamp 1698175906
transform 1 0 27776 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 4480 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 8064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_88
timestamp 1698175906
transform 1 0 11200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_124
timestamp 1698175906
transform 1 0 15232 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_128
timestamp 1698175906
transform 1 0 15680 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698175906
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_157
timestamp 1698175906
transform 1 0 18928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_161
timestamp 1698175906
transform 1 0 19376 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_198
timestamp 1698175906
transform 1 0 23520 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_202
timestamp 1698175906
transform 1 0 23968 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_241
timestamp 1698175906
transform 1 0 28336 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_245
timestamp 1698175906
transform 1 0 28784 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698175906
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 36512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 37408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_111
timestamp 1698175906
transform 1 0 13776 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_124
timestamp 1698175906
transform 1 0 15232 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_126
timestamp 1698175906
transform 1 0 15456 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_169
timestamp 1698175906
transform 1 0 20272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_173
timestamp 1698175906
transform 1 0 20720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_181
timestamp 1698175906
transform 1 0 21616 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_200
timestamp 1698175906
transform 1 0 23744 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_204
timestamp 1698175906
transform 1 0 24192 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_234
timestamp 1698175906
transform 1 0 27552 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_238
timestamp 1698175906
transform 1 0 28000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698175906
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 4480 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_136
timestamp 1698175906
transform 1 0 16576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_171
timestamp 1698175906
transform 1 0 20496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_175
timestamp 1698175906
transform 1 0 20944 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_205
timestamp 1698175906
transform 1 0 24304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_225
timestamp 1698175906
transform 1 0 26544 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_257
timestamp 1698175906
transform 1 0 30128 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_273
timestamp 1698175906
transform 1 0 31920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 32368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 36512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 37408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698175906
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698175906
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698175906
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_158
timestamp 1698175906
transform 1 0 19040 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_162
timestamp 1698175906
transform 1 0 19488 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_189
timestamp 1698175906
transform 1 0 22512 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_205
timestamp 1698175906
transform 1 0 24304 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita48_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita48_26
timestamp 1698175906
transform 1 0 39984 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform -1 0 4480 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 37520 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 21616 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 37520 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 37520 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 37520 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform -1 0 4480 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 24192 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 21280 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform -1 0 4480 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 4480 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform -1 0 20384 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 4480 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 19600 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 41200 17472 42000 17584 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 41200 16800 42000 16912 0 FreeSans 448 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 41200 5376 42000 5488 0 FreeSans 448 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 41200 25536 42000 25648 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 41200 24864 42000 24976 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 41200 24192 42000 24304 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 15456 800 15568 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 41200 20160 42000 20272 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 18144 41200 18256 42000 0 FreeSans 448 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 41200 21504 42000 21616 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 19488 41200 19600 42000 0 FreeSans 448 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 23520 41200 23632 42000 0 FreeSans 448 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 19096 25872 19096 25872 0 _000_
rlabel metal2 26208 18648 26208 18648 0 _001_
rlabel metal3 17136 24920 17136 24920 0 _002_
rlabel metal2 22008 25872 22008 25872 0 _003_
rlabel metal3 21560 20664 21560 20664 0 _004_
rlabel metal2 15736 15568 15736 15568 0 _005_
rlabel metal3 13104 20552 13104 20552 0 _006_
rlabel metal2 12040 21896 12040 21896 0 _007_
rlabel metal2 12600 24248 12600 24248 0 _008_
rlabel metal2 13776 23240 13776 23240 0 _009_
rlabel metal2 19544 14504 19544 14504 0 _010_
rlabel metal2 21448 24080 21448 24080 0 _011_
rlabel metal3 13720 15176 13720 15176 0 _012_
rlabel metal2 25368 24696 25368 24696 0 _013_
rlabel metal2 14224 13832 14224 13832 0 _014_
rlabel metal2 12824 17080 12824 17080 0 _015_
rlabel metal2 17976 22736 17976 22736 0 _016_
rlabel metal2 21896 18872 21896 18872 0 _017_
rlabel metal2 22120 21952 22120 21952 0 _018_
rlabel metal2 26600 20804 26600 20804 0 _019_
rlabel metal2 26264 23968 26264 23968 0 _020_
rlabel metal2 25032 16240 25032 16240 0 _021_
rlabel metal3 25592 16968 25592 16968 0 _022_
rlabel metal2 18872 16744 18872 16744 0 _023_
rlabel metal2 22120 23912 22120 23912 0 _024_
rlabel metal2 14616 15120 14616 15120 0 _025_
rlabel metal2 14672 15288 14672 15288 0 _026_
rlabel metal2 25928 25088 25928 25088 0 _027_
rlabel metal2 14784 14392 14784 14392 0 _028_
rlabel metal3 15288 16184 15288 16184 0 _029_
rlabel metal2 14504 16800 14504 16800 0 _030_
rlabel metal2 15064 17024 15064 17024 0 _031_
rlabel metal3 18480 22232 18480 22232 0 _032_
rlabel metal2 23128 21336 23128 21336 0 _033_
rlabel metal2 22568 21560 22568 21560 0 _034_
rlabel metal3 27384 21560 27384 21560 0 _035_
rlabel metal2 26600 23520 26600 23520 0 _036_
rlabel metal2 24360 16912 24360 16912 0 _037_
rlabel metal2 24024 17136 24024 17136 0 _038_
rlabel metal3 25760 17528 25760 17528 0 _039_
rlabel metal2 24808 17976 24808 17976 0 _040_
rlabel metal3 21952 18424 21952 18424 0 _041_
rlabel metal3 22456 17864 22456 17864 0 _042_
rlabel metal2 21448 17920 21448 17920 0 _043_
rlabel metal2 18872 18704 18872 18704 0 _044_
rlabel metal2 26824 18088 26824 18088 0 _045_
rlabel metal3 17080 21560 17080 21560 0 _046_
rlabel metal2 20328 18816 20328 18816 0 _047_
rlabel metal2 21672 23408 21672 23408 0 _048_
rlabel metal3 17136 19992 17136 19992 0 _049_
rlabel metal2 23016 24192 23016 24192 0 _050_
rlabel metal2 18760 24864 18760 24864 0 _051_
rlabel metal2 19824 25704 19824 25704 0 _052_
rlabel metal2 26376 23632 26376 23632 0 _053_
rlabel metal2 26656 19320 26656 19320 0 _054_
rlabel metal3 23576 21448 23576 21448 0 _055_
rlabel metal2 20552 21168 20552 21168 0 _056_
rlabel metal2 20216 21280 20216 21280 0 _057_
rlabel metal2 25480 21168 25480 21168 0 _058_
rlabel metal2 25816 19880 25816 19880 0 _059_
rlabel metal2 15624 17976 15624 17976 0 _060_
rlabel metal2 16520 17808 16520 17808 0 _061_
rlabel metal2 17472 22344 17472 22344 0 _062_
rlabel metal2 26096 21560 26096 21560 0 _063_
rlabel metal2 19488 21672 19488 21672 0 _064_
rlabel metal2 17080 21784 17080 21784 0 _065_
rlabel metal2 21896 24584 21896 24584 0 _066_
rlabel metal2 18424 24752 18424 24752 0 _067_
rlabel metal2 26376 25648 26376 25648 0 _068_
rlabel metal2 22568 25536 22568 25536 0 _069_
rlabel metal2 18368 15512 18368 15512 0 _070_
rlabel metal2 15512 15232 15512 15232 0 _071_
rlabel metal2 26152 23128 26152 23128 0 _072_
rlabel metal2 14840 18816 14840 18816 0 _073_
rlabel metal2 13944 22176 13944 22176 0 _074_
rlabel metal2 14280 18032 14280 18032 0 _075_
rlabel metal3 13552 23800 13552 23800 0 _076_
rlabel metal2 13944 24304 13944 24304 0 _077_
rlabel metal2 21448 22904 21448 22904 0 _078_
rlabel metal2 19432 15624 19432 15624 0 _079_
rlabel metal2 15624 16408 15624 16408 0 _080_
rlabel metal2 20216 17248 20216 17248 0 _081_
rlabel metal2 15960 18368 15960 18368 0 _082_
rlabel metal3 16744 15064 16744 15064 0 _083_
rlabel metal3 2478 23576 2478 23576 0 clk
rlabel metal2 21896 20440 21896 20440 0 clknet_0_clk
rlabel metal2 11368 23128 11368 23128 0 clknet_1_0__leaf_clk
rlabel metal3 25032 22120 25032 22120 0 clknet_1_1__leaf_clk
rlabel metal3 21392 15176 21392 15176 0 dut48.count\[0\]
rlabel metal3 19264 15288 19264 15288 0 dut48.count\[1\]
rlabel metal2 15176 21728 15176 21728 0 dut48.count\[2\]
rlabel metal2 14168 21504 14168 21504 0 dut48.count\[3\]
rlabel metal2 14056 26208 14056 26208 0 net1
rlabel metal2 27720 20944 27720 20944 0 net10
rlabel metal2 27608 23856 27608 23856 0 net11
rlabel metal2 28168 24136 28168 24136 0 net12
rlabel metal2 11032 15624 11032 15624 0 net13
rlabel metal3 23856 21672 23856 21672 0 net14
rlabel metal3 23576 21784 23576 21784 0 net15
rlabel metal3 23296 25256 23296 25256 0 net16
rlabel metal2 21784 3808 21784 3808 0 net17
rlabel metal2 14728 25816 14728 25816 0 net18
rlabel metal2 14504 24640 14504 24640 0 net19
rlabel metal2 25928 17584 25928 17584 0 net2
rlabel metal2 18648 26096 18648 26096 0 net20
rlabel metal3 27776 21672 27776 21672 0 net21
rlabel metal2 17416 23072 17416 23072 0 net22
rlabel metal2 20216 26488 20216 26488 0 net23
rlabel metal3 23800 25368 23800 25368 0 net24
rlabel metal2 15512 2030 15512 2030 0 net25
rlabel metal2 40264 5712 40264 5712 0 net26
rlabel metal2 16296 13552 16296 13552 0 net3
rlabel metal2 10696 16856 10696 16856 0 net4
rlabel metal2 28168 16800 28168 16800 0 net5
rlabel metal2 21896 9296 21896 9296 0 net6
rlabel metal2 4312 25200 4312 25200 0 net7
rlabel metal2 21336 6748 21336 6748 0 net8
rlabel metal2 26264 25984 26264 25984 0 net9
rlabel metal3 1358 26264 1358 26264 0 segm[0]
rlabel metal2 40040 17640 40040 17640 0 segm[10]
rlabel metal2 16184 2086 16184 2086 0 segm[11]
rlabel metal3 1358 16856 1358 16856 0 segm[12]
rlabel metal2 40040 16800 40040 16800 0 segm[13]
rlabel metal2 21560 2422 21560 2422 0 segm[2]
rlabel metal3 1414 24920 1414 24920 0 segm[3]
rlabel metal2 20888 2982 20888 2982 0 segm[5]
rlabel metal2 39928 25872 39928 25872 0 segm[6]
rlabel metal3 40642 20888 40642 20888 0 segm[7]
rlabel metal2 40040 25256 40040 25256 0 segm[8]
rlabel metal2 40040 24360 40040 24360 0 segm[9]
rlabel metal3 1358 15512 1358 15512 0 sel[0]
rlabel metal3 40642 20216 40642 20216 0 sel[10]
rlabel metal2 40040 22344 40040 22344 0 sel[11]
rlabel metal2 22232 39690 22232 39690 0 sel[1]
rlabel metal2 22232 2030 22232 2030 0 sel[2]
rlabel metal3 1358 25592 1358 25592 0 sel[3]
rlabel metal3 1358 24248 1358 24248 0 sel[4]
rlabel metal2 18200 39690 18200 39690 0 sel[5]
rlabel metal2 40040 21504 40040 21504 0 sel[6]
rlabel metal3 1358 22904 1358 22904 0 sel[7]
rlabel metal2 19544 39354 19544 39354 0 sel[8]
rlabel metal2 23576 39746 23576 39746 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
