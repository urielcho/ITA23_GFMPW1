magic
tech gf180mcuD
magscale 1 5
timestamp 1699643938
<< obsm1 >>
rect 672 1538 20328 19238
<< metal2 >>
rect 8400 20600 8456 21000
rect 8736 20600 8792 21000
rect 9744 20600 9800 21000
rect 10416 20600 10472 21000
rect 11424 20600 11480 21000
rect 12768 20600 12824 21000
rect 8736 0 8792 400
rect 9744 0 9800 400
rect 10080 0 10136 400
rect 11088 0 11144 400
rect 11760 0 11816 400
rect 12432 0 12488 400
<< obsm2 >>
rect 966 20570 8370 20600
rect 8486 20570 8706 20600
rect 8822 20570 9714 20600
rect 9830 20570 10386 20600
rect 10502 20570 11394 20600
rect 11510 20570 12738 20600
rect 12854 20570 20146 20600
rect 966 430 20146 20570
rect 966 400 8706 430
rect 8822 400 9714 430
rect 9830 400 10050 430
rect 10166 400 11058 430
rect 11174 400 11730 430
rect 11846 400 12402 430
rect 12518 400 20146 430
<< metal3 >>
rect 20600 17136 21000 17192
rect 0 14112 400 14168
rect 0 11760 400 11816
rect 20600 11760 21000 11816
rect 20600 11424 21000 11480
rect 20600 11088 21000 11144
rect 20600 10080 21000 10136
rect 20600 9744 21000 9800
rect 20600 9408 21000 9464
rect 20600 9072 21000 9128
rect 0 8736 400 8792
rect 20600 8736 21000 8792
rect 0 8064 400 8120
rect 0 7728 400 7784
rect 20600 7728 21000 7784
<< obsm3 >>
rect 400 17222 20600 19306
rect 400 17106 20570 17222
rect 400 14198 20600 17106
rect 430 14082 20600 14198
rect 400 11846 20600 14082
rect 430 11730 20570 11846
rect 400 11510 20600 11730
rect 400 11394 20570 11510
rect 400 11174 20600 11394
rect 400 11058 20570 11174
rect 400 10166 20600 11058
rect 400 10050 20570 10166
rect 400 9830 20600 10050
rect 400 9714 20570 9830
rect 400 9494 20600 9714
rect 400 9378 20570 9494
rect 400 9158 20600 9378
rect 400 9042 20570 9158
rect 400 8822 20600 9042
rect 430 8706 20570 8822
rect 400 8150 20600 8706
rect 430 8034 20600 8150
rect 400 7814 20600 8034
rect 430 7698 20570 7814
rect 400 1554 20600 7698
<< metal4 >>
rect 2224 1538 2384 19238
rect 9904 1538 10064 19238
rect 17584 1538 17744 19238
<< labels >>
rlabel metal3 s 0 14112 400 14168 6 clk
port 1 nsew signal input
rlabel metal2 s 9744 20600 9800 21000 6 segm[0]
port 2 nsew signal output
rlabel metal3 s 20600 9072 21000 9128 6 segm[10]
port 3 nsew signal output
rlabel metal3 s 0 8736 400 8792 6 segm[11]
port 4 nsew signal output
rlabel metal3 s 0 8064 400 8120 6 segm[12]
port 5 nsew signal output
rlabel metal2 s 10080 0 10136 400 6 segm[13]
port 6 nsew signal output
rlabel metal3 s 20600 11424 21000 11480 6 segm[1]
port 7 nsew signal output
rlabel metal3 s 20600 10080 21000 10136 6 segm[2]
port 8 nsew signal output
rlabel metal3 s 20600 17136 21000 17192 6 segm[3]
port 9 nsew signal output
rlabel metal3 s 20600 11760 21000 11816 6 segm[4]
port 10 nsew signal output
rlabel metal3 s 20600 9408 21000 9464 6 segm[5]
port 11 nsew signal output
rlabel metal3 s 0 7728 400 7784 6 segm[6]
port 12 nsew signal output
rlabel metal2 s 8736 0 8792 400 6 segm[7]
port 13 nsew signal output
rlabel metal2 s 12432 0 12488 400 6 segm[8]
port 14 nsew signal output
rlabel metal2 s 11760 0 11816 400 6 segm[9]
port 15 nsew signal output
rlabel metal2 s 8400 20600 8456 21000 6 sel[0]
port 16 nsew signal output
rlabel metal2 s 9744 0 9800 400 6 sel[10]
port 17 nsew signal output
rlabel metal3 s 20600 7728 21000 7784 6 sel[11]
port 18 nsew signal output
rlabel metal2 s 12768 20600 12824 21000 6 sel[1]
port 19 nsew signal output
rlabel metal2 s 10416 20600 10472 21000 6 sel[2]
port 20 nsew signal output
rlabel metal2 s 8736 20600 8792 21000 6 sel[3]
port 21 nsew signal output
rlabel metal3 s 20600 9744 21000 9800 6 sel[4]
port 22 nsew signal output
rlabel metal3 s 20600 11088 21000 11144 6 sel[5]
port 23 nsew signal output
rlabel metal3 s 20600 8736 21000 8792 6 sel[6]
port 24 nsew signal output
rlabel metal3 s 0 11760 400 11816 6 sel[7]
port 25 nsew signal output
rlabel metal2 s 11424 20600 11480 21000 6 sel[8]
port 26 nsew signal output
rlabel metal2 s 11088 0 11144 400 6 sel[9]
port 27 nsew signal output
rlabel metal4 s 2224 1538 2384 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 19238 6 vss
port 29 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 21000 21000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 507902
string GDS_FILE /home/urielcho/Proyectos_caravel/ITA23_GFMPW1b/openlane/ita20/runs/23_11_10_13_17/results/signoff/ita20.magic.gds
string GDS_START 170444
<< end >>

