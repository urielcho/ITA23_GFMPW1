magic
tech gf180mcuD
magscale 1 10
timestamp 1699643110
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 22430 38274 22482 38286
rect 22430 38210 22482 38222
rect 26126 38274 26178 38286
rect 26126 38210 26178 38222
rect 18834 38110 18846 38162
rect 18898 38110 18910 38162
rect 18050 37998 18062 38050
rect 18114 37998 18126 38050
rect 21522 37998 21534 38050
rect 21586 37998 21598 38050
rect 25218 37998 25230 38050
rect 25282 37998 25294 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 21422 37490 21474 37502
rect 21422 37426 21474 37438
rect 25790 37490 25842 37502
rect 25790 37426 25842 37438
rect 18274 37326 18286 37378
rect 18338 37326 18350 37378
rect 19618 37214 19630 37266
rect 19682 37214 19694 37266
rect 20514 37214 20526 37266
rect 20578 37214 20590 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 17602 27806 17614 27858
rect 17666 27806 17678 27858
rect 20974 27746 21026 27758
rect 18386 27694 18398 27746
rect 18450 27694 18462 27746
rect 20514 27694 20526 27746
rect 20578 27694 20590 27746
rect 20974 27682 21026 27694
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 25566 27298 25618 27310
rect 19394 27246 19406 27298
rect 19458 27295 19470 27298
rect 19730 27295 19742 27298
rect 19458 27249 19742 27295
rect 19458 27246 19470 27249
rect 19730 27246 19742 27249
rect 19794 27246 19806 27298
rect 25566 27234 25618 27246
rect 40014 27186 40066 27198
rect 18610 27134 18622 27186
rect 18674 27134 18686 27186
rect 25106 27134 25118 27186
rect 25170 27134 25182 27186
rect 40014 27122 40066 27134
rect 18846 27074 18898 27086
rect 15698 27022 15710 27074
rect 15762 27022 15774 27074
rect 18846 27010 18898 27022
rect 19182 27074 19234 27086
rect 19182 27010 19234 27022
rect 19854 27074 19906 27086
rect 26126 27074 26178 27086
rect 22306 27022 22318 27074
rect 22370 27022 22382 27074
rect 37650 27022 37662 27074
rect 37714 27022 37726 27074
rect 19854 27010 19906 27022
rect 26126 27010 26178 27022
rect 19070 26962 19122 26974
rect 16482 26910 16494 26962
rect 16546 26910 16558 26962
rect 19070 26898 19122 26910
rect 20078 26962 20130 26974
rect 20078 26898 20130 26910
rect 20190 26962 20242 26974
rect 20190 26898 20242 26910
rect 20638 26962 20690 26974
rect 20638 26898 20690 26910
rect 20750 26962 20802 26974
rect 20750 26898 20802 26910
rect 21310 26962 21362 26974
rect 21310 26898 21362 26910
rect 21534 26962 21586 26974
rect 21534 26898 21586 26910
rect 21646 26962 21698 26974
rect 25566 26962 25618 26974
rect 22978 26910 22990 26962
rect 23042 26910 23054 26962
rect 21646 26898 21698 26910
rect 25566 26898 25618 26910
rect 25678 26962 25730 26974
rect 25678 26898 25730 26910
rect 19630 26850 19682 26862
rect 19630 26786 19682 26798
rect 20414 26850 20466 26862
rect 20414 26786 20466 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 17390 26514 17442 26526
rect 23214 26514 23266 26526
rect 18386 26462 18398 26514
rect 18450 26462 18462 26514
rect 17390 26450 17442 26462
rect 23214 26450 23266 26462
rect 24110 26514 24162 26526
rect 24110 26450 24162 26462
rect 23438 26402 23490 26414
rect 20290 26350 20302 26402
rect 20354 26350 20366 26402
rect 23438 26338 23490 26350
rect 24222 26402 24274 26414
rect 26002 26350 26014 26402
rect 26066 26350 26078 26402
rect 24222 26338 24274 26350
rect 17726 26290 17778 26302
rect 17726 26226 17778 26238
rect 18734 26290 18786 26302
rect 23550 26290 23602 26302
rect 19618 26238 19630 26290
rect 19682 26238 19694 26290
rect 18734 26226 18786 26238
rect 23550 26226 23602 26238
rect 23886 26290 23938 26302
rect 25218 26238 25230 26290
rect 25282 26238 25294 26290
rect 23886 26226 23938 26238
rect 19182 26178 19234 26190
rect 28590 26178 28642 26190
rect 22418 26126 22430 26178
rect 22482 26126 22494 26178
rect 28130 26126 28142 26178
rect 28194 26126 28206 26178
rect 19182 26114 19234 26126
rect 28590 26114 28642 26126
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 25902 25730 25954 25742
rect 25902 25666 25954 25678
rect 1934 25618 1986 25630
rect 40014 25618 40066 25630
rect 13458 25566 13470 25618
rect 13522 25566 13534 25618
rect 1934 25554 1986 25566
rect 40014 25554 40066 25566
rect 25790 25506 25842 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 16258 25454 16270 25506
rect 16322 25454 16334 25506
rect 25218 25454 25230 25506
rect 25282 25454 25294 25506
rect 37650 25454 37662 25506
rect 37714 25454 37726 25506
rect 25790 25442 25842 25454
rect 20526 25394 20578 25406
rect 25902 25394 25954 25406
rect 15586 25342 15598 25394
rect 15650 25342 15662 25394
rect 24994 25342 25006 25394
rect 25058 25342 25070 25394
rect 20526 25330 20578 25342
rect 25902 25330 25954 25342
rect 16830 25282 16882 25294
rect 16830 25218 16882 25230
rect 20638 25282 20690 25294
rect 20638 25218 20690 25230
rect 20862 25282 20914 25294
rect 20862 25218 20914 25230
rect 22206 25282 22258 25294
rect 22206 25218 22258 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 16046 24946 16098 24958
rect 16046 24882 16098 24894
rect 16158 24946 16210 24958
rect 16158 24882 16210 24894
rect 29150 24946 29202 24958
rect 29150 24882 29202 24894
rect 15262 24834 15314 24846
rect 15262 24770 15314 24782
rect 15038 24722 15090 24734
rect 4274 24670 4286 24722
rect 4338 24670 4350 24722
rect 11554 24670 11566 24722
rect 11618 24670 11630 24722
rect 15038 24658 15090 24670
rect 15598 24722 15650 24734
rect 15598 24658 15650 24670
rect 19630 24722 19682 24734
rect 19954 24670 19966 24722
rect 20018 24670 20030 24722
rect 25890 24670 25902 24722
rect 25954 24670 25966 24722
rect 19630 24658 19682 24670
rect 15486 24610 15538 24622
rect 12226 24558 12238 24610
rect 12290 24558 12302 24610
rect 14354 24558 14366 24610
rect 14418 24558 14430 24610
rect 20738 24558 20750 24610
rect 20802 24558 20814 24610
rect 22866 24558 22878 24610
rect 22930 24558 22942 24610
rect 26562 24558 26574 24610
rect 26626 24558 26638 24610
rect 28690 24558 28702 24610
rect 28754 24558 28766 24610
rect 15486 24546 15538 24558
rect 1934 24498 1986 24510
rect 1934 24434 1986 24446
rect 15934 24498 15986 24510
rect 15934 24434 15986 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 12574 24162 12626 24174
rect 12574 24098 12626 24110
rect 17838 24162 17890 24174
rect 17838 24098 17890 24110
rect 21758 24050 21810 24062
rect 18610 23998 18622 24050
rect 18674 23998 18686 24050
rect 21758 23986 21810 23998
rect 23662 24050 23714 24062
rect 23662 23986 23714 23998
rect 26126 24050 26178 24062
rect 26126 23986 26178 23998
rect 40014 24050 40066 24062
rect 40014 23986 40066 23998
rect 14030 23938 14082 23950
rect 14030 23874 14082 23886
rect 14254 23938 14306 23950
rect 14254 23874 14306 23886
rect 14702 23938 14754 23950
rect 17278 23938 17330 23950
rect 17042 23886 17054 23938
rect 17106 23886 17118 23938
rect 14702 23874 14754 23886
rect 17278 23874 17330 23886
rect 17502 23938 17554 23950
rect 17502 23874 17554 23886
rect 17726 23938 17778 23950
rect 17726 23874 17778 23886
rect 19070 23938 19122 23950
rect 21198 23938 21250 23950
rect 19730 23886 19742 23938
rect 19794 23886 19806 23938
rect 20626 23886 20638 23938
rect 20690 23886 20702 23938
rect 19070 23874 19122 23886
rect 21198 23874 21250 23886
rect 21646 23938 21698 23950
rect 24222 23938 24274 23950
rect 22530 23886 22542 23938
rect 22594 23886 22606 23938
rect 23426 23886 23438 23938
rect 23490 23886 23502 23938
rect 21646 23874 21698 23886
rect 24222 23874 24274 23886
rect 26686 23938 26738 23950
rect 26686 23874 26738 23886
rect 26910 23938 26962 23950
rect 26910 23874 26962 23886
rect 27694 23938 27746 23950
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 27694 23874 27746 23886
rect 12910 23826 12962 23838
rect 12910 23762 12962 23774
rect 14142 23826 14194 23838
rect 23774 23826 23826 23838
rect 22306 23774 22318 23826
rect 22370 23774 22382 23826
rect 22978 23774 22990 23826
rect 23042 23774 23054 23826
rect 14142 23762 14194 23774
rect 23774 23762 23826 23774
rect 26238 23826 26290 23838
rect 27918 23826 27970 23838
rect 27234 23774 27246 23826
rect 27298 23774 27310 23826
rect 26238 23762 26290 23774
rect 27918 23762 27970 23774
rect 28030 23826 28082 23838
rect 28030 23762 28082 23774
rect 29262 23826 29314 23838
rect 29262 23762 29314 23774
rect 29374 23826 29426 23838
rect 29374 23762 29426 23774
rect 12686 23714 12738 23726
rect 12686 23650 12738 23662
rect 15038 23714 15090 23726
rect 15038 23650 15090 23662
rect 18622 23714 18674 23726
rect 18622 23650 18674 23662
rect 18734 23714 18786 23726
rect 18734 23650 18786 23662
rect 18958 23714 19010 23726
rect 21870 23714 21922 23726
rect 19506 23662 19518 23714
rect 19570 23662 19582 23714
rect 20402 23662 20414 23714
rect 20466 23662 20478 23714
rect 18958 23650 19010 23662
rect 21870 23650 21922 23662
rect 24110 23714 24162 23726
rect 24110 23650 24162 23662
rect 26014 23714 26066 23726
rect 26014 23650 26066 23662
rect 29038 23714 29090 23726
rect 29038 23650 29090 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 16942 23378 16994 23390
rect 24446 23378 24498 23390
rect 23538 23326 23550 23378
rect 23602 23326 23614 23378
rect 16942 23314 16994 23326
rect 24446 23314 24498 23326
rect 27470 23378 27522 23390
rect 27470 23314 27522 23326
rect 18286 23266 18338 23278
rect 21310 23266 21362 23278
rect 20514 23214 20526 23266
rect 20578 23214 20590 23266
rect 22978 23214 22990 23266
rect 23042 23214 23054 23266
rect 23202 23214 23214 23266
rect 23266 23214 23278 23266
rect 18286 23202 18338 23214
rect 21310 23202 21362 23214
rect 17390 23154 17442 23166
rect 4274 23102 4286 23154
rect 4338 23102 4350 23154
rect 13794 23102 13806 23154
rect 13858 23102 13870 23154
rect 14466 23102 14478 23154
rect 14530 23102 14542 23154
rect 17390 23090 17442 23102
rect 17502 23154 17554 23166
rect 17502 23090 17554 23102
rect 17614 23154 17666 23166
rect 17614 23090 17666 23102
rect 18062 23154 18114 23166
rect 21086 23154 21138 23166
rect 18498 23102 18510 23154
rect 18562 23102 18574 23154
rect 18722 23102 18734 23154
rect 18786 23102 18798 23154
rect 19282 23102 19294 23154
rect 19346 23102 19358 23154
rect 20178 23102 20190 23154
rect 20242 23102 20254 23154
rect 18062 23090 18114 23102
rect 21086 23090 21138 23102
rect 21422 23154 21474 23166
rect 23998 23154 24050 23166
rect 22194 23102 22206 23154
rect 22258 23102 22270 23154
rect 22642 23102 22654 23154
rect 22706 23102 22718 23154
rect 21422 23090 21474 23102
rect 23998 23090 24050 23102
rect 24670 23154 24722 23166
rect 27794 23102 27806 23154
rect 27858 23102 27870 23154
rect 24670 23090 24722 23102
rect 14254 23042 14306 23054
rect 10882 22990 10894 23042
rect 10946 22990 10958 23042
rect 13010 22990 13022 23042
rect 13074 22990 13086 23042
rect 14254 22978 14306 22990
rect 14926 23042 14978 23054
rect 21758 23042 21810 23054
rect 19506 22990 19518 23042
rect 19570 22990 19582 23042
rect 20402 22990 20414 23042
rect 20466 22990 20478 23042
rect 14926 22978 14978 22990
rect 21758 22978 21810 22990
rect 24558 23042 24610 23054
rect 28578 22990 28590 23042
rect 28642 22990 28654 23042
rect 30706 22990 30718 23042
rect 30770 22990 30782 23042
rect 24558 22978 24610 22990
rect 1934 22930 1986 22942
rect 1934 22866 1986 22878
rect 14142 22930 14194 22942
rect 14142 22866 14194 22878
rect 18174 22930 18226 22942
rect 18174 22866 18226 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 19630 22594 19682 22606
rect 19630 22530 19682 22542
rect 20414 22594 20466 22606
rect 20414 22530 20466 22542
rect 26462 22594 26514 22606
rect 26462 22530 26514 22542
rect 28478 22594 28530 22606
rect 28478 22530 28530 22542
rect 14030 22482 14082 22494
rect 14030 22418 14082 22430
rect 17166 22482 17218 22494
rect 19854 22482 19906 22494
rect 17714 22430 17726 22482
rect 17778 22430 17790 22482
rect 17166 22418 17218 22430
rect 19854 22418 19906 22430
rect 20750 22482 20802 22494
rect 26574 22482 26626 22494
rect 25890 22430 25902 22482
rect 25954 22430 25966 22482
rect 20750 22418 20802 22430
rect 26574 22418 26626 22430
rect 13582 22370 13634 22382
rect 13582 22306 13634 22318
rect 13806 22370 13858 22382
rect 23886 22370 23938 22382
rect 28590 22370 28642 22382
rect 17602 22318 17614 22370
rect 17666 22318 17678 22370
rect 18498 22318 18510 22370
rect 18562 22318 18574 22370
rect 22082 22318 22094 22370
rect 22146 22318 22158 22370
rect 24994 22318 25006 22370
rect 25058 22318 25070 22370
rect 25554 22318 25566 22370
rect 25618 22318 25630 22370
rect 13806 22306 13858 22318
rect 23886 22306 23938 22318
rect 28590 22306 28642 22318
rect 14142 22258 14194 22270
rect 16830 22258 16882 22270
rect 20526 22258 20578 22270
rect 22654 22258 22706 22270
rect 28030 22258 28082 22270
rect 16034 22206 16046 22258
rect 16098 22206 16110 22258
rect 17938 22206 17950 22258
rect 18002 22206 18014 22258
rect 21410 22206 21422 22258
rect 21474 22206 21486 22258
rect 25666 22206 25678 22258
rect 25730 22206 25742 22258
rect 14142 22194 14194 22206
rect 16830 22194 16882 22206
rect 20526 22194 20578 22206
rect 22654 22194 22706 22206
rect 28030 22194 28082 22206
rect 28478 22258 28530 22270
rect 28478 22194 28530 22206
rect 16382 22146 16434 22158
rect 16382 22082 16434 22094
rect 17054 22146 17106 22158
rect 17054 22082 17106 22094
rect 17278 22146 17330 22158
rect 21758 22146 21810 22158
rect 19282 22094 19294 22146
rect 19346 22094 19358 22146
rect 17278 22082 17330 22094
rect 21758 22082 21810 22094
rect 24446 22146 24498 22158
rect 24446 22082 24498 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 16270 21810 16322 21822
rect 23326 21810 23378 21822
rect 22978 21758 22990 21810
rect 23042 21758 23054 21810
rect 16270 21746 16322 21758
rect 23326 21746 23378 21758
rect 17602 21646 17614 21698
rect 17666 21646 17678 21698
rect 27346 21646 27358 21698
rect 27410 21646 27422 21698
rect 29374 21586 29426 21598
rect 22642 21534 22654 21586
rect 22706 21534 22718 21586
rect 28018 21534 28030 21586
rect 28082 21534 28094 21586
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 29374 21522 29426 21534
rect 16830 21474 16882 21486
rect 28926 21474 28978 21486
rect 25218 21422 25230 21474
rect 25282 21422 25294 21474
rect 16830 21410 16882 21422
rect 28926 21410 28978 21422
rect 28814 21362 28866 21374
rect 28814 21298 28866 21310
rect 40014 21362 40066 21374
rect 40014 21298 40066 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 16382 21026 16434 21038
rect 18610 20974 18622 21026
rect 18674 20974 18686 21026
rect 19394 20974 19406 21026
rect 19458 20974 19470 21026
rect 21858 20974 21870 21026
rect 21922 20974 21934 21026
rect 16382 20962 16434 20974
rect 19618 20862 19630 20914
rect 19682 20862 19694 20914
rect 22866 20862 22878 20914
rect 22930 20862 22942 20914
rect 27906 20862 27918 20914
rect 27970 20862 27982 20914
rect 29250 20862 29262 20914
rect 29314 20862 29326 20914
rect 39778 20862 39790 20914
rect 39842 20862 39854 20914
rect 14478 20802 14530 20814
rect 14478 20738 14530 20750
rect 14702 20802 14754 20814
rect 20078 20802 20130 20814
rect 17490 20750 17502 20802
rect 17554 20750 17566 20802
rect 18274 20750 18286 20802
rect 18338 20750 18350 20802
rect 18722 20750 18734 20802
rect 18786 20750 18798 20802
rect 19842 20750 19854 20802
rect 19906 20750 19918 20802
rect 14702 20738 14754 20750
rect 20078 20738 20130 20750
rect 21310 20802 21362 20814
rect 21310 20738 21362 20750
rect 21534 20802 21586 20814
rect 22530 20750 22542 20802
rect 22594 20750 22606 20802
rect 23314 20750 23326 20802
rect 23378 20750 23390 20802
rect 29138 20750 29150 20802
rect 29202 20750 29214 20802
rect 29810 20750 29822 20802
rect 29874 20750 29886 20802
rect 37650 20750 37662 20802
rect 37714 20750 37726 20802
rect 21534 20738 21586 20750
rect 14030 20690 14082 20702
rect 14030 20626 14082 20638
rect 16494 20690 16546 20702
rect 30158 20690 30210 20702
rect 17602 20638 17614 20690
rect 17666 20638 17678 20690
rect 16494 20626 16546 20638
rect 30158 20626 30210 20638
rect 13918 20578 13970 20590
rect 13918 20514 13970 20526
rect 14254 20578 14306 20590
rect 14254 20514 14306 20526
rect 29374 20578 29426 20590
rect 29374 20514 29426 20526
rect 29598 20578 29650 20590
rect 29598 20514 29650 20526
rect 30270 20578 30322 20590
rect 30270 20514 30322 20526
rect 30494 20578 30546 20590
rect 30494 20514 30546 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 40238 20242 40290 20254
rect 40238 20178 40290 20190
rect 16830 20130 16882 20142
rect 16830 20066 16882 20078
rect 18734 20130 18786 20142
rect 18734 20066 18786 20078
rect 19070 20130 19122 20142
rect 27134 20130 27186 20142
rect 23314 20078 23326 20130
rect 23378 20078 23390 20130
rect 28578 20078 28590 20130
rect 28642 20078 28654 20130
rect 19070 20066 19122 20078
rect 27134 20066 27186 20078
rect 16494 20018 16546 20030
rect 11554 19966 11566 20018
rect 11618 19966 11630 20018
rect 16494 19954 16546 19966
rect 17390 20018 17442 20030
rect 17390 19954 17442 19966
rect 18398 20018 18450 20030
rect 26910 20018 26962 20030
rect 19394 19966 19406 20018
rect 19458 19966 19470 20018
rect 18398 19954 18450 19966
rect 26910 19954 26962 19966
rect 27582 20018 27634 20030
rect 27794 19966 27806 20018
rect 27858 19966 27870 20018
rect 27582 19954 27634 19966
rect 14814 19906 14866 19918
rect 12226 19854 12238 19906
rect 12290 19854 12302 19906
rect 14354 19854 14366 19906
rect 14418 19854 14430 19906
rect 14814 19842 14866 19854
rect 17950 19906 18002 19918
rect 17950 19842 18002 19854
rect 27022 19906 27074 19918
rect 30706 19854 30718 19906
rect 30770 19854 30782 19906
rect 27022 19842 27074 19854
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 19630 19458 19682 19470
rect 19630 19394 19682 19406
rect 21646 19458 21698 19470
rect 21646 19394 21698 19406
rect 21870 19458 21922 19470
rect 26898 19406 26910 19458
rect 26962 19455 26974 19458
rect 27122 19455 27134 19458
rect 26962 19409 27134 19455
rect 26962 19406 26974 19409
rect 27122 19406 27134 19409
rect 27186 19406 27198 19458
rect 21870 19394 21922 19406
rect 20750 19346 20802 19358
rect 20750 19282 20802 19294
rect 21422 19346 21474 19358
rect 21422 19282 21474 19294
rect 14366 19234 14418 19246
rect 14130 19182 14142 19234
rect 14194 19182 14206 19234
rect 14366 19170 14418 19182
rect 16494 19234 16546 19246
rect 16494 19170 16546 19182
rect 18286 19234 18338 19246
rect 18286 19170 18338 19182
rect 18958 19234 19010 19246
rect 23662 19234 23714 19246
rect 20290 19182 20302 19234
rect 20354 19182 20366 19234
rect 23202 19182 23214 19234
rect 23266 19182 23278 19234
rect 18958 19170 19010 19182
rect 23662 19170 23714 19182
rect 12574 19122 12626 19134
rect 12574 19058 12626 19070
rect 12910 19122 12962 19134
rect 12910 19058 12962 19070
rect 13470 19122 13522 19134
rect 13470 19058 13522 19070
rect 16046 19122 16098 19134
rect 16046 19058 16098 19070
rect 16830 19122 16882 19134
rect 16830 19058 16882 19070
rect 18174 19122 18226 19134
rect 22978 19070 22990 19122
rect 23042 19070 23054 19122
rect 18174 19058 18226 19070
rect 16158 19010 16210 19022
rect 17502 19010 17554 19022
rect 17154 18958 17166 19010
rect 17218 18958 17230 19010
rect 16158 18946 16210 18958
rect 17502 18946 17554 18958
rect 17950 19010 18002 19022
rect 19406 19010 19458 19022
rect 18610 18958 18622 19010
rect 18674 18958 18686 19010
rect 17950 18946 18002 18958
rect 19406 18946 19458 18958
rect 19518 19010 19570 19022
rect 19518 18946 19570 18958
rect 22318 19010 22370 19022
rect 22318 18946 22370 18958
rect 23774 19010 23826 19022
rect 23774 18946 23826 18958
rect 23998 19010 24050 19022
rect 23998 18946 24050 18958
rect 26910 19010 26962 19022
rect 26910 18946 26962 18958
rect 27470 19010 27522 19022
rect 27470 18946 27522 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 19182 18674 19234 18686
rect 22206 18674 22258 18686
rect 19618 18622 19630 18674
rect 19682 18622 19694 18674
rect 21074 18622 21086 18674
rect 21138 18622 21150 18674
rect 25554 18622 25566 18674
rect 25618 18622 25630 18674
rect 19182 18610 19234 18622
rect 22206 18610 22258 18622
rect 18846 18562 18898 18574
rect 21982 18562 22034 18574
rect 20402 18510 20414 18562
rect 20466 18510 20478 18562
rect 18846 18498 18898 18510
rect 21982 18498 22034 18510
rect 22654 18562 22706 18574
rect 22654 18498 22706 18510
rect 22766 18562 22818 18574
rect 28018 18510 28030 18562
rect 28082 18510 28094 18562
rect 22766 18498 22818 18510
rect 16158 18450 16210 18462
rect 19070 18450 19122 18462
rect 20750 18450 20802 18462
rect 12786 18398 12798 18450
rect 12850 18398 12862 18450
rect 13570 18398 13582 18450
rect 13634 18398 13646 18450
rect 18610 18398 18622 18450
rect 18674 18398 18686 18450
rect 19842 18398 19854 18450
rect 19906 18398 19918 18450
rect 16158 18386 16210 18398
rect 19070 18386 19122 18398
rect 20750 18386 20802 18398
rect 22094 18450 22146 18462
rect 25902 18450 25954 18462
rect 25218 18398 25230 18450
rect 25282 18398 25294 18450
rect 25442 18398 25454 18450
rect 25506 18398 25518 18450
rect 22094 18386 22146 18398
rect 25902 18386 25954 18398
rect 26126 18450 26178 18462
rect 27234 18398 27246 18450
rect 27298 18398 27310 18450
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 26126 18386 26178 18398
rect 18958 18338 19010 18350
rect 15698 18286 15710 18338
rect 15762 18286 15774 18338
rect 18958 18274 19010 18286
rect 21422 18338 21474 18350
rect 21422 18274 21474 18286
rect 21646 18338 21698 18350
rect 21646 18274 21698 18286
rect 25678 18338 25730 18350
rect 25678 18274 25730 18286
rect 26910 18338 26962 18350
rect 30146 18286 30158 18338
rect 30210 18286 30222 18338
rect 26910 18274 26962 18286
rect 22766 18226 22818 18238
rect 22766 18162 22818 18174
rect 26798 18226 26850 18238
rect 26798 18162 26850 18174
rect 40014 18226 40066 18238
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 28254 17890 28306 17902
rect 28254 17826 28306 17838
rect 1934 17778 1986 17790
rect 40014 17778 40066 17790
rect 25666 17726 25678 17778
rect 25730 17726 25742 17778
rect 27794 17726 27806 17778
rect 27858 17726 27870 17778
rect 1934 17714 1986 17726
rect 40014 17714 40066 17726
rect 14814 17666 14866 17678
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 14814 17602 14866 17614
rect 21646 17666 21698 17678
rect 24994 17614 25006 17666
rect 25058 17614 25070 17666
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 21646 17602 21698 17614
rect 14142 17554 14194 17566
rect 14142 17490 14194 17502
rect 14254 17554 14306 17566
rect 14254 17490 14306 17502
rect 14702 17554 14754 17566
rect 14702 17490 14754 17502
rect 20078 17554 20130 17566
rect 20078 17490 20130 17502
rect 28142 17554 28194 17566
rect 28142 17490 28194 17502
rect 28254 17554 28306 17566
rect 28254 17490 28306 17502
rect 13918 17442 13970 17454
rect 13918 17378 13970 17390
rect 14478 17442 14530 17454
rect 14478 17378 14530 17390
rect 20190 17442 20242 17454
rect 20190 17378 20242 17390
rect 20414 17442 20466 17454
rect 29262 17442 29314 17454
rect 21298 17390 21310 17442
rect 21362 17390 21374 17442
rect 20414 17378 20466 17390
rect 29262 17378 29314 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 15598 17106 15650 17118
rect 15598 17042 15650 17054
rect 23102 17106 23154 17118
rect 23102 17042 23154 17054
rect 24446 17106 24498 17118
rect 24446 17042 24498 17054
rect 18958 16994 19010 17006
rect 18958 16930 19010 16942
rect 19294 16994 19346 17006
rect 19294 16930 19346 16942
rect 22206 16994 22258 17006
rect 23326 16994 23378 17006
rect 22418 16942 22430 16994
rect 22482 16942 22494 16994
rect 22206 16930 22258 16942
rect 23326 16930 23378 16942
rect 23438 16994 23490 17006
rect 23438 16930 23490 16942
rect 24110 16994 24162 17006
rect 24110 16930 24162 16942
rect 30046 16994 30098 17006
rect 30046 16930 30098 16942
rect 14478 16882 14530 16894
rect 4274 16830 4286 16882
rect 4338 16830 4350 16882
rect 13458 16830 13470 16882
rect 13522 16830 13534 16882
rect 14130 16830 14142 16882
rect 14194 16830 14206 16882
rect 14478 16818 14530 16830
rect 14702 16882 14754 16894
rect 14702 16818 14754 16830
rect 14814 16882 14866 16894
rect 14814 16818 14866 16830
rect 15150 16882 15202 16894
rect 15150 16818 15202 16830
rect 22766 16882 22818 16894
rect 22766 16818 22818 16830
rect 24446 16882 24498 16894
rect 24446 16818 24498 16830
rect 24782 16882 24834 16894
rect 26674 16830 26686 16882
rect 26738 16830 26750 16882
rect 37874 16830 37886 16882
rect 37938 16830 37950 16882
rect 24782 16818 24834 16830
rect 21982 16770 22034 16782
rect 40014 16770 40066 16782
rect 11330 16718 11342 16770
rect 11394 16718 11406 16770
rect 27458 16718 27470 16770
rect 27522 16718 27534 16770
rect 29586 16718 29598 16770
rect 29650 16718 29662 16770
rect 21982 16706 22034 16718
rect 40014 16706 40066 16718
rect 1934 16658 1986 16670
rect 1934 16594 1986 16606
rect 22990 16658 23042 16670
rect 22990 16594 23042 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 14814 16322 14866 16334
rect 14814 16258 14866 16270
rect 19518 16322 19570 16334
rect 19518 16258 19570 16270
rect 27358 16210 27410 16222
rect 24210 16158 24222 16210
rect 24274 16158 24286 16210
rect 26338 16158 26350 16210
rect 26402 16158 26414 16210
rect 27358 16146 27410 16158
rect 40014 16210 40066 16222
rect 40014 16146 40066 16158
rect 13806 16098 13858 16110
rect 13806 16034 13858 16046
rect 14030 16098 14082 16110
rect 14030 16034 14082 16046
rect 14366 16098 14418 16110
rect 14366 16034 14418 16046
rect 14702 16098 14754 16110
rect 14702 16034 14754 16046
rect 18734 16098 18786 16110
rect 26910 16098 26962 16110
rect 19842 16046 19854 16098
rect 19906 16046 19918 16098
rect 23538 16046 23550 16098
rect 23602 16046 23614 16098
rect 18734 16034 18786 16046
rect 26910 16034 26962 16046
rect 27582 16098 27634 16110
rect 29250 16046 29262 16098
rect 29314 16046 29326 16098
rect 37650 16046 37662 16098
rect 37714 16046 37726 16098
rect 27582 16034 27634 16046
rect 14814 15986 14866 15998
rect 14814 15922 14866 15934
rect 17950 15986 18002 15998
rect 17950 15922 18002 15934
rect 27134 15986 27186 15998
rect 27134 15922 27186 15934
rect 13918 15874 13970 15886
rect 13918 15810 13970 15822
rect 17614 15874 17666 15886
rect 17614 15810 17666 15822
rect 17838 15874 17890 15886
rect 17838 15810 17890 15822
rect 18398 15874 18450 15886
rect 18398 15810 18450 15822
rect 19182 15874 19234 15886
rect 19182 15810 19234 15822
rect 19630 15874 19682 15886
rect 29474 15822 29486 15874
rect 29538 15822 29550 15874
rect 19630 15810 19682 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 14702 15538 14754 15550
rect 14702 15474 14754 15486
rect 16606 15538 16658 15550
rect 16606 15474 16658 15486
rect 18510 15538 18562 15550
rect 18510 15474 18562 15486
rect 18846 15538 18898 15550
rect 18846 15474 18898 15486
rect 20414 15538 20466 15550
rect 20414 15474 20466 15486
rect 20862 15538 20914 15550
rect 20862 15474 20914 15486
rect 23886 15538 23938 15550
rect 23886 15474 23938 15486
rect 25118 15538 25170 15550
rect 25118 15474 25170 15486
rect 26574 15538 26626 15550
rect 26574 15474 26626 15486
rect 17502 15426 17554 15438
rect 13458 15374 13470 15426
rect 13522 15374 13534 15426
rect 17502 15362 17554 15374
rect 17726 15426 17778 15438
rect 17726 15362 17778 15374
rect 20638 15426 20690 15438
rect 20638 15362 20690 15374
rect 22766 15426 22818 15438
rect 22766 15362 22818 15374
rect 25342 15426 25394 15438
rect 25342 15362 25394 15374
rect 25454 15426 25506 15438
rect 25454 15362 25506 15374
rect 16270 15314 16322 15326
rect 14242 15262 14254 15314
rect 14306 15262 14318 15314
rect 16270 15250 16322 15262
rect 16606 15314 16658 15326
rect 16606 15250 16658 15262
rect 16942 15314 16994 15326
rect 16942 15250 16994 15262
rect 17950 15314 18002 15326
rect 17950 15250 18002 15262
rect 18174 15314 18226 15326
rect 18174 15250 18226 15262
rect 18622 15314 18674 15326
rect 18622 15250 18674 15262
rect 18734 15314 18786 15326
rect 19294 15314 19346 15326
rect 19854 15314 19906 15326
rect 19058 15262 19070 15314
rect 19122 15262 19134 15314
rect 19618 15262 19630 15314
rect 19682 15262 19694 15314
rect 18734 15250 18786 15262
rect 19294 15250 19346 15262
rect 19854 15250 19906 15262
rect 20078 15314 20130 15326
rect 20078 15250 20130 15262
rect 20302 15314 20354 15326
rect 22978 15262 22990 15314
rect 23042 15262 23054 15314
rect 20302 15250 20354 15262
rect 23998 15202 24050 15214
rect 11330 15150 11342 15202
rect 11394 15150 11406 15202
rect 23998 15138 24050 15150
rect 20974 15090 21026 15102
rect 20974 15026 21026 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 25342 14642 25394 14654
rect 17042 14590 17054 14642
rect 17106 14590 17118 14642
rect 19170 14590 19182 14642
rect 19234 14590 19246 14642
rect 22754 14590 22766 14642
rect 22818 14590 22830 14642
rect 24882 14590 24894 14642
rect 24946 14590 24958 14642
rect 25342 14578 25394 14590
rect 19630 14530 19682 14542
rect 16258 14478 16270 14530
rect 16322 14478 16334 14530
rect 22082 14478 22094 14530
rect 22146 14478 22158 14530
rect 19630 14466 19682 14478
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 21074 13806 21086 13858
rect 21138 13806 21150 13858
rect 22318 13746 22370 13758
rect 21858 13694 21870 13746
rect 21922 13694 21934 13746
rect 22318 13682 22370 13694
rect 18946 13582 18958 13634
rect 19010 13582 19022 13634
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 18286 13074 18338 13086
rect 15586 13022 15598 13074
rect 15650 13022 15662 13074
rect 17714 13022 17726 13074
rect 17778 13022 17790 13074
rect 18286 13010 18338 13022
rect 14802 12910 14814 12962
rect 14866 12910 14878 12962
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 18398 4450 18450 4462
rect 18398 4386 18450 4398
rect 19058 4286 19070 4338
rect 19122 4286 19134 4338
rect 20078 4114 20130 4126
rect 20078 4050 20130 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 18622 3666 18674 3678
rect 18622 3602 18674 3614
rect 22094 3666 22146 3678
rect 22094 3602 22146 3614
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 17602 3502 17614 3554
rect 17666 3502 17678 3554
rect 21074 3502 21086 3554
rect 21138 3502 21150 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 22430 38222 22482 38274
rect 26126 38222 26178 38274
rect 18846 38110 18898 38162
rect 18062 37998 18114 38050
rect 21534 37998 21586 38050
rect 25230 37998 25282 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 21422 37438 21474 37490
rect 25790 37438 25842 37490
rect 18286 37326 18338 37378
rect 19630 37214 19682 37266
rect 20526 37214 20578 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 17614 27806 17666 27858
rect 18398 27694 18450 27746
rect 20526 27694 20578 27746
rect 20974 27694 21026 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 19406 27246 19458 27298
rect 19742 27246 19794 27298
rect 25566 27246 25618 27298
rect 18622 27134 18674 27186
rect 25118 27134 25170 27186
rect 40014 27134 40066 27186
rect 15710 27022 15762 27074
rect 18846 27022 18898 27074
rect 19182 27022 19234 27074
rect 19854 27022 19906 27074
rect 22318 27022 22370 27074
rect 26126 27022 26178 27074
rect 37662 27022 37714 27074
rect 16494 26910 16546 26962
rect 19070 26910 19122 26962
rect 20078 26910 20130 26962
rect 20190 26910 20242 26962
rect 20638 26910 20690 26962
rect 20750 26910 20802 26962
rect 21310 26910 21362 26962
rect 21534 26910 21586 26962
rect 21646 26910 21698 26962
rect 22990 26910 23042 26962
rect 25566 26910 25618 26962
rect 25678 26910 25730 26962
rect 19630 26798 19682 26850
rect 20414 26798 20466 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 17390 26462 17442 26514
rect 18398 26462 18450 26514
rect 23214 26462 23266 26514
rect 24110 26462 24162 26514
rect 20302 26350 20354 26402
rect 23438 26350 23490 26402
rect 24222 26350 24274 26402
rect 26014 26350 26066 26402
rect 17726 26238 17778 26290
rect 18734 26238 18786 26290
rect 19630 26238 19682 26290
rect 23550 26238 23602 26290
rect 23886 26238 23938 26290
rect 25230 26238 25282 26290
rect 19182 26126 19234 26178
rect 22430 26126 22482 26178
rect 28142 26126 28194 26178
rect 28590 26126 28642 26178
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 25902 25678 25954 25730
rect 1934 25566 1986 25618
rect 13470 25566 13522 25618
rect 40014 25566 40066 25618
rect 4286 25454 4338 25506
rect 16270 25454 16322 25506
rect 25230 25454 25282 25506
rect 25790 25454 25842 25506
rect 37662 25454 37714 25506
rect 15598 25342 15650 25394
rect 20526 25342 20578 25394
rect 25006 25342 25058 25394
rect 25902 25342 25954 25394
rect 16830 25230 16882 25282
rect 20638 25230 20690 25282
rect 20862 25230 20914 25282
rect 22206 25230 22258 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 16046 24894 16098 24946
rect 16158 24894 16210 24946
rect 29150 24894 29202 24946
rect 15262 24782 15314 24834
rect 4286 24670 4338 24722
rect 11566 24670 11618 24722
rect 15038 24670 15090 24722
rect 15598 24670 15650 24722
rect 19630 24670 19682 24722
rect 19966 24670 20018 24722
rect 25902 24670 25954 24722
rect 12238 24558 12290 24610
rect 14366 24558 14418 24610
rect 15486 24558 15538 24610
rect 20750 24558 20802 24610
rect 22878 24558 22930 24610
rect 26574 24558 26626 24610
rect 28702 24558 28754 24610
rect 1934 24446 1986 24498
rect 15934 24446 15986 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 12574 24110 12626 24162
rect 17838 24110 17890 24162
rect 18622 23998 18674 24050
rect 21758 23998 21810 24050
rect 23662 23998 23714 24050
rect 26126 23998 26178 24050
rect 40014 23998 40066 24050
rect 14030 23886 14082 23938
rect 14254 23886 14306 23938
rect 14702 23886 14754 23938
rect 17054 23886 17106 23938
rect 17278 23886 17330 23938
rect 17502 23886 17554 23938
rect 17726 23886 17778 23938
rect 19070 23886 19122 23938
rect 19742 23886 19794 23938
rect 20638 23886 20690 23938
rect 21198 23886 21250 23938
rect 21646 23886 21698 23938
rect 22542 23886 22594 23938
rect 23438 23886 23490 23938
rect 24222 23886 24274 23938
rect 26686 23886 26738 23938
rect 26910 23886 26962 23938
rect 27694 23886 27746 23938
rect 37662 23886 37714 23938
rect 12910 23774 12962 23826
rect 14142 23774 14194 23826
rect 22318 23774 22370 23826
rect 22990 23774 23042 23826
rect 23774 23774 23826 23826
rect 26238 23774 26290 23826
rect 27246 23774 27298 23826
rect 27918 23774 27970 23826
rect 28030 23774 28082 23826
rect 29262 23774 29314 23826
rect 29374 23774 29426 23826
rect 12686 23662 12738 23714
rect 15038 23662 15090 23714
rect 18622 23662 18674 23714
rect 18734 23662 18786 23714
rect 18958 23662 19010 23714
rect 19518 23662 19570 23714
rect 20414 23662 20466 23714
rect 21870 23662 21922 23714
rect 24110 23662 24162 23714
rect 26014 23662 26066 23714
rect 29038 23662 29090 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 16942 23326 16994 23378
rect 23550 23326 23602 23378
rect 24446 23326 24498 23378
rect 27470 23326 27522 23378
rect 18286 23214 18338 23266
rect 20526 23214 20578 23266
rect 21310 23214 21362 23266
rect 22990 23214 23042 23266
rect 23214 23214 23266 23266
rect 4286 23102 4338 23154
rect 13806 23102 13858 23154
rect 14478 23102 14530 23154
rect 17390 23102 17442 23154
rect 17502 23102 17554 23154
rect 17614 23102 17666 23154
rect 18062 23102 18114 23154
rect 18510 23102 18562 23154
rect 18734 23102 18786 23154
rect 19294 23102 19346 23154
rect 20190 23102 20242 23154
rect 21086 23102 21138 23154
rect 21422 23102 21474 23154
rect 22206 23102 22258 23154
rect 22654 23102 22706 23154
rect 23998 23102 24050 23154
rect 24670 23102 24722 23154
rect 27806 23102 27858 23154
rect 10894 22990 10946 23042
rect 13022 22990 13074 23042
rect 14254 22990 14306 23042
rect 14926 22990 14978 23042
rect 19518 22990 19570 23042
rect 20414 22990 20466 23042
rect 21758 22990 21810 23042
rect 24558 22990 24610 23042
rect 28590 22990 28642 23042
rect 30718 22990 30770 23042
rect 1934 22878 1986 22930
rect 14142 22878 14194 22930
rect 18174 22878 18226 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 19630 22542 19682 22594
rect 20414 22542 20466 22594
rect 26462 22542 26514 22594
rect 28478 22542 28530 22594
rect 14030 22430 14082 22482
rect 17166 22430 17218 22482
rect 17726 22430 17778 22482
rect 19854 22430 19906 22482
rect 20750 22430 20802 22482
rect 25902 22430 25954 22482
rect 26574 22430 26626 22482
rect 13582 22318 13634 22370
rect 13806 22318 13858 22370
rect 17614 22318 17666 22370
rect 18510 22318 18562 22370
rect 22094 22318 22146 22370
rect 23886 22318 23938 22370
rect 25006 22318 25058 22370
rect 25566 22318 25618 22370
rect 28590 22318 28642 22370
rect 14142 22206 14194 22258
rect 16046 22206 16098 22258
rect 16830 22206 16882 22258
rect 17950 22206 18002 22258
rect 20526 22206 20578 22258
rect 21422 22206 21474 22258
rect 22654 22206 22706 22258
rect 25678 22206 25730 22258
rect 28030 22206 28082 22258
rect 28478 22206 28530 22258
rect 16382 22094 16434 22146
rect 17054 22094 17106 22146
rect 17278 22094 17330 22146
rect 19294 22094 19346 22146
rect 21758 22094 21810 22146
rect 24446 22094 24498 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 16270 21758 16322 21810
rect 22990 21758 23042 21810
rect 23326 21758 23378 21810
rect 17614 21646 17666 21698
rect 27358 21646 27410 21698
rect 22654 21534 22706 21586
rect 28030 21534 28082 21586
rect 29374 21534 29426 21586
rect 37662 21534 37714 21586
rect 16830 21422 16882 21474
rect 25230 21422 25282 21474
rect 28926 21422 28978 21474
rect 28814 21310 28866 21362
rect 40014 21310 40066 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 16382 20974 16434 21026
rect 18622 20974 18674 21026
rect 19406 20974 19458 21026
rect 21870 20974 21922 21026
rect 19630 20862 19682 20914
rect 22878 20862 22930 20914
rect 27918 20862 27970 20914
rect 29262 20862 29314 20914
rect 39790 20862 39842 20914
rect 14478 20750 14530 20802
rect 14702 20750 14754 20802
rect 17502 20750 17554 20802
rect 18286 20750 18338 20802
rect 18734 20750 18786 20802
rect 19854 20750 19906 20802
rect 20078 20750 20130 20802
rect 21310 20750 21362 20802
rect 21534 20750 21586 20802
rect 22542 20750 22594 20802
rect 23326 20750 23378 20802
rect 29150 20750 29202 20802
rect 29822 20750 29874 20802
rect 37662 20750 37714 20802
rect 14030 20638 14082 20690
rect 16494 20638 16546 20690
rect 17614 20638 17666 20690
rect 30158 20638 30210 20690
rect 13918 20526 13970 20578
rect 14254 20526 14306 20578
rect 29374 20526 29426 20578
rect 29598 20526 29650 20578
rect 30270 20526 30322 20578
rect 30494 20526 30546 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 40238 20190 40290 20242
rect 16830 20078 16882 20130
rect 18734 20078 18786 20130
rect 19070 20078 19122 20130
rect 23326 20078 23378 20130
rect 27134 20078 27186 20130
rect 28590 20078 28642 20130
rect 11566 19966 11618 20018
rect 16494 19966 16546 20018
rect 17390 19966 17442 20018
rect 18398 19966 18450 20018
rect 19406 19966 19458 20018
rect 26910 19966 26962 20018
rect 27582 19966 27634 20018
rect 27806 19966 27858 20018
rect 12238 19854 12290 19906
rect 14366 19854 14418 19906
rect 14814 19854 14866 19906
rect 17950 19854 18002 19906
rect 27022 19854 27074 19906
rect 30718 19854 30770 19906
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 19630 19406 19682 19458
rect 21646 19406 21698 19458
rect 21870 19406 21922 19458
rect 26910 19406 26962 19458
rect 27134 19406 27186 19458
rect 20750 19294 20802 19346
rect 21422 19294 21474 19346
rect 14142 19182 14194 19234
rect 14366 19182 14418 19234
rect 16494 19182 16546 19234
rect 18286 19182 18338 19234
rect 18958 19182 19010 19234
rect 20302 19182 20354 19234
rect 23214 19182 23266 19234
rect 23662 19182 23714 19234
rect 12574 19070 12626 19122
rect 12910 19070 12962 19122
rect 13470 19070 13522 19122
rect 16046 19070 16098 19122
rect 16830 19070 16882 19122
rect 18174 19070 18226 19122
rect 22990 19070 23042 19122
rect 16158 18958 16210 19010
rect 17166 18958 17218 19010
rect 17502 18958 17554 19010
rect 17950 18958 18002 19010
rect 18622 18958 18674 19010
rect 19406 18958 19458 19010
rect 19518 18958 19570 19010
rect 22318 18958 22370 19010
rect 23774 18958 23826 19010
rect 23998 18958 24050 19010
rect 26910 18958 26962 19010
rect 27470 18958 27522 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 19182 18622 19234 18674
rect 19630 18622 19682 18674
rect 21086 18622 21138 18674
rect 22206 18622 22258 18674
rect 25566 18622 25618 18674
rect 18846 18510 18898 18562
rect 20414 18510 20466 18562
rect 21982 18510 22034 18562
rect 22654 18510 22706 18562
rect 22766 18510 22818 18562
rect 28030 18510 28082 18562
rect 12798 18398 12850 18450
rect 13582 18398 13634 18450
rect 16158 18398 16210 18450
rect 18622 18398 18674 18450
rect 19070 18398 19122 18450
rect 19854 18398 19906 18450
rect 20750 18398 20802 18450
rect 22094 18398 22146 18450
rect 25230 18398 25282 18450
rect 25454 18398 25506 18450
rect 25902 18398 25954 18450
rect 26126 18398 26178 18450
rect 27246 18398 27298 18450
rect 37662 18398 37714 18450
rect 15710 18286 15762 18338
rect 18958 18286 19010 18338
rect 21422 18286 21474 18338
rect 21646 18286 21698 18338
rect 25678 18286 25730 18338
rect 26910 18286 26962 18338
rect 30158 18286 30210 18338
rect 22766 18174 22818 18226
rect 26798 18174 26850 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 28254 17838 28306 17890
rect 1934 17726 1986 17778
rect 25678 17726 25730 17778
rect 27806 17726 27858 17778
rect 40014 17726 40066 17778
rect 4286 17614 4338 17666
rect 14814 17614 14866 17666
rect 21646 17614 21698 17666
rect 25006 17614 25058 17666
rect 37662 17614 37714 17666
rect 14142 17502 14194 17554
rect 14254 17502 14306 17554
rect 14702 17502 14754 17554
rect 20078 17502 20130 17554
rect 28142 17502 28194 17554
rect 28254 17502 28306 17554
rect 13918 17390 13970 17442
rect 14478 17390 14530 17442
rect 20190 17390 20242 17442
rect 20414 17390 20466 17442
rect 21310 17390 21362 17442
rect 29262 17390 29314 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 15598 17054 15650 17106
rect 23102 17054 23154 17106
rect 24446 17054 24498 17106
rect 18958 16942 19010 16994
rect 19294 16942 19346 16994
rect 22206 16942 22258 16994
rect 22430 16942 22482 16994
rect 23326 16942 23378 16994
rect 23438 16942 23490 16994
rect 24110 16942 24162 16994
rect 30046 16942 30098 16994
rect 4286 16830 4338 16882
rect 13470 16830 13522 16882
rect 14142 16830 14194 16882
rect 14478 16830 14530 16882
rect 14702 16830 14754 16882
rect 14814 16830 14866 16882
rect 15150 16830 15202 16882
rect 22766 16830 22818 16882
rect 24446 16830 24498 16882
rect 24782 16830 24834 16882
rect 26686 16830 26738 16882
rect 37886 16830 37938 16882
rect 11342 16718 11394 16770
rect 21982 16718 22034 16770
rect 27470 16718 27522 16770
rect 29598 16718 29650 16770
rect 40014 16718 40066 16770
rect 1934 16606 1986 16658
rect 22990 16606 23042 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 14814 16270 14866 16322
rect 19518 16270 19570 16322
rect 24222 16158 24274 16210
rect 26350 16158 26402 16210
rect 27358 16158 27410 16210
rect 40014 16158 40066 16210
rect 13806 16046 13858 16098
rect 14030 16046 14082 16098
rect 14366 16046 14418 16098
rect 14702 16046 14754 16098
rect 18734 16046 18786 16098
rect 19854 16046 19906 16098
rect 23550 16046 23602 16098
rect 26910 16046 26962 16098
rect 27582 16046 27634 16098
rect 29262 16046 29314 16098
rect 37662 16046 37714 16098
rect 14814 15934 14866 15986
rect 17950 15934 18002 15986
rect 27134 15934 27186 15986
rect 13918 15822 13970 15874
rect 17614 15822 17666 15874
rect 17838 15822 17890 15874
rect 18398 15822 18450 15874
rect 19182 15822 19234 15874
rect 19630 15822 19682 15874
rect 29486 15822 29538 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 14702 15486 14754 15538
rect 16606 15486 16658 15538
rect 18510 15486 18562 15538
rect 18846 15486 18898 15538
rect 20414 15486 20466 15538
rect 20862 15486 20914 15538
rect 23886 15486 23938 15538
rect 25118 15486 25170 15538
rect 26574 15486 26626 15538
rect 13470 15374 13522 15426
rect 17502 15374 17554 15426
rect 17726 15374 17778 15426
rect 20638 15374 20690 15426
rect 22766 15374 22818 15426
rect 25342 15374 25394 15426
rect 25454 15374 25506 15426
rect 14254 15262 14306 15314
rect 16270 15262 16322 15314
rect 16606 15262 16658 15314
rect 16942 15262 16994 15314
rect 17950 15262 18002 15314
rect 18174 15262 18226 15314
rect 18622 15262 18674 15314
rect 18734 15262 18786 15314
rect 19070 15262 19122 15314
rect 19294 15262 19346 15314
rect 19630 15262 19682 15314
rect 19854 15262 19906 15314
rect 20078 15262 20130 15314
rect 20302 15262 20354 15314
rect 22990 15262 23042 15314
rect 11342 15150 11394 15202
rect 23998 15150 24050 15202
rect 20974 15038 21026 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 17054 14590 17106 14642
rect 19182 14590 19234 14642
rect 22766 14590 22818 14642
rect 24894 14590 24946 14642
rect 25342 14590 25394 14642
rect 16270 14478 16322 14530
rect 19630 14478 19682 14530
rect 22094 14478 22146 14530
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 21086 13806 21138 13858
rect 21870 13694 21922 13746
rect 22318 13694 22370 13746
rect 18958 13582 19010 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 15598 13022 15650 13074
rect 17726 13022 17778 13074
rect 18286 13022 18338 13074
rect 14814 12910 14866 12962
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 18398 4398 18450 4450
rect 19070 4286 19122 4338
rect 20078 4062 20130 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18622 3614 18674 3666
rect 22094 3614 22146 3666
rect 25566 3614 25618 3666
rect 17614 3502 17666 3554
rect 21086 3502 21138 3554
rect 24558 3502 24610 3554
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 18144 41200 18256 42000
rect 18816 41200 18928 42000
rect 20160 41200 20272 42000
rect 22176 41200 22288 42000
rect 24864 41200 24976 42000
rect 25536 41200 25648 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 18060 38050 18116 38062
rect 18060 37998 18062 38050
rect 18114 37998 18116 38050
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 18060 31948 18116 37998
rect 18172 37380 18228 41200
rect 18844 38162 18900 41200
rect 18844 38110 18846 38162
rect 18898 38110 18900 38162
rect 18844 38098 18900 38110
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20188 37492 20244 41200
rect 22204 38276 22260 41200
rect 22428 38276 22484 38286
rect 22204 38274 22484 38276
rect 22204 38222 22430 38274
rect 22482 38222 22484 38274
rect 22204 38220 22484 38222
rect 22428 38210 22484 38220
rect 24892 38276 24948 41200
rect 24892 38210 24948 38220
rect 21532 38050 21588 38062
rect 21532 37998 21534 38050
rect 21586 37998 21588 38050
rect 20188 37426 20244 37436
rect 21420 37492 21476 37502
rect 21420 37398 21476 37436
rect 18284 37380 18340 37390
rect 18172 37378 18340 37380
rect 18172 37326 18286 37378
rect 18338 37326 18340 37378
rect 18172 37324 18340 37326
rect 18284 37314 18340 37324
rect 19628 37266 19684 37278
rect 19628 37214 19630 37266
rect 19682 37214 19684 37266
rect 19628 31948 19684 37214
rect 20524 37266 20580 37278
rect 20524 37214 20526 37266
rect 20578 37214 20580 37266
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 18060 31892 18340 31948
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 17612 27858 17668 27870
rect 17612 27806 17614 27858
rect 17666 27806 17668 27858
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 15708 27076 15764 27086
rect 15708 26982 15764 27020
rect 16380 27076 16436 27086
rect 4172 26964 4228 26974
rect 1932 25618 1988 25630
rect 1932 25566 1934 25618
rect 1986 25566 1988 25618
rect 1932 24948 1988 25566
rect 1932 24882 1988 24892
rect 1932 24500 1988 24510
rect 1932 24406 1988 24444
rect 1932 22932 1988 22942
rect 1932 22838 1988 22876
rect 4172 19908 4228 26908
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 13468 25618 13524 25630
rect 13468 25566 13470 25618
rect 13522 25566 13524 25618
rect 4284 25508 4340 25518
rect 4284 25414 4340 25452
rect 13468 25508 13524 25566
rect 13468 25442 13524 25452
rect 15260 25508 15316 25518
rect 15260 24834 15316 25452
rect 16268 25506 16324 25518
rect 16268 25454 16270 25506
rect 16322 25454 16324 25506
rect 15596 25396 15652 25406
rect 15596 25394 16100 25396
rect 15596 25342 15598 25394
rect 15650 25342 16100 25394
rect 15596 25340 16100 25342
rect 15596 25330 15652 25340
rect 16044 24946 16100 25340
rect 16268 25284 16324 25454
rect 16380 25284 16436 27020
rect 17612 27076 17668 27806
rect 17612 27010 17668 27020
rect 16492 26962 16548 26974
rect 16492 26910 16494 26962
rect 16546 26910 16548 26962
rect 16492 26516 16548 26910
rect 16492 26450 16548 26460
rect 17388 26516 17444 26526
rect 18284 26516 18340 31892
rect 19516 31892 19684 31948
rect 18396 27748 18452 27758
rect 18396 27746 18900 27748
rect 18396 27694 18398 27746
rect 18450 27694 18900 27746
rect 18396 27692 18900 27694
rect 18396 27682 18452 27692
rect 18732 27524 18788 27534
rect 18620 27468 18732 27524
rect 18620 27186 18676 27468
rect 18732 27458 18788 27468
rect 18620 27134 18622 27186
rect 18674 27134 18676 27186
rect 18620 26908 18676 27134
rect 18844 27074 18900 27692
rect 19516 27524 19572 31892
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19516 27458 19572 27468
rect 19628 27748 19684 27758
rect 20524 27748 20580 37214
rect 19404 27300 19460 27310
rect 19180 27298 19460 27300
rect 19180 27246 19406 27298
rect 19458 27246 19460 27298
rect 19180 27244 19460 27246
rect 18844 27022 18846 27074
rect 18898 27022 18900 27074
rect 18844 27010 18900 27022
rect 18956 27076 19012 27086
rect 18620 26852 18788 26908
rect 18396 26516 18452 26526
rect 18284 26514 18452 26516
rect 18284 26462 18398 26514
rect 18450 26462 18452 26514
rect 18284 26460 18452 26462
rect 17388 26422 17444 26460
rect 18396 26450 18452 26460
rect 18508 26404 18564 26414
rect 17724 26290 17780 26302
rect 17724 26238 17726 26290
rect 17778 26238 17780 26290
rect 16828 25284 16884 25294
rect 16268 25282 16884 25284
rect 16268 25230 16830 25282
rect 16882 25230 16884 25282
rect 16268 25228 16884 25230
rect 16044 24894 16046 24946
rect 16098 24894 16100 24946
rect 16044 24882 16100 24894
rect 16156 24948 16212 24958
rect 16156 24854 16212 24892
rect 15260 24782 15262 24834
rect 15314 24782 15316 24834
rect 15260 24770 15316 24782
rect 4284 24722 4340 24734
rect 4284 24670 4286 24722
rect 4338 24670 4340 24722
rect 4284 24612 4340 24670
rect 4284 24546 4340 24556
rect 11564 24722 11620 24734
rect 11564 24670 11566 24722
rect 11618 24670 11620 24722
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 11564 23604 11620 24670
rect 14700 24724 14756 24734
rect 12236 24612 12292 24622
rect 14364 24612 14420 24622
rect 12236 24610 12628 24612
rect 12236 24558 12238 24610
rect 12290 24558 12628 24610
rect 12236 24556 12628 24558
rect 12236 24546 12292 24556
rect 12572 24162 12628 24556
rect 12572 24110 12574 24162
rect 12626 24110 12628 24162
rect 12572 24098 12628 24110
rect 14252 24556 14364 24612
rect 14028 24052 14084 24062
rect 14028 23938 14084 23996
rect 14028 23886 14030 23938
rect 14082 23886 14084 23938
rect 14028 23874 14084 23886
rect 14252 23938 14308 24556
rect 14364 24518 14420 24556
rect 14476 24052 14532 24062
rect 14532 23996 14644 24052
rect 14476 23986 14532 23996
rect 14252 23886 14254 23938
rect 14306 23886 14308 23938
rect 14252 23874 14308 23886
rect 12908 23828 12964 23838
rect 12908 23734 12964 23772
rect 14140 23828 14196 23838
rect 14140 23734 14196 23772
rect 11564 23538 11620 23548
rect 12684 23714 12740 23726
rect 12684 23662 12686 23714
rect 12738 23662 12740 23714
rect 4284 23156 4340 23166
rect 4284 23062 4340 23100
rect 10892 23044 10948 23054
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 10892 22372 10948 22988
rect 12684 22932 12740 23662
rect 13804 23604 13860 23614
rect 13804 23154 13860 23548
rect 13804 23102 13806 23154
rect 13858 23102 13860 23154
rect 13804 23090 13860 23102
rect 14476 23156 14532 23166
rect 14476 23062 14532 23100
rect 13020 23044 13076 23054
rect 13020 22950 13076 22988
rect 14252 23044 14308 23054
rect 14252 22950 14308 22988
rect 12684 22866 12740 22876
rect 13580 22932 13636 22942
rect 10892 22306 10948 22316
rect 13580 22484 13636 22876
rect 14140 22930 14196 22942
rect 14140 22878 14142 22930
rect 14194 22878 14196 22930
rect 13580 22370 13636 22428
rect 14028 22484 14084 22494
rect 14140 22484 14196 22878
rect 14028 22482 14196 22484
rect 14028 22430 14030 22482
rect 14082 22430 14196 22482
rect 14028 22428 14196 22430
rect 14028 22418 14084 22428
rect 13580 22318 13582 22370
rect 13634 22318 13636 22370
rect 13580 22306 13636 22318
rect 13804 22372 13860 22382
rect 13804 22278 13860 22316
rect 14140 22258 14196 22270
rect 14140 22206 14142 22258
rect 14194 22206 14196 22258
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 13692 20748 14084 20804
rect 4172 19842 4228 19852
rect 11564 20018 11620 20030
rect 11564 19966 11566 20018
rect 11618 19966 11620 20018
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 11564 18452 11620 19966
rect 12236 19908 12292 19918
rect 12236 19906 12628 19908
rect 12236 19854 12238 19906
rect 12290 19854 12628 19906
rect 12236 19852 12628 19854
rect 12236 19842 12292 19852
rect 12572 19122 12628 19852
rect 12572 19070 12574 19122
rect 12626 19070 12628 19122
rect 12572 19058 12628 19070
rect 12908 19124 12964 19134
rect 13468 19124 13524 19134
rect 12908 19122 13524 19124
rect 12908 19070 12910 19122
rect 12962 19070 13470 19122
rect 13522 19070 13524 19122
rect 12908 19068 13524 19070
rect 12908 19058 12964 19068
rect 13468 19058 13524 19068
rect 11564 18386 11620 18396
rect 12796 18452 12852 18462
rect 12796 18358 12852 18396
rect 13580 18452 13636 18462
rect 13692 18452 13748 20748
rect 14028 20690 14084 20748
rect 14028 20638 14030 20690
rect 14082 20638 14084 20690
rect 14028 20626 14084 20638
rect 13916 20578 13972 20590
rect 13916 20526 13918 20578
rect 13970 20526 13972 20578
rect 13916 20188 13972 20526
rect 14140 20188 14196 22206
rect 14476 20804 14532 20814
rect 14588 20804 14644 23996
rect 14476 20802 14644 20804
rect 14476 20750 14478 20802
rect 14530 20750 14644 20802
rect 14476 20748 14644 20750
rect 14700 23938 14756 24668
rect 15036 24722 15092 24734
rect 15036 24670 15038 24722
rect 15090 24670 15092 24722
rect 15036 24052 15092 24670
rect 15596 24724 15652 24734
rect 16268 24724 16324 25228
rect 16828 25218 16884 25228
rect 15596 24630 15652 24668
rect 16156 24668 16324 24724
rect 17052 24948 17108 24958
rect 15484 24610 15540 24622
rect 15484 24558 15486 24610
rect 15538 24558 15540 24610
rect 15484 24500 15540 24558
rect 15932 24500 15988 24510
rect 15484 24498 15988 24500
rect 15484 24446 15934 24498
rect 15986 24446 15988 24498
rect 15484 24444 15988 24446
rect 15932 24434 15988 24444
rect 15036 23986 15092 23996
rect 14700 23886 14702 23938
rect 14754 23886 14756 23938
rect 14700 22148 14756 23886
rect 15036 23716 15092 23726
rect 14700 20802 14756 22092
rect 14700 20750 14702 20802
rect 14754 20750 14756 20802
rect 14476 20738 14532 20748
rect 14700 20738 14756 20750
rect 14924 23714 15092 23716
rect 14924 23662 15038 23714
rect 15090 23662 15092 23714
rect 14924 23660 15092 23662
rect 14924 23604 14980 23660
rect 15036 23650 15092 23660
rect 14924 23042 14980 23548
rect 16156 23604 16212 24668
rect 17052 23940 17108 24892
rect 17724 24164 17780 26238
rect 17836 24164 17892 24174
rect 17724 24162 17892 24164
rect 17724 24110 17838 24162
rect 17890 24110 17892 24162
rect 17724 24108 17892 24110
rect 17836 24098 17892 24108
rect 18060 24164 18116 24174
rect 17276 23940 17332 23950
rect 17052 23938 17220 23940
rect 17052 23886 17054 23938
rect 17106 23886 17220 23938
rect 17052 23884 17220 23886
rect 17052 23874 17108 23884
rect 16156 23538 16212 23548
rect 16940 23604 16996 23614
rect 16940 23378 16996 23548
rect 16940 23326 16942 23378
rect 16994 23326 16996 23378
rect 16940 23314 16996 23326
rect 14924 22990 14926 23042
rect 14978 22990 14980 23042
rect 14924 21700 14980 22990
rect 17052 22932 17108 22942
rect 16940 22876 17052 22932
rect 16828 22820 16884 22830
rect 16380 22372 16436 22382
rect 16268 22316 16380 22372
rect 16044 22260 16100 22270
rect 16044 22166 16100 22204
rect 16268 21812 16324 22316
rect 16380 22306 16436 22316
rect 16828 22258 16884 22764
rect 16828 22206 16830 22258
rect 16882 22206 16884 22258
rect 16828 22194 16884 22206
rect 16380 22148 16436 22158
rect 16380 22054 16436 22092
rect 16268 21810 16436 21812
rect 16268 21758 16270 21810
rect 16322 21758 16436 21810
rect 16268 21756 16436 21758
rect 16268 21746 16324 21756
rect 13580 18450 13748 18452
rect 13580 18398 13582 18450
rect 13634 18398 13748 18450
rect 13580 18396 13748 18398
rect 13580 18386 13636 18396
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1932 17778 1988 17790
rect 1932 17726 1934 17778
rect 1986 17726 1988 17778
rect 1932 16884 1988 17726
rect 4284 17668 4340 17678
rect 4284 17574 4340 17612
rect 11228 17668 11284 17678
rect 1932 16818 1988 16828
rect 4284 16882 4340 16894
rect 4284 16830 4286 16882
rect 4338 16830 4340 16882
rect 4284 16772 4340 16830
rect 4284 16706 4340 16716
rect 1932 16658 1988 16670
rect 1932 16606 1934 16658
rect 1986 16606 1988 16658
rect 1932 16212 1988 16606
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 1932 16146 1988 16156
rect 11228 15204 11284 17612
rect 13692 17556 13748 18396
rect 13692 17490 13748 17500
rect 13804 20132 13972 20188
rect 14028 20132 14196 20188
rect 14252 20578 14308 20590
rect 14252 20526 14254 20578
rect 14306 20526 14308 20578
rect 13468 16884 13524 16894
rect 13468 16790 13524 16828
rect 11340 16772 11396 16782
rect 11340 15988 11396 16716
rect 13804 16098 13860 20132
rect 14028 18788 14084 20132
rect 14140 19234 14196 19246
rect 14140 19182 14142 19234
rect 14194 19182 14196 19234
rect 14140 19012 14196 19182
rect 14252 19236 14308 20526
rect 14364 20020 14420 20030
rect 14364 19906 14420 19964
rect 14364 19854 14366 19906
rect 14418 19854 14420 19906
rect 14364 19842 14420 19854
rect 14812 19908 14868 19918
rect 14924 19908 14980 21644
rect 16380 21026 16436 21756
rect 16380 20974 16382 21026
rect 16434 20974 16436 21026
rect 16380 20962 16436 20974
rect 16828 21474 16884 21486
rect 16828 21422 16830 21474
rect 16882 21422 16884 21474
rect 16828 20804 16884 21422
rect 16828 20738 16884 20748
rect 16492 20690 16548 20702
rect 16492 20638 16494 20690
rect 16546 20638 16548 20690
rect 16492 20020 16548 20638
rect 16828 20132 16884 20142
rect 16828 20038 16884 20076
rect 16492 19926 16548 19964
rect 14812 19906 14980 19908
rect 14812 19854 14814 19906
rect 14866 19854 14980 19906
rect 14812 19852 14980 19854
rect 14364 19236 14420 19246
rect 14252 19234 14420 19236
rect 14252 19182 14366 19234
rect 14418 19182 14420 19234
rect 14252 19180 14420 19182
rect 14364 19124 14420 19180
rect 14364 19058 14420 19068
rect 14140 18946 14196 18956
rect 14028 18732 14196 18788
rect 14028 18452 14084 18462
rect 13804 16046 13806 16098
rect 13858 16046 13860 16098
rect 13804 16034 13860 16046
rect 13916 17442 13972 17454
rect 13916 17390 13918 17442
rect 13970 17390 13972 17442
rect 13916 16100 13972 17390
rect 14028 16884 14084 18396
rect 14140 17892 14196 18732
rect 14812 18452 14868 19852
rect 16828 19348 16884 19358
rect 16492 19236 16548 19246
rect 16044 19234 16548 19236
rect 16044 19182 16494 19234
rect 16546 19182 16548 19234
rect 16044 19180 16548 19182
rect 16044 19122 16100 19180
rect 16492 19170 16548 19180
rect 16044 19070 16046 19122
rect 16098 19070 16100 19122
rect 14812 18386 14868 18396
rect 14924 18564 14980 18574
rect 14140 17836 14308 17892
rect 14140 17668 14196 17678
rect 14140 17554 14196 17612
rect 14140 17502 14142 17554
rect 14194 17502 14196 17554
rect 14140 17490 14196 17502
rect 14252 17554 14308 17836
rect 14812 17668 14868 17678
rect 14924 17668 14980 18508
rect 14812 17666 14980 17668
rect 14812 17614 14814 17666
rect 14866 17614 14980 17666
rect 14812 17612 14980 17614
rect 15596 18452 15652 18462
rect 14812 17602 14868 17612
rect 14252 17502 14254 17554
rect 14306 17502 14308 17554
rect 14252 17444 14308 17502
rect 14700 17556 14756 17566
rect 14700 17462 14756 17500
rect 14252 17378 14308 17388
rect 14476 17442 14532 17454
rect 14476 17390 14478 17442
rect 14530 17390 14532 17442
rect 14140 16884 14196 16894
rect 14028 16882 14308 16884
rect 14028 16830 14142 16882
rect 14194 16830 14308 16882
rect 14028 16828 14308 16830
rect 14140 16818 14196 16828
rect 14028 16100 14084 16110
rect 13916 16098 14084 16100
rect 13916 16046 14030 16098
rect 14082 16046 14084 16098
rect 13916 16044 14084 16046
rect 14028 16034 14084 16044
rect 11340 15922 11396 15932
rect 13916 15874 13972 15886
rect 13916 15822 13918 15874
rect 13970 15822 13972 15874
rect 13916 15540 13972 15822
rect 13468 15484 13972 15540
rect 14252 15540 14308 16828
rect 14476 16882 14532 17390
rect 14476 16830 14478 16882
rect 14530 16830 14532 16882
rect 14476 16818 14532 16830
rect 14588 17444 14644 17454
rect 14364 16100 14420 16110
rect 14588 16100 14644 17388
rect 15596 17106 15652 18396
rect 15708 18340 15764 18350
rect 16044 18340 16100 19070
rect 16828 19122 16884 19292
rect 16828 19070 16830 19122
rect 16882 19070 16884 19122
rect 16828 19058 16884 19070
rect 16156 19012 16212 19022
rect 16156 18918 16212 18956
rect 16156 18452 16212 18462
rect 16156 18358 16212 18396
rect 15708 18338 16100 18340
rect 15708 18286 15710 18338
rect 15762 18286 16100 18338
rect 15708 18284 16100 18286
rect 15708 18274 15764 18284
rect 15596 17054 15598 17106
rect 15650 17054 15652 17106
rect 15596 17042 15652 17054
rect 14700 16884 14756 16894
rect 14700 16790 14756 16828
rect 14812 16882 14868 16894
rect 14812 16830 14814 16882
rect 14866 16830 14868 16882
rect 14812 16322 14868 16830
rect 14812 16270 14814 16322
rect 14866 16270 14868 16322
rect 14812 16258 14868 16270
rect 15148 16882 15204 16894
rect 15148 16830 15150 16882
rect 15202 16830 15204 16882
rect 14700 16100 14756 16110
rect 14588 16098 14756 16100
rect 14588 16046 14702 16098
rect 14754 16046 14756 16098
rect 14588 16044 14756 16046
rect 14364 16006 14420 16044
rect 14700 16034 14756 16044
rect 15148 16100 15204 16830
rect 14812 15988 14868 15998
rect 14812 15894 14868 15932
rect 14700 15540 14756 15550
rect 14252 15538 14756 15540
rect 14252 15486 14702 15538
rect 14754 15486 14756 15538
rect 14252 15484 14756 15486
rect 13468 15426 13524 15484
rect 13468 15374 13470 15426
rect 13522 15374 13524 15426
rect 13468 15362 13524 15374
rect 14252 15314 14308 15484
rect 14252 15262 14254 15314
rect 14306 15262 14308 15314
rect 14252 15250 14308 15262
rect 11340 15204 11396 15214
rect 11228 15202 11396 15204
rect 11228 15150 11342 15202
rect 11394 15150 11396 15202
rect 11228 15148 11396 15150
rect 11340 15138 11396 15148
rect 14700 15092 14756 15484
rect 15148 15316 15204 16044
rect 16604 15540 16660 15550
rect 15148 15250 15204 15260
rect 15596 15538 16660 15540
rect 15596 15486 16606 15538
rect 16658 15486 16660 15538
rect 15596 15484 16660 15486
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 14700 12964 14756 15036
rect 15596 13074 15652 15484
rect 16604 15474 16660 15484
rect 16268 15316 16324 15326
rect 16268 15222 16324 15260
rect 16604 15316 16660 15326
rect 16604 15222 16660 15260
rect 16940 15314 16996 22876
rect 17052 22866 17108 22876
rect 17164 22482 17220 23884
rect 17276 23846 17332 23884
rect 17500 23938 17556 23950
rect 17500 23886 17502 23938
rect 17554 23886 17556 23938
rect 17164 22430 17166 22482
rect 17218 22430 17220 22482
rect 17164 22418 17220 22430
rect 17388 23154 17444 23166
rect 17388 23102 17390 23154
rect 17442 23102 17444 23154
rect 17388 22260 17444 23102
rect 17500 23156 17556 23886
rect 17724 23938 17780 23950
rect 17724 23886 17726 23938
rect 17778 23886 17780 23938
rect 17724 23828 17780 23886
rect 17724 23762 17780 23772
rect 18060 23604 18116 24108
rect 17500 23062 17556 23100
rect 17612 23154 17668 23166
rect 17612 23102 17614 23154
rect 17666 23102 17668 23154
rect 17612 22596 17668 23102
rect 17388 22194 17444 22204
rect 17500 22540 17668 22596
rect 18060 23154 18116 23548
rect 18060 23102 18062 23154
rect 18114 23102 18116 23154
rect 17052 22146 17108 22158
rect 17052 22094 17054 22146
rect 17106 22094 17108 22146
rect 17052 19572 17108 22094
rect 17276 22146 17332 22158
rect 17276 22094 17278 22146
rect 17330 22094 17332 22146
rect 17276 22036 17332 22094
rect 17276 21970 17332 21980
rect 17500 21812 17556 22540
rect 17724 22484 17780 22522
rect 17724 22418 17780 22428
rect 17612 22372 17668 22382
rect 17612 22278 17668 22316
rect 17500 21476 17556 21756
rect 17948 22258 18004 22270
rect 17948 22206 17950 22258
rect 18002 22206 18004 22258
rect 17612 21700 17668 21710
rect 17612 21606 17668 21644
rect 17500 21420 17668 21476
rect 17500 20802 17556 20814
rect 17500 20750 17502 20802
rect 17554 20750 17556 20802
rect 17052 19506 17108 19516
rect 17388 20018 17444 20030
rect 17388 19966 17390 20018
rect 17442 19966 17444 20018
rect 17388 19460 17444 19966
rect 17388 19394 17444 19404
rect 17164 19010 17220 19022
rect 17164 18958 17166 19010
rect 17218 18958 17220 19010
rect 17164 18452 17220 18958
rect 17500 19012 17556 20750
rect 17612 20690 17668 21420
rect 17612 20638 17614 20690
rect 17666 20638 17668 20690
rect 17612 20626 17668 20638
rect 17948 20916 18004 22206
rect 18060 21588 18116 23102
rect 18284 23266 18340 23278
rect 18284 23214 18286 23266
rect 18338 23214 18340 23266
rect 18172 22932 18228 22942
rect 18172 22838 18228 22876
rect 18284 22820 18340 23214
rect 18508 23156 18564 26348
rect 18732 26290 18788 26852
rect 18732 26238 18734 26290
rect 18786 26238 18788 26290
rect 18620 24050 18676 24062
rect 18620 23998 18622 24050
rect 18674 23998 18676 24050
rect 18620 23940 18676 23998
rect 18732 23940 18788 26238
rect 18956 26180 19012 27020
rect 19180 27074 19236 27244
rect 19404 27234 19460 27244
rect 19180 27022 19182 27074
rect 19234 27022 19236 27074
rect 19180 27010 19236 27022
rect 19068 26962 19124 26974
rect 19068 26910 19070 26962
rect 19122 26910 19124 26962
rect 19068 26404 19124 26910
rect 19068 26338 19124 26348
rect 19628 26850 19684 27692
rect 20076 27746 20580 27748
rect 20076 27694 20526 27746
rect 20578 27694 20580 27746
rect 20076 27692 20580 27694
rect 19740 27298 19796 27310
rect 19740 27246 19742 27298
rect 19794 27246 19796 27298
rect 19740 27076 19796 27246
rect 19852 27076 19908 27086
rect 19740 27074 19908 27076
rect 19740 27022 19854 27074
rect 19906 27022 19908 27074
rect 19740 27020 19908 27022
rect 19852 27010 19908 27020
rect 20076 26962 20132 27692
rect 20524 27682 20580 27692
rect 20972 27748 21028 27758
rect 20972 27654 21028 27692
rect 20076 26910 20078 26962
rect 20130 26910 20132 26962
rect 20076 26898 20132 26910
rect 20188 26962 20244 26974
rect 20188 26910 20190 26962
rect 20242 26910 20244 26962
rect 19628 26798 19630 26850
rect 19682 26798 19684 26850
rect 19628 26290 19684 26798
rect 20188 26852 20244 26910
rect 20636 26962 20692 26974
rect 20636 26910 20638 26962
rect 20690 26910 20692 26962
rect 20188 26786 20244 26796
rect 20412 26850 20468 26862
rect 20412 26798 20414 26850
rect 20466 26798 20468 26850
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20300 26404 20356 26414
rect 20412 26404 20468 26798
rect 20300 26402 20468 26404
rect 20300 26350 20302 26402
rect 20354 26350 20468 26402
rect 20300 26348 20468 26350
rect 20300 26338 20356 26348
rect 19628 26238 19630 26290
rect 19682 26238 19684 26290
rect 19180 26180 19236 26190
rect 19628 26180 19684 26238
rect 18956 26178 19684 26180
rect 18956 26126 19182 26178
rect 19234 26126 19684 26178
rect 18956 26124 19684 26126
rect 19180 26114 19236 26124
rect 19292 25396 19348 25406
rect 19180 25340 19292 25396
rect 19068 23940 19124 23950
rect 18732 23938 19124 23940
rect 18732 23886 19070 23938
rect 19122 23886 19124 23938
rect 18732 23884 19124 23886
rect 18620 23874 18676 23884
rect 19068 23874 19124 23884
rect 18620 23714 18676 23726
rect 18620 23662 18622 23714
rect 18674 23662 18676 23714
rect 18620 23604 18676 23662
rect 18732 23716 18788 23726
rect 18956 23716 19012 23726
rect 18732 23714 18900 23716
rect 18732 23662 18734 23714
rect 18786 23662 18900 23714
rect 18732 23660 18900 23662
rect 18732 23650 18788 23660
rect 18620 23538 18676 23548
rect 18732 23156 18788 23166
rect 18508 23154 18676 23156
rect 18508 23102 18510 23154
rect 18562 23102 18676 23154
rect 18508 23100 18676 23102
rect 18508 23090 18564 23100
rect 18284 22754 18340 22764
rect 18508 22372 18564 22382
rect 18060 21532 18228 21588
rect 17948 19908 18004 20860
rect 17948 19906 18116 19908
rect 17948 19854 17950 19906
rect 18002 19854 18116 19906
rect 17948 19852 18116 19854
rect 17948 19842 18004 19852
rect 18060 19124 18116 19852
rect 18172 19796 18228 21532
rect 18284 20804 18340 20814
rect 18284 20710 18340 20748
rect 18396 20020 18452 20030
rect 18396 19926 18452 19964
rect 18172 19740 18452 19796
rect 18284 19236 18340 19246
rect 18284 19142 18340 19180
rect 18172 19124 18228 19134
rect 18060 19068 18172 19124
rect 18172 19030 18228 19068
rect 17500 18918 17556 18956
rect 17948 19010 18004 19022
rect 18396 19012 18452 19740
rect 17948 18958 17950 19010
rect 18002 18958 18004 19010
rect 17164 17556 17220 18396
rect 17948 18228 18004 18958
rect 17948 18162 18004 18172
rect 18284 18956 18452 19012
rect 17164 17490 17220 17500
rect 17948 15988 18004 15998
rect 17948 15986 18228 15988
rect 17948 15934 17950 15986
rect 18002 15934 18228 15986
rect 17948 15932 18228 15934
rect 17948 15922 18004 15932
rect 17612 15874 17668 15886
rect 17612 15822 17614 15874
rect 17666 15822 17668 15874
rect 17500 15428 17556 15438
rect 17500 15334 17556 15372
rect 16940 15262 16942 15314
rect 16994 15262 16996 15314
rect 16940 15250 16996 15262
rect 17612 15316 17668 15822
rect 17724 15876 17780 15886
rect 17724 15426 17780 15820
rect 17836 15874 17892 15886
rect 17836 15822 17838 15874
rect 17890 15822 17892 15874
rect 17836 15540 17892 15822
rect 18172 15540 18228 15932
rect 18284 15876 18340 18956
rect 18508 18004 18564 22316
rect 18620 21026 18676 23100
rect 18732 22484 18788 23100
rect 18732 22418 18788 22428
rect 18620 20974 18622 21026
rect 18674 20974 18676 21026
rect 18620 20962 18676 20974
rect 18732 22148 18788 22158
rect 18732 20802 18788 22092
rect 18732 20750 18734 20802
rect 18786 20750 18788 20802
rect 18732 20738 18788 20750
rect 18732 20132 18788 20142
rect 18732 20038 18788 20076
rect 18620 19460 18676 19470
rect 18620 19010 18676 19404
rect 18620 18958 18622 19010
rect 18674 18958 18676 19010
rect 18620 18676 18676 18958
rect 18844 18900 18900 23660
rect 18956 23622 19012 23660
rect 19068 22484 19124 22494
rect 18956 22428 19068 22484
rect 18956 20132 19012 22428
rect 19068 22418 19124 22428
rect 19180 22148 19236 25340
rect 19292 25330 19348 25340
rect 19628 24724 19684 26124
rect 20636 25620 20692 26910
rect 20748 26964 20804 26974
rect 21308 26964 21364 26974
rect 20748 26962 21364 26964
rect 20748 26910 20750 26962
rect 20802 26910 21310 26962
rect 21362 26910 21364 26962
rect 20748 26908 21364 26910
rect 20748 26898 20804 26908
rect 21308 26898 21364 26908
rect 21532 26964 21588 37998
rect 25228 38050 25284 38062
rect 25228 37998 25230 38050
rect 25282 37998 25284 38050
rect 25228 28532 25284 37998
rect 25564 37492 25620 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 26124 38276 26180 38286
rect 26124 38182 26180 38220
rect 25788 37492 25844 37502
rect 25564 37490 25844 37492
rect 25564 37438 25790 37490
rect 25842 37438 25844 37490
rect 25564 37436 25844 37438
rect 25788 37426 25844 37436
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 25116 28476 25284 28532
rect 24108 27188 24164 27198
rect 22316 27076 22372 27086
rect 22316 26982 22372 27020
rect 21532 26870 21588 26908
rect 21644 26962 21700 26974
rect 21644 26910 21646 26962
rect 21698 26910 21700 26962
rect 21644 26852 21700 26910
rect 21644 26786 21700 26796
rect 22428 26964 22484 26974
rect 22428 26178 22484 26908
rect 22988 26964 23044 26974
rect 22988 26962 23268 26964
rect 22988 26910 22990 26962
rect 23042 26910 23268 26962
rect 22988 26908 23268 26910
rect 22988 26898 23044 26908
rect 23212 26514 23268 26908
rect 23212 26462 23214 26514
rect 23266 26462 23268 26514
rect 23212 26450 23268 26462
rect 24108 26514 24164 27132
rect 25116 27188 25172 28476
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 25564 27300 25620 27310
rect 25564 27298 26068 27300
rect 25564 27246 25566 27298
rect 25618 27246 26068 27298
rect 25564 27244 26068 27246
rect 25564 27234 25620 27244
rect 25116 27094 25172 27132
rect 25228 27076 25284 27086
rect 24108 26462 24110 26514
rect 24162 26462 24164 26514
rect 24108 26450 24164 26462
rect 24220 26852 24276 26862
rect 22428 26126 22430 26178
rect 22482 26126 22484 26178
rect 22428 26114 22484 26126
rect 23436 26402 23492 26414
rect 23436 26350 23438 26402
rect 23490 26350 23492 26402
rect 20412 25564 20692 25620
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20412 24948 20468 25564
rect 20524 25396 20580 25406
rect 20524 25302 20580 25340
rect 20076 24892 20468 24948
rect 20636 25282 20692 25294
rect 20636 25230 20638 25282
rect 20690 25230 20692 25282
rect 19964 24724 20020 24734
rect 19628 24722 20020 24724
rect 19628 24670 19630 24722
rect 19682 24670 19966 24722
rect 20018 24670 20020 24722
rect 19628 24668 20020 24670
rect 19628 24658 19684 24668
rect 19964 24658 20020 24668
rect 19740 23940 19796 23950
rect 19628 23938 19796 23940
rect 19628 23886 19742 23938
rect 19794 23886 19796 23938
rect 19628 23884 19796 23886
rect 19404 23828 19460 23838
rect 19292 23156 19348 23166
rect 19292 23062 19348 23100
rect 19292 22148 19348 22158
rect 19180 22092 19292 22148
rect 19292 22054 19348 22092
rect 19404 21026 19460 23772
rect 19404 20974 19406 21026
rect 19458 20974 19460 21026
rect 19404 20962 19460 20974
rect 19516 23714 19572 23726
rect 19516 23662 19518 23714
rect 19570 23662 19572 23714
rect 19516 23604 19572 23662
rect 19516 23042 19572 23548
rect 19516 22990 19518 23042
rect 19570 22990 19572 23042
rect 19516 20244 19572 22990
rect 19628 22596 19684 23884
rect 19740 23874 19796 23884
rect 20076 23716 20132 24892
rect 20636 24164 20692 25230
rect 20860 25284 20916 25294
rect 20860 25190 20916 25228
rect 22204 25282 22260 25294
rect 22204 25230 22206 25282
rect 22258 25230 22260 25282
rect 20748 24612 20804 24622
rect 20748 24610 21812 24612
rect 20748 24558 20750 24610
rect 20802 24558 21812 24610
rect 20748 24556 21812 24558
rect 20748 24546 20804 24556
rect 20076 23650 20132 23660
rect 20188 24108 20692 24164
rect 21196 24164 21252 24174
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19628 22502 19684 22540
rect 19852 23268 19908 23278
rect 19852 22484 19908 23212
rect 19852 22390 19908 22428
rect 20188 23154 20244 24108
rect 20636 23940 20692 23950
rect 20412 23716 20468 23726
rect 20188 23102 20190 23154
rect 20242 23102 20244 23154
rect 19628 22148 19684 22158
rect 19628 20914 19684 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20076 21588 20132 21598
rect 19628 20862 19630 20914
rect 19682 20862 19684 20914
rect 19628 20850 19684 20862
rect 19740 20916 19796 20926
rect 19796 20860 19908 20916
rect 19740 20850 19796 20860
rect 19852 20802 19908 20860
rect 19852 20750 19854 20802
rect 19906 20750 19908 20802
rect 19852 20738 19908 20750
rect 20076 20804 20132 21532
rect 20076 20710 20132 20748
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19292 20188 19572 20244
rect 19068 20132 19124 20142
rect 18956 20130 19124 20132
rect 18956 20078 19070 20130
rect 19122 20078 19124 20130
rect 18956 20076 19124 20078
rect 18956 19236 19012 20076
rect 19068 20066 19124 20076
rect 18956 19142 19012 19180
rect 18620 18610 18676 18620
rect 18732 18844 18844 18900
rect 18620 18452 18676 18462
rect 18620 18358 18676 18396
rect 18732 18228 18788 18844
rect 18844 18834 18900 18844
rect 19180 18900 19236 18910
rect 19180 18674 19236 18844
rect 19292 18788 19348 20188
rect 19628 20132 19684 20142
rect 19404 20020 19460 20030
rect 19404 19926 19460 19964
rect 19628 19460 19684 20076
rect 20188 20132 20244 23102
rect 20300 23714 20468 23716
rect 20300 23662 20414 23714
rect 20466 23662 20468 23714
rect 20300 23660 20468 23662
rect 20300 22372 20356 23660
rect 20412 23650 20468 23660
rect 20524 23492 20580 23502
rect 20524 23266 20580 23436
rect 20524 23214 20526 23266
rect 20578 23214 20580 23266
rect 20524 23202 20580 23214
rect 20412 23042 20468 23054
rect 20412 22990 20414 23042
rect 20466 22990 20468 23042
rect 20412 22820 20468 22990
rect 20412 22754 20468 22764
rect 20412 22596 20468 22606
rect 20412 22502 20468 22540
rect 20300 22306 20356 22316
rect 20524 22260 20580 22270
rect 20636 22260 20692 23884
rect 21196 23938 21252 24108
rect 21644 24052 21700 24062
rect 21644 23940 21700 23996
rect 21756 24050 21812 24556
rect 22204 24164 22260 25230
rect 23436 25284 23492 26350
rect 24220 26402 24276 26796
rect 24220 26350 24222 26402
rect 24274 26350 24276 26402
rect 24220 26338 24276 26350
rect 25004 26852 25060 26862
rect 23548 26292 23604 26302
rect 23884 26292 23940 26302
rect 23548 26290 23940 26292
rect 23548 26238 23550 26290
rect 23602 26238 23886 26290
rect 23938 26238 23940 26290
rect 23548 26236 23940 26238
rect 23548 26226 23604 26236
rect 23884 26226 23940 26236
rect 25004 25508 25060 26796
rect 25228 26290 25284 27020
rect 25564 26964 25620 26974
rect 25228 26238 25230 26290
rect 25282 26238 25284 26290
rect 25228 26226 25284 26238
rect 25452 26962 25620 26964
rect 25452 26910 25566 26962
rect 25618 26910 25620 26962
rect 25452 26908 25620 26910
rect 25004 25394 25060 25452
rect 25004 25342 25006 25394
rect 25058 25342 25060 25394
rect 25004 25330 25060 25342
rect 25228 25506 25284 25518
rect 25228 25454 25230 25506
rect 25282 25454 25284 25506
rect 23492 25228 24052 25284
rect 23436 25190 23492 25228
rect 22204 24098 22260 24108
rect 22876 24610 22932 24622
rect 22876 24558 22878 24610
rect 22930 24558 22932 24610
rect 21756 23998 21758 24050
rect 21810 23998 21812 24050
rect 21756 23986 21812 23998
rect 21196 23886 21198 23938
rect 21250 23886 21252 23938
rect 21196 23874 21252 23886
rect 21532 23938 21700 23940
rect 21532 23886 21646 23938
rect 21698 23886 21700 23938
rect 21532 23884 21700 23886
rect 20972 23716 21028 23726
rect 20748 22484 20804 22494
rect 20748 22390 20804 22428
rect 20524 22258 20692 22260
rect 20524 22206 20526 22258
rect 20578 22206 20692 22258
rect 20524 22204 20692 22206
rect 20524 22194 20580 22204
rect 20188 20066 20244 20076
rect 20748 20132 20804 20142
rect 19628 19366 19684 19404
rect 20300 19348 20356 19358
rect 20300 19234 20356 19292
rect 20748 19346 20804 20076
rect 20748 19294 20750 19346
rect 20802 19294 20804 19346
rect 20748 19282 20804 19294
rect 20300 19182 20302 19234
rect 20354 19182 20356 19234
rect 20300 19170 20356 19182
rect 19404 19012 19460 19022
rect 19404 18918 19460 18956
rect 19516 19010 19572 19022
rect 19516 18958 19518 19010
rect 19570 18958 19572 19010
rect 19292 18732 19460 18788
rect 19180 18622 19182 18674
rect 19234 18622 19236 18674
rect 19180 18610 19236 18622
rect 18844 18564 18900 18574
rect 18844 18470 18900 18508
rect 19068 18450 19124 18462
rect 19068 18398 19070 18450
rect 19122 18398 19124 18450
rect 18956 18338 19012 18350
rect 18956 18286 18958 18338
rect 19010 18286 19012 18338
rect 18732 18172 18900 18228
rect 18508 17938 18564 17948
rect 18732 16996 18788 17006
rect 18732 16098 18788 16940
rect 18732 16046 18734 16098
rect 18786 16046 18788 16098
rect 18732 16034 18788 16046
rect 18284 15810 18340 15820
rect 18396 15874 18452 15886
rect 18396 15822 18398 15874
rect 18450 15822 18452 15874
rect 18284 15540 18340 15550
rect 17836 15484 18116 15540
rect 18172 15484 18284 15540
rect 17724 15374 17726 15426
rect 17778 15374 17780 15426
rect 17724 15362 17780 15374
rect 17948 15316 18004 15326
rect 17612 15250 17668 15260
rect 17836 15314 18004 15316
rect 17836 15262 17950 15314
rect 18002 15262 18004 15314
rect 17836 15260 18004 15262
rect 16268 15092 16324 15102
rect 16268 14532 16324 15036
rect 17836 14868 17892 15260
rect 17948 15250 18004 15260
rect 18060 15148 18116 15484
rect 18284 15474 18340 15484
rect 18396 15428 18452 15822
rect 18508 15540 18564 15550
rect 18508 15446 18564 15484
rect 18844 15538 18900 18172
rect 18956 17332 19012 18286
rect 18956 17266 19012 17276
rect 18844 15486 18846 15538
rect 18898 15486 18900 15538
rect 18396 15362 18452 15372
rect 18844 15428 18900 15486
rect 18956 16994 19012 17006
rect 18956 16942 18958 16994
rect 19010 16942 19012 16994
rect 18956 15540 19012 16942
rect 19068 16996 19124 18398
rect 19292 18004 19348 18014
rect 19068 16930 19124 16940
rect 19180 17220 19236 17230
rect 19180 16100 19236 17164
rect 19292 16994 19348 17948
rect 19292 16942 19294 16994
rect 19346 16942 19348 16994
rect 19292 16930 19348 16942
rect 19180 16034 19236 16044
rect 19180 15876 19236 15886
rect 19180 15782 19236 15820
rect 18956 15474 19012 15484
rect 18844 15362 18900 15372
rect 18172 15316 18228 15326
rect 18172 15222 18228 15260
rect 18620 15314 18676 15326
rect 18620 15262 18622 15314
rect 18674 15262 18676 15314
rect 17052 14812 17892 14868
rect 17948 15092 18116 15148
rect 17052 14642 17108 14812
rect 17052 14590 17054 14642
rect 17106 14590 17108 14642
rect 17052 14578 17108 14590
rect 16268 14438 16324 14476
rect 17724 13076 17780 13086
rect 17948 13076 18004 15092
rect 18620 14644 18676 15262
rect 18732 15316 18788 15326
rect 18732 15222 18788 15260
rect 19068 15316 19124 15326
rect 19292 15316 19348 15326
rect 19404 15316 19460 18732
rect 19516 18340 19572 18958
rect 19628 18900 19684 18910
rect 19628 18674 19684 18844
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 18622 19630 18674
rect 19682 18622 19684 18674
rect 19628 18610 19684 18622
rect 20188 18676 20244 18686
rect 20972 18676 21028 23660
rect 21308 23268 21364 23278
rect 21308 23174 21364 23212
rect 21084 23154 21140 23166
rect 21084 23102 21086 23154
rect 21138 23102 21140 23154
rect 21084 22820 21140 23102
rect 21084 22754 21140 22764
rect 21420 23154 21476 23166
rect 21420 23102 21422 23154
rect 21474 23102 21476 23154
rect 21420 22596 21476 23102
rect 21420 22530 21476 22540
rect 21420 22260 21476 22270
rect 21532 22260 21588 23884
rect 21644 23874 21700 23884
rect 22540 23938 22596 23950
rect 22540 23886 22542 23938
rect 22594 23886 22596 23938
rect 22316 23826 22372 23838
rect 22316 23774 22318 23826
rect 22370 23774 22372 23826
rect 21868 23714 21924 23726
rect 21868 23662 21870 23714
rect 21922 23662 21924 23714
rect 21868 23156 21924 23662
rect 22204 23156 22260 23166
rect 21756 23044 21812 23054
rect 21420 22258 21588 22260
rect 21420 22206 21422 22258
rect 21474 22206 21588 22258
rect 21420 22204 21588 22206
rect 21644 23042 21812 23044
rect 21644 22990 21758 23042
rect 21810 22990 21812 23042
rect 21644 22988 21812 22990
rect 21644 22260 21700 22988
rect 21756 22978 21812 22988
rect 21420 22194 21476 22204
rect 21644 22194 21700 22204
rect 21756 22148 21812 22158
rect 21756 22054 21812 22092
rect 21868 21026 21924 23100
rect 21868 20974 21870 21026
rect 21922 20974 21924 21026
rect 21868 20962 21924 20974
rect 21980 23154 22260 23156
rect 21980 23102 22206 23154
rect 22258 23102 22260 23154
rect 21980 23100 22260 23102
rect 21308 20804 21364 20814
rect 21532 20804 21588 20814
rect 21308 20802 21476 20804
rect 21308 20750 21310 20802
rect 21362 20750 21476 20802
rect 21308 20748 21476 20750
rect 21308 20738 21364 20748
rect 21420 19348 21476 20748
rect 21532 20802 21700 20804
rect 21532 20750 21534 20802
rect 21586 20750 21700 20802
rect 21532 20748 21700 20750
rect 21532 20738 21588 20748
rect 21644 19460 21700 20748
rect 21980 20244 22036 23100
rect 22204 23090 22260 23100
rect 22092 22370 22148 22382
rect 22092 22318 22094 22370
rect 22146 22318 22148 22370
rect 22092 21812 22148 22318
rect 22316 22036 22372 23774
rect 22540 22260 22596 23886
rect 22876 23940 22932 24558
rect 23436 24164 23492 24174
rect 23492 24108 23604 24164
rect 23436 24098 23492 24108
rect 23436 23940 23492 23950
rect 22876 23874 22932 23884
rect 23100 23938 23492 23940
rect 23100 23886 23438 23938
rect 23490 23886 23492 23938
rect 23100 23884 23492 23886
rect 22988 23828 23044 23838
rect 23100 23828 23156 23884
rect 23436 23874 23492 23884
rect 22988 23826 23156 23828
rect 22988 23774 22990 23826
rect 23042 23774 23156 23826
rect 22988 23772 23156 23774
rect 22988 23762 23044 23772
rect 22988 23266 23044 23278
rect 22988 23214 22990 23266
rect 23042 23214 23044 23266
rect 22652 23156 22708 23166
rect 22652 23062 22708 23100
rect 22988 22596 23044 23214
rect 23100 23268 23156 23772
rect 23548 23378 23604 24108
rect 23660 24052 23716 24062
rect 23660 23958 23716 23996
rect 23548 23326 23550 23378
rect 23602 23326 23604 23378
rect 23212 23268 23268 23278
rect 23100 23266 23268 23268
rect 23100 23214 23214 23266
rect 23266 23214 23268 23266
rect 23100 23212 23268 23214
rect 22764 22540 23044 22596
rect 22652 22260 22708 22270
rect 22540 22204 22652 22260
rect 22652 22166 22708 22204
rect 22316 21970 22372 21980
rect 22092 21746 22148 21756
rect 22540 21924 22596 21934
rect 22540 20804 22596 21868
rect 21644 19366 21700 19404
rect 21868 19460 21924 19470
rect 21980 19460 22036 20188
rect 21868 19458 22036 19460
rect 21868 19406 21870 19458
rect 21922 19406 22036 19458
rect 21868 19404 22036 19406
rect 22204 20802 22596 20804
rect 22204 20750 22542 20802
rect 22594 20750 22596 20802
rect 22204 20748 22596 20750
rect 21868 19394 21924 19404
rect 21420 19254 21476 19292
rect 22092 19124 22148 19134
rect 21980 19068 22092 19124
rect 21084 18676 21140 18686
rect 20972 18674 21140 18676
rect 20972 18622 21086 18674
rect 21138 18622 21140 18674
rect 20972 18620 21140 18622
rect 19852 18564 19908 18574
rect 19852 18450 19908 18508
rect 19852 18398 19854 18450
rect 19906 18398 19908 18450
rect 19852 18340 19908 18398
rect 19516 18284 19908 18340
rect 19516 18116 19572 18126
rect 19516 16322 19572 18060
rect 20076 17556 20132 17566
rect 19628 17554 20132 17556
rect 19628 17502 20078 17554
rect 20130 17502 20132 17554
rect 19628 17500 20132 17502
rect 19628 16996 19684 17500
rect 20076 17490 20132 17500
rect 20188 17442 20244 18620
rect 21084 18610 21140 18620
rect 20412 18562 20468 18574
rect 20412 18510 20414 18562
rect 20466 18510 20468 18562
rect 20412 17668 20468 18510
rect 21980 18562 22036 19068
rect 22092 19058 22148 19068
rect 22204 18674 22260 20748
rect 22540 20738 22596 20748
rect 22652 21586 22708 21598
rect 22652 21534 22654 21586
rect 22706 21534 22708 21586
rect 22652 20804 22708 21534
rect 22652 20738 22708 20748
rect 22764 20692 22820 22540
rect 22988 22484 23044 22540
rect 22988 22418 23044 22428
rect 22876 22372 22932 22382
rect 22876 21812 22932 22316
rect 22876 20914 22932 21756
rect 22988 22148 23044 22158
rect 23212 22148 23268 23212
rect 23548 23044 23604 23326
rect 23772 23826 23828 23838
rect 23772 23774 23774 23826
rect 23826 23774 23828 23826
rect 23772 23380 23828 23774
rect 23772 23314 23828 23324
rect 23996 23154 24052 25228
rect 25228 24052 25284 25454
rect 25228 23986 25284 23996
rect 24220 23940 24276 23950
rect 24220 23846 24276 23884
rect 23996 23102 23998 23154
rect 24050 23102 24052 23154
rect 23996 23090 24052 23102
rect 24108 23714 24164 23726
rect 24108 23662 24110 23714
rect 24162 23662 24164 23714
rect 23548 22978 23604 22988
rect 23044 22092 23268 22148
rect 23884 22370 23940 22382
rect 23884 22318 23886 22370
rect 23938 22318 23940 22370
rect 23884 22260 23940 22318
rect 22988 21810 23044 22092
rect 23660 22036 23716 22046
rect 22988 21758 22990 21810
rect 23042 21758 23044 21810
rect 22988 21746 23044 21758
rect 23324 21924 23380 21934
rect 23324 21810 23380 21868
rect 23324 21758 23326 21810
rect 23378 21758 23380 21810
rect 23324 21746 23380 21758
rect 22876 20862 22878 20914
rect 22930 20862 22932 20914
rect 22876 20850 22932 20862
rect 23324 20804 23380 20814
rect 22764 20636 23044 20692
rect 22988 19124 23044 20636
rect 23212 20244 23268 20254
rect 23212 19234 23268 20188
rect 23324 20130 23380 20748
rect 23324 20078 23326 20130
rect 23378 20078 23380 20130
rect 23324 20066 23380 20078
rect 23212 19182 23214 19234
rect 23266 19182 23268 19234
rect 23212 19170 23268 19182
rect 23660 19234 23716 21980
rect 23884 21588 23940 22204
rect 24108 21924 24164 23662
rect 25452 23492 25508 26908
rect 25564 26898 25620 26908
rect 25676 26964 25732 26974
rect 25676 26962 25956 26964
rect 25676 26910 25678 26962
rect 25730 26910 25956 26962
rect 25676 26908 25956 26910
rect 25676 26898 25732 26908
rect 25900 25730 25956 26908
rect 26012 26402 26068 27244
rect 40012 27186 40068 27198
rect 40012 27134 40014 27186
rect 40066 27134 40068 27186
rect 26012 26350 26014 26402
rect 26066 26350 26068 26402
rect 26012 26338 26068 26350
rect 26124 27076 26180 27086
rect 25900 25678 25902 25730
rect 25954 25678 25956 25730
rect 25900 25666 25956 25678
rect 26124 25620 26180 27020
rect 37660 27074 37716 27086
rect 37660 27022 37662 27074
rect 37714 27022 37716 27074
rect 26012 25564 26180 25620
rect 28140 26180 28196 26190
rect 25788 25508 25844 25518
rect 25788 25414 25844 25452
rect 25900 25396 25956 25406
rect 25900 25302 25956 25340
rect 25900 25060 25956 25070
rect 26012 25060 26068 25564
rect 28140 25396 28196 26124
rect 28140 25330 28196 25340
rect 28588 26178 28644 26190
rect 28588 26126 28590 26178
rect 28642 26126 28644 26178
rect 25956 25004 26068 25060
rect 27468 25172 27524 25182
rect 25900 24722 25956 25004
rect 25900 24670 25902 24722
rect 25954 24670 25956 24722
rect 25900 24658 25956 24670
rect 26572 24612 26628 24622
rect 26124 24610 26628 24612
rect 26124 24558 26574 24610
rect 26626 24558 26628 24610
rect 26124 24556 26628 24558
rect 26124 24050 26180 24556
rect 26572 24546 26628 24556
rect 26124 23998 26126 24050
rect 26178 23998 26180 24050
rect 26124 23986 26180 23998
rect 26908 24052 26964 24062
rect 26684 23940 26740 23950
rect 26684 23846 26740 23884
rect 26908 23938 26964 23996
rect 26908 23886 26910 23938
rect 26962 23886 26964 23938
rect 26908 23874 26964 23886
rect 26236 23828 26292 23838
rect 26236 23734 26292 23772
rect 27244 23828 27300 23838
rect 27244 23734 27300 23772
rect 25452 23426 25508 23436
rect 26012 23714 26068 23726
rect 26012 23662 26014 23714
rect 26066 23662 26068 23714
rect 26012 23492 26068 23662
rect 26012 23426 26068 23436
rect 24444 23380 24500 23390
rect 24444 23286 24500 23324
rect 25564 23380 25620 23390
rect 24668 23156 24724 23166
rect 24668 23062 24724 23100
rect 24556 23042 24612 23054
rect 24556 22990 24558 23042
rect 24610 22990 24612 23042
rect 24108 21858 24164 21868
rect 24444 22146 24500 22158
rect 24444 22094 24446 22146
rect 24498 22094 24500 22146
rect 23884 21522 23940 21532
rect 24444 20580 24500 22094
rect 24556 21700 24612 22990
rect 25564 22596 25620 23324
rect 27468 23380 27524 25116
rect 28588 25172 28644 26126
rect 37660 26180 37716 27022
rect 40012 26292 40068 27134
rect 40012 26226 40068 26236
rect 37660 26114 37716 26124
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 40012 25618 40068 25630
rect 40012 25566 40014 25618
rect 40066 25566 40068 25618
rect 37660 25506 37716 25518
rect 37660 25454 37662 25506
rect 37714 25454 37716 25506
rect 28588 25106 28644 25116
rect 29148 25172 29204 25182
rect 29148 24946 29204 25116
rect 29148 24894 29150 24946
rect 29202 24894 29204 24946
rect 29148 24882 29204 24894
rect 27916 24612 27972 24622
rect 27692 23940 27748 23950
rect 27692 23846 27748 23884
rect 27916 23826 27972 24556
rect 28700 24612 28756 24622
rect 28700 24518 28756 24556
rect 37660 24612 37716 25454
rect 40012 24948 40068 25566
rect 40012 24882 40068 24892
rect 37660 24546 37716 24556
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 29260 23940 29316 23950
rect 27916 23774 27918 23826
rect 27970 23774 27972 23826
rect 27916 23762 27972 23774
rect 28028 23828 28084 23838
rect 28028 23734 28084 23772
rect 29260 23826 29316 23884
rect 30716 23940 30772 23950
rect 29260 23774 29262 23826
rect 29314 23774 29316 23826
rect 29260 23762 29316 23774
rect 29372 23828 29428 23838
rect 29428 23772 29540 23828
rect 29372 23734 29428 23772
rect 29036 23716 29092 23726
rect 28700 23714 29092 23716
rect 28700 23662 29038 23714
rect 29090 23662 29092 23714
rect 28700 23660 29092 23662
rect 27468 23378 27860 23380
rect 27468 23326 27470 23378
rect 27522 23326 27860 23378
rect 27468 23324 27860 23326
rect 27468 23314 27524 23324
rect 27804 23156 27860 23324
rect 27804 23154 27972 23156
rect 27804 23102 27806 23154
rect 27858 23102 27972 23154
rect 27804 23100 27972 23102
rect 27804 23090 27860 23100
rect 25004 22372 25060 22382
rect 25004 22278 25060 22316
rect 25564 22370 25620 22540
rect 26460 22596 26516 22606
rect 26460 22502 26516 22540
rect 25564 22318 25566 22370
rect 25618 22318 25620 22370
rect 25564 22306 25620 22318
rect 25900 22482 25956 22494
rect 25900 22430 25902 22482
rect 25954 22430 25956 22482
rect 25676 22260 25732 22270
rect 25676 22166 25732 22204
rect 24556 21634 24612 21644
rect 25228 21474 25284 21486
rect 25228 21422 25230 21474
rect 25282 21422 25284 21474
rect 24444 20514 24500 20524
rect 25116 20580 25172 20590
rect 23660 19182 23662 19234
rect 23714 19182 23716 19234
rect 23660 19170 23716 19182
rect 22988 19030 23044 19068
rect 22204 18622 22206 18674
rect 22258 18622 22260 18674
rect 22204 18610 22260 18622
rect 22316 19012 22372 19022
rect 21980 18510 21982 18562
rect 22034 18510 22036 18562
rect 21980 18498 22036 18510
rect 20748 18452 20804 18462
rect 20748 18358 20804 18396
rect 22092 18452 22148 18462
rect 22092 18358 22148 18396
rect 21420 18340 21476 18350
rect 21420 18246 21476 18284
rect 21644 18338 21700 18350
rect 21644 18286 21646 18338
rect 21698 18286 21700 18338
rect 20188 17390 20190 17442
rect 20242 17390 20244 17442
rect 20188 17378 20244 17390
rect 20300 17612 20468 17668
rect 21644 18004 21700 18286
rect 22316 18340 22372 18956
rect 23772 19012 23828 19022
rect 22652 18564 22708 18574
rect 22652 18470 22708 18508
rect 22764 18562 22820 18574
rect 23772 18564 23828 18956
rect 22764 18510 22766 18562
rect 22818 18510 22820 18562
rect 22764 18452 22820 18510
rect 22764 18386 22820 18396
rect 23436 18508 23828 18564
rect 23996 19010 24052 19022
rect 23996 18958 23998 19010
rect 24050 18958 24052 19010
rect 22316 18274 22372 18284
rect 21644 17666 21700 17948
rect 21644 17614 21646 17666
rect 21698 17614 21700 17666
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 16930 19684 16940
rect 20300 16996 20356 17612
rect 21644 17602 21700 17614
rect 22764 18226 22820 18238
rect 22764 18174 22766 18226
rect 22818 18174 22820 18226
rect 20300 16930 20356 16940
rect 20412 17442 20468 17454
rect 20412 17390 20414 17442
rect 20466 17390 20468 17442
rect 20412 16884 20468 17390
rect 21308 17444 21364 17454
rect 21308 17350 21364 17388
rect 21980 17444 22036 17454
rect 20412 16818 20468 16828
rect 20860 16996 20916 17006
rect 19516 16270 19518 16322
rect 19570 16270 19572 16322
rect 19516 16258 19572 16270
rect 19852 16098 19908 16110
rect 19852 16046 19854 16098
rect 19906 16046 19908 16098
rect 19628 15874 19684 15886
rect 19628 15822 19630 15874
rect 19682 15822 19684 15874
rect 19628 15540 19684 15822
rect 19852 15876 19908 16046
rect 19852 15820 20244 15876
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20076 15540 20132 15550
rect 20188 15540 20244 15820
rect 19628 15484 19908 15540
rect 19516 15428 19572 15438
rect 19572 15372 19684 15428
rect 19516 15362 19572 15372
rect 19068 15314 19460 15316
rect 19068 15262 19070 15314
rect 19122 15262 19294 15314
rect 19346 15262 19460 15314
rect 19068 15260 19460 15262
rect 19628 15314 19684 15372
rect 19628 15262 19630 15314
rect 19682 15262 19684 15314
rect 19068 15250 19124 15260
rect 19292 15250 19348 15260
rect 19628 15250 19684 15262
rect 19852 15314 19908 15484
rect 19852 15262 19854 15314
rect 19906 15262 19908 15314
rect 19852 15250 19908 15262
rect 20132 15484 20244 15540
rect 20412 15540 20468 15550
rect 20412 15538 20692 15540
rect 20412 15486 20414 15538
rect 20466 15486 20692 15538
rect 20412 15484 20692 15486
rect 20076 15314 20132 15484
rect 20412 15474 20468 15484
rect 20636 15426 20692 15484
rect 20860 15538 20916 16940
rect 21980 16770 22036 17388
rect 22764 17444 22820 18174
rect 22764 17378 22820 17388
rect 22204 17164 23156 17220
rect 22204 16994 22260 17164
rect 23100 17106 23156 17164
rect 23100 17054 23102 17106
rect 23154 17054 23156 17106
rect 23100 17042 23156 17054
rect 22204 16942 22206 16994
rect 22258 16942 22260 16994
rect 22204 16930 22260 16942
rect 22428 16994 22484 17006
rect 22428 16942 22430 16994
rect 22482 16942 22484 16994
rect 22428 16884 22484 16942
rect 23324 16994 23380 17006
rect 23324 16942 23326 16994
rect 23378 16942 23380 16994
rect 22428 16818 22484 16828
rect 22764 16884 22820 16894
rect 22764 16790 22820 16828
rect 21980 16718 21982 16770
rect 22034 16718 22036 16770
rect 21980 16706 22036 16718
rect 22988 16658 23044 16670
rect 22988 16606 22990 16658
rect 23042 16606 23044 16658
rect 20860 15486 20862 15538
rect 20914 15486 20916 15538
rect 20860 15474 20916 15486
rect 22092 15988 22148 15998
rect 20636 15374 20638 15426
rect 20690 15374 20692 15426
rect 20636 15362 20692 15374
rect 20076 15262 20078 15314
rect 20130 15262 20132 15314
rect 20076 15250 20132 15262
rect 20300 15314 20356 15326
rect 20300 15262 20302 15314
rect 20354 15262 20356 15314
rect 19180 14644 19236 14654
rect 18620 14642 19236 14644
rect 18620 14590 19182 14642
rect 19234 14590 19236 14642
rect 18620 14588 19236 14590
rect 15596 13022 15598 13074
rect 15650 13022 15652 13074
rect 15596 13010 15652 13022
rect 17612 13074 18004 13076
rect 17612 13022 17726 13074
rect 17778 13022 18004 13074
rect 17612 13020 18004 13022
rect 18284 14532 18340 14542
rect 18284 13074 18340 14476
rect 18956 13634 19012 13646
rect 18956 13582 18958 13634
rect 19010 13582 19012 13634
rect 18956 13524 19012 13582
rect 18956 13458 19012 13468
rect 18284 13022 18286 13074
rect 18338 13022 18340 13074
rect 14812 12964 14868 12974
rect 14700 12962 14868 12964
rect 14700 12910 14814 12962
rect 14866 12910 14868 12962
rect 14700 12908 14868 12910
rect 14812 12898 14868 12908
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 17500 3668 17556 3678
rect 17500 800 17556 3612
rect 17612 3554 17668 13020
rect 17724 13010 17780 13020
rect 18284 13010 18340 13022
rect 18396 4452 18452 4462
rect 17612 3502 17614 3554
rect 17666 3502 17668 3554
rect 17612 3490 17668 3502
rect 18172 4450 18452 4452
rect 18172 4398 18398 4450
rect 18450 4398 18452 4450
rect 18172 4396 18452 4398
rect 18172 800 18228 4396
rect 18396 4386 18452 4396
rect 19068 4338 19124 14588
rect 19180 14578 19236 14588
rect 19628 14532 19684 14542
rect 19628 14438 19684 14476
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20300 13524 20356 15262
rect 20972 15090 21028 15102
rect 20972 15038 20974 15090
rect 21026 15038 21028 15090
rect 20972 13860 21028 15038
rect 22092 14530 22148 15932
rect 22764 15426 22820 15438
rect 22764 15374 22766 15426
rect 22818 15374 22820 15426
rect 22764 14642 22820 15374
rect 22988 15314 23044 16606
rect 23324 16324 23380 16942
rect 23436 16994 23492 18508
rect 23996 18452 24052 18958
rect 23996 18386 24052 18396
rect 24220 18340 24276 18350
rect 23436 16942 23438 16994
rect 23490 16942 23492 16994
rect 23436 16930 23492 16942
rect 24108 18284 24220 18340
rect 24108 16994 24164 18284
rect 24220 18274 24276 18284
rect 25116 18340 25172 20524
rect 25228 20244 25284 21422
rect 25228 20178 25284 20188
rect 25564 18674 25620 18686
rect 25564 18622 25566 18674
rect 25618 18622 25620 18674
rect 25116 18274 25172 18284
rect 25228 18450 25284 18462
rect 25228 18398 25230 18450
rect 25282 18398 25284 18450
rect 25228 18228 25284 18398
rect 25452 18452 25508 18462
rect 25452 18358 25508 18396
rect 25228 18162 25284 18172
rect 25564 17780 25620 18622
rect 25900 18450 25956 22430
rect 26572 22484 26628 22494
rect 26572 22390 26628 22428
rect 27356 21700 27412 21710
rect 27356 21606 27412 21644
rect 27916 21588 27972 23100
rect 28028 23044 28084 23054
rect 28028 22260 28084 22988
rect 28588 23042 28644 23054
rect 28588 22990 28590 23042
rect 28642 22990 28644 23042
rect 28476 22596 28532 22606
rect 28588 22596 28644 22990
rect 28476 22594 28644 22596
rect 28476 22542 28478 22594
rect 28530 22542 28644 22594
rect 28476 22540 28644 22542
rect 28476 22530 28532 22540
rect 28588 22372 28644 22382
rect 28700 22372 28756 23660
rect 29036 23650 29092 23660
rect 28588 22370 28756 22372
rect 28588 22318 28590 22370
rect 28642 22318 28756 22370
rect 28588 22316 28756 22318
rect 28588 22306 28644 22316
rect 28476 22260 28532 22270
rect 28028 22258 28532 22260
rect 28028 22206 28030 22258
rect 28082 22206 28478 22258
rect 28530 22206 28532 22258
rect 28028 22204 28532 22206
rect 28028 22194 28084 22204
rect 28476 22194 28532 22204
rect 28028 21588 28084 21598
rect 27916 21532 28028 21588
rect 27916 20914 27972 21532
rect 28028 21494 28084 21532
rect 29372 21588 29428 21598
rect 29372 21494 29428 21532
rect 28924 21476 28980 21486
rect 28924 21474 29316 21476
rect 28924 21422 28926 21474
rect 28978 21422 29316 21474
rect 28924 21420 29316 21422
rect 28924 21410 28980 21420
rect 27916 20862 27918 20914
rect 27970 20862 27972 20914
rect 27580 20356 27636 20366
rect 27132 20132 27188 20142
rect 27132 20038 27188 20076
rect 26908 20018 26964 20030
rect 26908 19966 26910 20018
rect 26962 19966 26964 20018
rect 26908 19458 26964 19966
rect 27580 20018 27636 20300
rect 27916 20188 27972 20862
rect 28812 21362 28868 21374
rect 28812 21310 28814 21362
rect 28866 21310 28868 21362
rect 28812 20188 28868 21310
rect 29260 20914 29316 21420
rect 29260 20862 29262 20914
rect 29314 20862 29316 20914
rect 29260 20850 29316 20862
rect 29148 20802 29204 20814
rect 29148 20750 29150 20802
rect 29202 20750 29204 20802
rect 29148 20580 29204 20750
rect 29148 20514 29204 20524
rect 29372 20578 29428 20590
rect 29372 20526 29374 20578
rect 29426 20526 29428 20578
rect 27580 19966 27582 20018
rect 27634 19966 27636 20018
rect 27580 19954 27636 19966
rect 27804 20132 27972 20188
rect 28588 20132 28868 20188
rect 29372 20132 29428 20526
rect 29484 20580 29540 23772
rect 30716 23042 30772 23884
rect 37660 23940 37716 23950
rect 37660 23846 37716 23884
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 30716 22990 30718 23042
rect 30770 22990 30772 23042
rect 30716 22978 30772 22990
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 30716 21588 30772 21598
rect 29820 20804 29876 20814
rect 29820 20710 29876 20748
rect 30716 20804 30772 21532
rect 37660 21588 37716 21598
rect 37660 21494 37716 21532
rect 40012 21362 40068 21374
rect 40012 21310 40014 21362
rect 40066 21310 40068 21362
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 39788 20914 39844 20926
rect 39788 20862 39790 20914
rect 39842 20862 39844 20914
rect 30156 20690 30212 20702
rect 30156 20638 30158 20690
rect 30210 20638 30212 20690
rect 29596 20580 29652 20590
rect 30156 20580 30212 20638
rect 29484 20578 30212 20580
rect 29484 20526 29598 20578
rect 29650 20526 30212 20578
rect 29484 20524 30212 20526
rect 30268 20580 30324 20590
rect 29596 20514 29652 20524
rect 30268 20188 30324 20524
rect 30492 20578 30548 20590
rect 30492 20526 30494 20578
rect 30546 20526 30548 20578
rect 30492 20356 30548 20526
rect 30492 20290 30548 20300
rect 27804 20018 27860 20132
rect 28588 20130 28644 20132
rect 28588 20078 28590 20130
rect 28642 20078 28644 20130
rect 28588 20066 28644 20078
rect 29372 20066 29428 20076
rect 30156 20132 30324 20188
rect 27804 19966 27806 20018
rect 27858 19966 27860 20018
rect 26908 19406 26910 19458
rect 26962 19406 26964 19458
rect 26908 19394 26964 19406
rect 27020 19906 27076 19918
rect 27020 19854 27022 19906
rect 27074 19854 27076 19906
rect 26908 19010 26964 19022
rect 26908 18958 26910 19010
rect 26962 18958 26964 19010
rect 26908 18564 26964 18958
rect 26796 18508 26964 18564
rect 27020 18564 27076 19854
rect 25900 18398 25902 18450
rect 25954 18398 25956 18450
rect 25676 18340 25732 18350
rect 25732 18284 25844 18340
rect 25676 18246 25732 18284
rect 25676 17780 25732 17790
rect 25564 17778 25732 17780
rect 25564 17726 25678 17778
rect 25730 17726 25732 17778
rect 25564 17724 25732 17726
rect 25676 17714 25732 17724
rect 25004 17668 25060 17678
rect 25788 17668 25844 18284
rect 25004 17666 25172 17668
rect 25004 17614 25006 17666
rect 25058 17614 25172 17666
rect 25004 17612 25172 17614
rect 25004 17602 25060 17612
rect 24556 17444 24612 17454
rect 24444 17108 24500 17118
rect 24108 16942 24110 16994
rect 24162 16942 24164 16994
rect 24108 16930 24164 16942
rect 24220 17106 24500 17108
rect 24220 17054 24446 17106
rect 24498 17054 24500 17106
rect 24220 17052 24500 17054
rect 23324 16268 23940 16324
rect 23548 16100 23604 16110
rect 23436 16098 23604 16100
rect 23436 16046 23550 16098
rect 23602 16046 23604 16098
rect 23436 16044 23604 16046
rect 23436 15988 23492 16044
rect 23548 16034 23604 16044
rect 23436 15922 23492 15932
rect 23884 15538 23940 16268
rect 24220 16210 24276 17052
rect 24444 17042 24500 17052
rect 24444 16884 24500 16894
rect 24556 16884 24612 17388
rect 24444 16882 24612 16884
rect 24444 16830 24446 16882
rect 24498 16830 24612 16882
rect 24444 16828 24612 16830
rect 24780 16884 24836 16894
rect 24780 16882 25060 16884
rect 24780 16830 24782 16882
rect 24834 16830 25060 16882
rect 24780 16828 25060 16830
rect 24444 16818 24500 16828
rect 24780 16818 24836 16828
rect 24220 16158 24222 16210
rect 24274 16158 24276 16210
rect 24220 16146 24276 16158
rect 23884 15486 23886 15538
rect 23938 15486 23940 15538
rect 23884 15474 23940 15486
rect 25004 15540 25060 16828
rect 25116 15988 25172 17612
rect 25788 17602 25844 17612
rect 25452 17556 25508 17566
rect 25172 15932 25284 15988
rect 25116 15922 25172 15932
rect 25116 15540 25172 15550
rect 25004 15538 25172 15540
rect 25004 15486 25118 15538
rect 25170 15486 25172 15538
rect 25004 15484 25172 15486
rect 25116 15474 25172 15484
rect 22988 15262 22990 15314
rect 23042 15262 23044 15314
rect 22988 15250 23044 15262
rect 22764 14590 22766 14642
rect 22818 14590 22820 14642
rect 22764 14578 22820 14590
rect 23996 15202 24052 15214
rect 23996 15150 23998 15202
rect 24050 15150 24052 15202
rect 23996 14644 24052 15150
rect 24892 14644 24948 14654
rect 23996 14642 24948 14644
rect 23996 14590 24894 14642
rect 24946 14590 24948 14642
rect 23996 14588 24948 14590
rect 25228 14644 25284 15932
rect 25340 15428 25396 15438
rect 25340 15334 25396 15372
rect 25452 15426 25508 17500
rect 25900 17556 25956 18398
rect 26124 18450 26180 18462
rect 26124 18398 26126 18450
rect 26178 18398 26180 18450
rect 26124 18228 26180 18398
rect 26796 18452 26852 18508
rect 27020 18498 27076 18508
rect 27132 19458 27188 19470
rect 27132 19406 27134 19458
rect 27186 19406 27188 19458
rect 26796 18386 26852 18396
rect 26908 18338 26964 18350
rect 26908 18286 26910 18338
rect 26962 18286 26964 18338
rect 26796 18228 26852 18238
rect 26124 18226 26852 18228
rect 26124 18174 26798 18226
rect 26850 18174 26852 18226
rect 26124 18172 26852 18174
rect 26796 18162 26852 18172
rect 26908 17892 26964 18286
rect 26908 17826 26964 17836
rect 25900 17490 25956 17500
rect 26908 17668 26964 17678
rect 26684 16884 26740 16894
rect 26572 16828 26684 16884
rect 26348 16212 26404 16222
rect 25452 15374 25454 15426
rect 25506 15374 25508 15426
rect 25452 15362 25508 15374
rect 26236 16210 26404 16212
rect 26236 16158 26350 16210
rect 26402 16158 26404 16210
rect 26236 16156 26404 16158
rect 26236 15428 26292 16156
rect 26348 16146 26404 16156
rect 26348 15988 26404 15998
rect 26572 15988 26628 16828
rect 26684 16790 26740 16828
rect 26908 16098 26964 17612
rect 27132 16884 27188 19406
rect 27468 19012 27524 19022
rect 27804 19012 27860 19966
rect 27468 19010 27860 19012
rect 27468 18958 27470 19010
rect 27522 18958 27860 19010
rect 27468 18956 27860 18958
rect 27244 18452 27300 18462
rect 27468 18452 27524 18956
rect 28028 18564 28084 18574
rect 28028 18470 28084 18508
rect 27300 18396 27524 18452
rect 27244 16996 27300 18396
rect 30156 18338 30212 20132
rect 30716 19906 30772 20748
rect 37660 20804 37716 20814
rect 37660 20710 37716 20748
rect 39788 20244 39844 20862
rect 40012 20916 40068 21310
rect 40012 20850 40068 20860
rect 39788 20178 39844 20188
rect 40236 20242 40292 20254
rect 40236 20190 40238 20242
rect 40290 20190 40292 20242
rect 30716 19854 30718 19906
rect 30770 19854 30772 19906
rect 30716 19842 30772 19854
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 40236 19572 40292 20190
rect 40236 19506 40292 19516
rect 30156 18286 30158 18338
rect 30210 18286 30212 18338
rect 30156 18274 30212 18286
rect 37660 18450 37716 18462
rect 37660 18398 37662 18450
rect 37714 18398 37716 18450
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 27804 17892 27860 17902
rect 28252 17892 28308 17902
rect 27804 17778 27860 17836
rect 27804 17726 27806 17778
rect 27858 17726 27860 17778
rect 27804 17714 27860 17726
rect 27916 17890 28308 17892
rect 27916 17838 28254 17890
rect 28306 17838 28308 17890
rect 27916 17836 28308 17838
rect 27244 16930 27300 16940
rect 27132 16818 27188 16828
rect 27468 16770 27524 16782
rect 27468 16718 27470 16770
rect 27522 16718 27524 16770
rect 27356 16212 27412 16222
rect 27468 16212 27524 16718
rect 27916 16660 27972 17836
rect 28252 17826 28308 17836
rect 37660 17892 37716 18398
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 37660 17826 37716 17836
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 28252 17668 28308 17678
rect 28140 17556 28196 17566
rect 28140 17462 28196 17500
rect 28252 17554 28308 17612
rect 28252 17502 28254 17554
rect 28306 17502 28308 17554
rect 28252 17490 28308 17502
rect 29596 17668 29652 17678
rect 29260 17442 29316 17454
rect 29260 17390 29262 17442
rect 29314 17390 29316 17442
rect 29260 16996 29316 17390
rect 29260 16930 29316 16940
rect 29596 16772 29652 17612
rect 37660 17668 37716 17678
rect 37660 17574 37716 17612
rect 40012 17556 40068 17726
rect 40012 17490 40068 17500
rect 30044 16996 30100 17006
rect 30044 16902 30100 16940
rect 27356 16210 27524 16212
rect 27356 16158 27358 16210
rect 27410 16158 27524 16210
rect 27356 16156 27524 16158
rect 27580 16604 27972 16660
rect 29260 16770 29652 16772
rect 29260 16718 29598 16770
rect 29650 16718 29652 16770
rect 29260 16716 29652 16718
rect 27356 16146 27412 16156
rect 26908 16046 26910 16098
rect 26962 16046 26964 16098
rect 26908 16034 26964 16046
rect 27580 16098 27636 16604
rect 27580 16046 27582 16098
rect 27634 16046 27636 16098
rect 27580 16034 27636 16046
rect 29260 16098 29316 16716
rect 29596 16706 29652 16716
rect 37884 16882 37940 16894
rect 37884 16830 37886 16882
rect 37938 16830 37940 16882
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 29260 16046 29262 16098
rect 29314 16046 29316 16098
rect 29260 16034 29316 16046
rect 37660 16098 37716 16110
rect 37660 16046 37662 16098
rect 37714 16046 37716 16098
rect 26404 15932 26628 15988
rect 26348 15922 26404 15932
rect 26572 15538 26628 15932
rect 27132 15988 27188 15998
rect 27132 15894 27188 15932
rect 29484 15876 29540 15886
rect 29484 15782 29540 15820
rect 26572 15486 26574 15538
rect 26626 15486 26628 15538
rect 26572 15474 26628 15486
rect 26348 15428 26404 15438
rect 26236 15372 26348 15428
rect 26348 15362 26404 15372
rect 37660 15428 37716 16046
rect 37884 15876 37940 16830
rect 40012 16884 40068 16894
rect 40012 16770 40068 16828
rect 40012 16718 40014 16770
rect 40066 16718 40068 16770
rect 40012 16706 40068 16718
rect 40012 16212 40068 16222
rect 40012 16118 40068 16156
rect 37884 15810 37940 15820
rect 37660 15362 37716 15372
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 25340 14644 25396 14654
rect 25228 14642 25396 14644
rect 25228 14590 25342 14642
rect 25394 14590 25396 14642
rect 25228 14588 25396 14590
rect 22092 14478 22094 14530
rect 22146 14478 22148 14530
rect 21084 13860 21140 13870
rect 20972 13858 21140 13860
rect 20972 13806 21086 13858
rect 21138 13806 21140 13858
rect 20972 13804 21140 13806
rect 21084 13794 21140 13804
rect 21868 13748 21924 13758
rect 22092 13748 22148 14478
rect 22316 13748 22372 13758
rect 21868 13746 22372 13748
rect 21868 13694 21870 13746
rect 21922 13694 22318 13746
rect 22370 13694 22372 13746
rect 21868 13692 22372 13694
rect 21868 13682 21924 13692
rect 22316 13682 22372 13692
rect 20300 13458 20356 13468
rect 21084 13524 21140 13534
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19068 4286 19070 4338
rect 19122 4286 19124 4338
rect 19068 4274 19124 4286
rect 18844 4116 18900 4126
rect 18620 3668 18676 3678
rect 18620 3574 18676 3612
rect 18844 800 18900 4060
rect 20076 4116 20132 4126
rect 20076 4022 20132 4060
rect 20860 3668 20916 3678
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20860 800 20916 3612
rect 21084 3554 21140 13468
rect 24892 8428 24948 14588
rect 25340 14578 25396 14588
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 24556 8372 24948 8428
rect 22092 3668 22148 3678
rect 22092 3574 22148 3612
rect 24220 3668 24276 3678
rect 21084 3502 21086 3554
rect 21138 3502 21140 3554
rect 21084 3490 21140 3502
rect 24220 800 24276 3612
rect 24556 3554 24612 8372
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 20832 0 20944 800
rect 24192 0 24304 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 24892 38220 24948 38276
rect 20188 37436 20244 37492
rect 21420 37490 21476 37492
rect 21420 37438 21422 37490
rect 21422 37438 21474 37490
rect 21474 37438 21476 37490
rect 21420 37436 21476 37438
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 15708 27074 15764 27076
rect 15708 27022 15710 27074
rect 15710 27022 15762 27074
rect 15762 27022 15764 27074
rect 15708 27020 15764 27022
rect 16380 27020 16436 27076
rect 4172 26908 4228 26964
rect 1932 24892 1988 24948
rect 1932 24498 1988 24500
rect 1932 24446 1934 24498
rect 1934 24446 1986 24498
rect 1986 24446 1988 24498
rect 1932 24444 1988 24446
rect 1932 22930 1988 22932
rect 1932 22878 1934 22930
rect 1934 22878 1986 22930
rect 1986 22878 1988 22930
rect 1932 22876 1988 22878
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4284 25506 4340 25508
rect 4284 25454 4286 25506
rect 4286 25454 4338 25506
rect 4338 25454 4340 25506
rect 4284 25452 4340 25454
rect 13468 25452 13524 25508
rect 15260 25452 15316 25508
rect 17612 27020 17668 27076
rect 16492 26460 16548 26516
rect 17388 26514 17444 26516
rect 17388 26462 17390 26514
rect 17390 26462 17442 26514
rect 17442 26462 17444 26514
rect 17388 26460 17444 26462
rect 18732 27468 18788 27524
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19516 27468 19572 27524
rect 19628 27692 19684 27748
rect 18956 27020 19012 27076
rect 18508 26348 18564 26404
rect 16156 24946 16212 24948
rect 16156 24894 16158 24946
rect 16158 24894 16210 24946
rect 16210 24894 16212 24946
rect 16156 24892 16212 24894
rect 4284 24556 4340 24612
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 14700 24668 14756 24724
rect 14364 24610 14420 24612
rect 14364 24558 14366 24610
rect 14366 24558 14418 24610
rect 14418 24558 14420 24610
rect 14364 24556 14420 24558
rect 14028 23996 14084 24052
rect 14476 23996 14532 24052
rect 12908 23826 12964 23828
rect 12908 23774 12910 23826
rect 12910 23774 12962 23826
rect 12962 23774 12964 23826
rect 12908 23772 12964 23774
rect 14140 23826 14196 23828
rect 14140 23774 14142 23826
rect 14142 23774 14194 23826
rect 14194 23774 14196 23826
rect 14140 23772 14196 23774
rect 11564 23548 11620 23604
rect 4284 23154 4340 23156
rect 4284 23102 4286 23154
rect 4286 23102 4338 23154
rect 4338 23102 4340 23154
rect 4284 23100 4340 23102
rect 10892 23042 10948 23044
rect 10892 22990 10894 23042
rect 10894 22990 10946 23042
rect 10946 22990 10948 23042
rect 10892 22988 10948 22990
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 13804 23548 13860 23604
rect 14476 23154 14532 23156
rect 14476 23102 14478 23154
rect 14478 23102 14530 23154
rect 14530 23102 14532 23154
rect 14476 23100 14532 23102
rect 13020 23042 13076 23044
rect 13020 22990 13022 23042
rect 13022 22990 13074 23042
rect 13074 22990 13076 23042
rect 13020 22988 13076 22990
rect 14252 23042 14308 23044
rect 14252 22990 14254 23042
rect 14254 22990 14306 23042
rect 14306 22990 14308 23042
rect 14252 22988 14308 22990
rect 12684 22876 12740 22932
rect 13580 22876 13636 22932
rect 10892 22316 10948 22372
rect 13580 22428 13636 22484
rect 13804 22370 13860 22372
rect 13804 22318 13806 22370
rect 13806 22318 13858 22370
rect 13858 22318 13860 22370
rect 13804 22316 13860 22318
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4172 19852 4228 19908
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 11564 18396 11620 18452
rect 12796 18450 12852 18452
rect 12796 18398 12798 18450
rect 12798 18398 12850 18450
rect 12850 18398 12852 18450
rect 12796 18396 12852 18398
rect 15596 24722 15652 24724
rect 15596 24670 15598 24722
rect 15598 24670 15650 24722
rect 15650 24670 15652 24722
rect 15596 24668 15652 24670
rect 17052 24892 17108 24948
rect 15036 23996 15092 24052
rect 14700 22092 14756 22148
rect 14924 23548 14980 23604
rect 18060 24108 18116 24164
rect 16156 23548 16212 23604
rect 16940 23548 16996 23604
rect 17052 22876 17108 22932
rect 16828 22764 16884 22820
rect 16380 22316 16436 22372
rect 16044 22258 16100 22260
rect 16044 22206 16046 22258
rect 16046 22206 16098 22258
rect 16098 22206 16100 22258
rect 16044 22204 16100 22206
rect 16380 22146 16436 22148
rect 16380 22094 16382 22146
rect 16382 22094 16434 22146
rect 16434 22094 16436 22146
rect 16380 22092 16436 22094
rect 14924 21644 14980 21700
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4284 17666 4340 17668
rect 4284 17614 4286 17666
rect 4286 17614 4338 17666
rect 4338 17614 4340 17666
rect 4284 17612 4340 17614
rect 11228 17612 11284 17668
rect 1932 16828 1988 16884
rect 4284 16716 4340 16772
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 1932 16156 1988 16212
rect 13692 17500 13748 17556
rect 13468 16882 13524 16884
rect 13468 16830 13470 16882
rect 13470 16830 13522 16882
rect 13522 16830 13524 16882
rect 13468 16828 13524 16830
rect 11340 16770 11396 16772
rect 11340 16718 11342 16770
rect 11342 16718 11394 16770
rect 11394 16718 11396 16770
rect 11340 16716 11396 16718
rect 14364 19964 14420 20020
rect 16828 20748 16884 20804
rect 16828 20130 16884 20132
rect 16828 20078 16830 20130
rect 16830 20078 16882 20130
rect 16882 20078 16884 20130
rect 16828 20076 16884 20078
rect 16492 20018 16548 20020
rect 16492 19966 16494 20018
rect 16494 19966 16546 20018
rect 16546 19966 16548 20018
rect 16492 19964 16548 19966
rect 14364 19068 14420 19124
rect 14140 18956 14196 19012
rect 14028 18396 14084 18452
rect 16828 19292 16884 19348
rect 14812 18396 14868 18452
rect 14924 18508 14980 18564
rect 14140 17612 14196 17668
rect 15596 18396 15652 18452
rect 14700 17554 14756 17556
rect 14700 17502 14702 17554
rect 14702 17502 14754 17554
rect 14754 17502 14756 17554
rect 14700 17500 14756 17502
rect 14252 17388 14308 17444
rect 11340 15932 11396 15988
rect 14588 17388 14644 17444
rect 14364 16098 14420 16100
rect 14364 16046 14366 16098
rect 14366 16046 14418 16098
rect 14418 16046 14420 16098
rect 14364 16044 14420 16046
rect 16156 19010 16212 19012
rect 16156 18958 16158 19010
rect 16158 18958 16210 19010
rect 16210 18958 16212 19010
rect 16156 18956 16212 18958
rect 16156 18450 16212 18452
rect 16156 18398 16158 18450
rect 16158 18398 16210 18450
rect 16210 18398 16212 18450
rect 16156 18396 16212 18398
rect 14700 16882 14756 16884
rect 14700 16830 14702 16882
rect 14702 16830 14754 16882
rect 14754 16830 14756 16882
rect 14700 16828 14756 16830
rect 15148 16044 15204 16100
rect 14812 15986 14868 15988
rect 14812 15934 14814 15986
rect 14814 15934 14866 15986
rect 14866 15934 14868 15986
rect 14812 15932 14868 15934
rect 15148 15260 15204 15316
rect 14700 15036 14756 15092
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 16268 15314 16324 15316
rect 16268 15262 16270 15314
rect 16270 15262 16322 15314
rect 16322 15262 16324 15314
rect 16268 15260 16324 15262
rect 16604 15314 16660 15316
rect 16604 15262 16606 15314
rect 16606 15262 16658 15314
rect 16658 15262 16660 15314
rect 16604 15260 16660 15262
rect 17276 23938 17332 23940
rect 17276 23886 17278 23938
rect 17278 23886 17330 23938
rect 17330 23886 17332 23938
rect 17276 23884 17332 23886
rect 17724 23772 17780 23828
rect 18060 23548 18116 23604
rect 17500 23154 17556 23156
rect 17500 23102 17502 23154
rect 17502 23102 17554 23154
rect 17554 23102 17556 23154
rect 17500 23100 17556 23102
rect 17388 22204 17444 22260
rect 17276 21980 17332 22036
rect 17724 22482 17780 22484
rect 17724 22430 17726 22482
rect 17726 22430 17778 22482
rect 17778 22430 17780 22482
rect 17724 22428 17780 22430
rect 17612 22370 17668 22372
rect 17612 22318 17614 22370
rect 17614 22318 17666 22370
rect 17666 22318 17668 22370
rect 17612 22316 17668 22318
rect 17500 21756 17556 21812
rect 17612 21698 17668 21700
rect 17612 21646 17614 21698
rect 17614 21646 17666 21698
rect 17666 21646 17668 21698
rect 17612 21644 17668 21646
rect 17052 19516 17108 19572
rect 17388 19404 17444 19460
rect 18172 22930 18228 22932
rect 18172 22878 18174 22930
rect 18174 22878 18226 22930
rect 18226 22878 18228 22930
rect 18172 22876 18228 22878
rect 18620 23884 18676 23940
rect 19068 26348 19124 26404
rect 20972 27746 21028 27748
rect 20972 27694 20974 27746
rect 20974 27694 21026 27746
rect 21026 27694 21028 27746
rect 20972 27692 21028 27694
rect 20188 26796 20244 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19292 25340 19348 25396
rect 18620 23548 18676 23604
rect 18284 22764 18340 22820
rect 18508 22370 18564 22372
rect 18508 22318 18510 22370
rect 18510 22318 18562 22370
rect 18562 22318 18564 22370
rect 18508 22316 18564 22318
rect 17948 20860 18004 20916
rect 18284 20802 18340 20804
rect 18284 20750 18286 20802
rect 18286 20750 18338 20802
rect 18338 20750 18340 20802
rect 18284 20748 18340 20750
rect 18396 20018 18452 20020
rect 18396 19966 18398 20018
rect 18398 19966 18450 20018
rect 18450 19966 18452 20018
rect 18396 19964 18452 19966
rect 18284 19234 18340 19236
rect 18284 19182 18286 19234
rect 18286 19182 18338 19234
rect 18338 19182 18340 19234
rect 18284 19180 18340 19182
rect 18172 19122 18228 19124
rect 18172 19070 18174 19122
rect 18174 19070 18226 19122
rect 18226 19070 18228 19122
rect 18172 19068 18228 19070
rect 17500 19010 17556 19012
rect 17500 18958 17502 19010
rect 17502 18958 17554 19010
rect 17554 18958 17556 19010
rect 17500 18956 17556 18958
rect 17164 18396 17220 18452
rect 17948 18172 18004 18228
rect 17164 17500 17220 17556
rect 17500 15426 17556 15428
rect 17500 15374 17502 15426
rect 17502 15374 17554 15426
rect 17554 15374 17556 15426
rect 17500 15372 17556 15374
rect 17724 15820 17780 15876
rect 18732 23154 18788 23156
rect 18732 23102 18734 23154
rect 18734 23102 18786 23154
rect 18786 23102 18788 23154
rect 18732 23100 18788 23102
rect 18732 22428 18788 22484
rect 18732 22092 18788 22148
rect 18732 20130 18788 20132
rect 18732 20078 18734 20130
rect 18734 20078 18786 20130
rect 18786 20078 18788 20130
rect 18732 20076 18788 20078
rect 18620 19404 18676 19460
rect 18956 23714 19012 23716
rect 18956 23662 18958 23714
rect 18958 23662 19010 23714
rect 19010 23662 19012 23714
rect 18956 23660 19012 23662
rect 19068 22428 19124 22484
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 26124 38274 26180 38276
rect 26124 38222 26126 38274
rect 26126 38222 26178 38274
rect 26178 38222 26180 38274
rect 26124 38220 26180 38222
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 24108 27132 24164 27188
rect 22316 27074 22372 27076
rect 22316 27022 22318 27074
rect 22318 27022 22370 27074
rect 22370 27022 22372 27074
rect 22316 27020 22372 27022
rect 21532 26962 21588 26964
rect 21532 26910 21534 26962
rect 21534 26910 21586 26962
rect 21586 26910 21588 26962
rect 21532 26908 21588 26910
rect 21644 26796 21700 26852
rect 22428 26908 22484 26964
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 25116 27186 25172 27188
rect 25116 27134 25118 27186
rect 25118 27134 25170 27186
rect 25170 27134 25172 27186
rect 25116 27132 25172 27134
rect 25228 27020 25284 27076
rect 24220 26796 24276 26852
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20524 25394 20580 25396
rect 20524 25342 20526 25394
rect 20526 25342 20578 25394
rect 20578 25342 20580 25394
rect 20524 25340 20580 25342
rect 19404 23772 19460 23828
rect 19292 23154 19348 23156
rect 19292 23102 19294 23154
rect 19294 23102 19346 23154
rect 19346 23102 19348 23154
rect 19292 23100 19348 23102
rect 19292 22146 19348 22148
rect 19292 22094 19294 22146
rect 19294 22094 19346 22146
rect 19346 22094 19348 22146
rect 19292 22092 19348 22094
rect 19516 23548 19572 23604
rect 20860 25282 20916 25284
rect 20860 25230 20862 25282
rect 20862 25230 20914 25282
rect 20914 25230 20916 25282
rect 20860 25228 20916 25230
rect 20076 23660 20132 23716
rect 21196 24108 21252 24164
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19628 22594 19684 22596
rect 19628 22542 19630 22594
rect 19630 22542 19682 22594
rect 19682 22542 19684 22594
rect 19628 22540 19684 22542
rect 19852 23212 19908 23268
rect 19852 22482 19908 22484
rect 19852 22430 19854 22482
rect 19854 22430 19906 22482
rect 19906 22430 19908 22482
rect 19852 22428 19908 22430
rect 20636 23938 20692 23940
rect 20636 23886 20638 23938
rect 20638 23886 20690 23938
rect 20690 23886 20692 23938
rect 20636 23884 20692 23886
rect 19628 22092 19684 22148
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20076 21532 20132 21588
rect 19740 20860 19796 20916
rect 20076 20802 20132 20804
rect 20076 20750 20078 20802
rect 20078 20750 20130 20802
rect 20130 20750 20132 20802
rect 20076 20748 20132 20750
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 18956 19234 19012 19236
rect 18956 19182 18958 19234
rect 18958 19182 19010 19234
rect 19010 19182 19012 19234
rect 18956 19180 19012 19182
rect 18620 18620 18676 18676
rect 18844 18844 18900 18900
rect 18620 18450 18676 18452
rect 18620 18398 18622 18450
rect 18622 18398 18674 18450
rect 18674 18398 18676 18450
rect 18620 18396 18676 18398
rect 19180 18844 19236 18900
rect 19628 20076 19684 20132
rect 19404 20018 19460 20020
rect 19404 19966 19406 20018
rect 19406 19966 19458 20018
rect 19458 19966 19460 20018
rect 19404 19964 19460 19966
rect 20524 23436 20580 23492
rect 20412 22764 20468 22820
rect 20412 22594 20468 22596
rect 20412 22542 20414 22594
rect 20414 22542 20466 22594
rect 20466 22542 20468 22594
rect 20412 22540 20468 22542
rect 20300 22316 20356 22372
rect 21644 23996 21700 24052
rect 25004 26796 25060 26852
rect 25004 25452 25060 25508
rect 23436 25228 23492 25284
rect 22204 24108 22260 24164
rect 20972 23660 21028 23716
rect 20748 22482 20804 22484
rect 20748 22430 20750 22482
rect 20750 22430 20802 22482
rect 20802 22430 20804 22482
rect 20748 22428 20804 22430
rect 20188 20076 20244 20132
rect 20748 20076 20804 20132
rect 19628 19458 19684 19460
rect 19628 19406 19630 19458
rect 19630 19406 19682 19458
rect 19682 19406 19684 19458
rect 19628 19404 19684 19406
rect 20300 19292 20356 19348
rect 19404 19010 19460 19012
rect 19404 18958 19406 19010
rect 19406 18958 19458 19010
rect 19458 18958 19460 19010
rect 19404 18956 19460 18958
rect 18844 18562 18900 18564
rect 18844 18510 18846 18562
rect 18846 18510 18898 18562
rect 18898 18510 18900 18562
rect 18844 18508 18900 18510
rect 18508 17948 18564 18004
rect 18732 16940 18788 16996
rect 18284 15820 18340 15876
rect 18284 15484 18340 15540
rect 17612 15260 17668 15316
rect 16268 15036 16324 15092
rect 18508 15538 18564 15540
rect 18508 15486 18510 15538
rect 18510 15486 18562 15538
rect 18562 15486 18564 15538
rect 18508 15484 18564 15486
rect 18956 17276 19012 17332
rect 18396 15372 18452 15428
rect 19292 17948 19348 18004
rect 19068 16940 19124 16996
rect 19180 17164 19236 17220
rect 19180 16044 19236 16100
rect 19180 15874 19236 15876
rect 19180 15822 19182 15874
rect 19182 15822 19234 15874
rect 19234 15822 19236 15874
rect 19180 15820 19236 15822
rect 18956 15484 19012 15540
rect 18844 15372 18900 15428
rect 18172 15314 18228 15316
rect 18172 15262 18174 15314
rect 18174 15262 18226 15314
rect 18226 15262 18228 15314
rect 18172 15260 18228 15262
rect 16268 14530 16324 14532
rect 16268 14478 16270 14530
rect 16270 14478 16322 14530
rect 16322 14478 16324 14530
rect 16268 14476 16324 14478
rect 18732 15314 18788 15316
rect 18732 15262 18734 15314
rect 18734 15262 18786 15314
rect 18786 15262 18788 15314
rect 18732 15260 18788 15262
rect 19628 18844 19684 18900
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20188 18620 20244 18676
rect 21308 23266 21364 23268
rect 21308 23214 21310 23266
rect 21310 23214 21362 23266
rect 21362 23214 21364 23266
rect 21308 23212 21364 23214
rect 21084 22764 21140 22820
rect 21420 22540 21476 22596
rect 21868 23100 21924 23156
rect 21644 22204 21700 22260
rect 21756 22146 21812 22148
rect 21756 22094 21758 22146
rect 21758 22094 21810 22146
rect 21810 22094 21812 22146
rect 21756 22092 21812 22094
rect 23436 24108 23492 24164
rect 22876 23884 22932 23940
rect 22652 23154 22708 23156
rect 22652 23102 22654 23154
rect 22654 23102 22706 23154
rect 22706 23102 22708 23154
rect 22652 23100 22708 23102
rect 23660 24050 23716 24052
rect 23660 23998 23662 24050
rect 23662 23998 23714 24050
rect 23714 23998 23716 24050
rect 23660 23996 23716 23998
rect 22652 22258 22708 22260
rect 22652 22206 22654 22258
rect 22654 22206 22706 22258
rect 22706 22206 22708 22258
rect 22652 22204 22708 22206
rect 22316 21980 22372 22036
rect 22092 21756 22148 21812
rect 22540 21868 22596 21924
rect 21980 20188 22036 20244
rect 21644 19458 21700 19460
rect 21644 19406 21646 19458
rect 21646 19406 21698 19458
rect 21698 19406 21700 19458
rect 21644 19404 21700 19406
rect 21420 19346 21476 19348
rect 21420 19294 21422 19346
rect 21422 19294 21474 19346
rect 21474 19294 21476 19346
rect 21420 19292 21476 19294
rect 22092 19068 22148 19124
rect 19852 18508 19908 18564
rect 19516 18060 19572 18116
rect 22652 20748 22708 20804
rect 22988 22428 23044 22484
rect 22876 22316 22932 22372
rect 22876 21756 22932 21812
rect 23772 23324 23828 23380
rect 25228 23996 25284 24052
rect 24220 23938 24276 23940
rect 24220 23886 24222 23938
rect 24222 23886 24274 23938
rect 24274 23886 24276 23938
rect 24220 23884 24276 23886
rect 23548 22988 23604 23044
rect 22988 22092 23044 22148
rect 23884 22204 23940 22260
rect 23660 21980 23716 22036
rect 23324 21868 23380 21924
rect 23324 20802 23380 20804
rect 23324 20750 23326 20802
rect 23326 20750 23378 20802
rect 23378 20750 23380 20802
rect 23324 20748 23380 20750
rect 23212 20188 23268 20244
rect 26124 27074 26180 27076
rect 26124 27022 26126 27074
rect 26126 27022 26178 27074
rect 26178 27022 26180 27074
rect 26124 27020 26180 27022
rect 28140 26178 28196 26180
rect 28140 26126 28142 26178
rect 28142 26126 28194 26178
rect 28194 26126 28196 26178
rect 28140 26124 28196 26126
rect 25788 25506 25844 25508
rect 25788 25454 25790 25506
rect 25790 25454 25842 25506
rect 25842 25454 25844 25506
rect 25788 25452 25844 25454
rect 25900 25394 25956 25396
rect 25900 25342 25902 25394
rect 25902 25342 25954 25394
rect 25954 25342 25956 25394
rect 25900 25340 25956 25342
rect 28140 25340 28196 25396
rect 25900 25004 25956 25060
rect 27468 25116 27524 25172
rect 26908 23996 26964 24052
rect 26684 23938 26740 23940
rect 26684 23886 26686 23938
rect 26686 23886 26738 23938
rect 26738 23886 26740 23938
rect 26684 23884 26740 23886
rect 26236 23826 26292 23828
rect 26236 23774 26238 23826
rect 26238 23774 26290 23826
rect 26290 23774 26292 23826
rect 26236 23772 26292 23774
rect 27244 23826 27300 23828
rect 27244 23774 27246 23826
rect 27246 23774 27298 23826
rect 27298 23774 27300 23826
rect 27244 23772 27300 23774
rect 25452 23436 25508 23492
rect 26012 23436 26068 23492
rect 24444 23378 24500 23380
rect 24444 23326 24446 23378
rect 24446 23326 24498 23378
rect 24498 23326 24500 23378
rect 24444 23324 24500 23326
rect 25564 23324 25620 23380
rect 24668 23154 24724 23156
rect 24668 23102 24670 23154
rect 24670 23102 24722 23154
rect 24722 23102 24724 23154
rect 24668 23100 24724 23102
rect 24108 21868 24164 21924
rect 23884 21532 23940 21588
rect 40012 26236 40068 26292
rect 37660 26124 37716 26180
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 28588 25116 28644 25172
rect 29148 25116 29204 25172
rect 27916 24556 27972 24612
rect 27692 23938 27748 23940
rect 27692 23886 27694 23938
rect 27694 23886 27746 23938
rect 27746 23886 27748 23938
rect 27692 23884 27748 23886
rect 28700 24610 28756 24612
rect 28700 24558 28702 24610
rect 28702 24558 28754 24610
rect 28754 24558 28756 24610
rect 28700 24556 28756 24558
rect 40012 24892 40068 24948
rect 37660 24556 37716 24612
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 29260 23884 29316 23940
rect 28028 23826 28084 23828
rect 28028 23774 28030 23826
rect 28030 23774 28082 23826
rect 28082 23774 28084 23826
rect 28028 23772 28084 23774
rect 30716 23884 30772 23940
rect 29372 23826 29428 23828
rect 29372 23774 29374 23826
rect 29374 23774 29426 23826
rect 29426 23774 29428 23826
rect 29372 23772 29428 23774
rect 25564 22540 25620 22596
rect 25004 22370 25060 22372
rect 25004 22318 25006 22370
rect 25006 22318 25058 22370
rect 25058 22318 25060 22370
rect 25004 22316 25060 22318
rect 26460 22594 26516 22596
rect 26460 22542 26462 22594
rect 26462 22542 26514 22594
rect 26514 22542 26516 22594
rect 26460 22540 26516 22542
rect 25676 22258 25732 22260
rect 25676 22206 25678 22258
rect 25678 22206 25730 22258
rect 25730 22206 25732 22258
rect 25676 22204 25732 22206
rect 24556 21644 24612 21700
rect 24444 20524 24500 20580
rect 25116 20524 25172 20580
rect 22988 19122 23044 19124
rect 22988 19070 22990 19122
rect 22990 19070 23042 19122
rect 23042 19070 23044 19122
rect 22988 19068 23044 19070
rect 22316 19010 22372 19012
rect 22316 18958 22318 19010
rect 22318 18958 22370 19010
rect 22370 18958 22372 19010
rect 22316 18956 22372 18958
rect 20748 18450 20804 18452
rect 20748 18398 20750 18450
rect 20750 18398 20802 18450
rect 20802 18398 20804 18450
rect 20748 18396 20804 18398
rect 22092 18450 22148 18452
rect 22092 18398 22094 18450
rect 22094 18398 22146 18450
rect 22146 18398 22148 18450
rect 22092 18396 22148 18398
rect 21420 18338 21476 18340
rect 21420 18286 21422 18338
rect 21422 18286 21474 18338
rect 21474 18286 21476 18338
rect 21420 18284 21476 18286
rect 23772 19010 23828 19012
rect 23772 18958 23774 19010
rect 23774 18958 23826 19010
rect 23826 18958 23828 19010
rect 23772 18956 23828 18958
rect 22652 18562 22708 18564
rect 22652 18510 22654 18562
rect 22654 18510 22706 18562
rect 22706 18510 22708 18562
rect 22652 18508 22708 18510
rect 22764 18396 22820 18452
rect 22316 18284 22372 18340
rect 21644 17948 21700 18004
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19628 16940 19684 16996
rect 20300 16940 20356 16996
rect 21308 17442 21364 17444
rect 21308 17390 21310 17442
rect 21310 17390 21362 17442
rect 21362 17390 21364 17442
rect 21308 17388 21364 17390
rect 21980 17388 22036 17444
rect 20412 16828 20468 16884
rect 20860 16940 20916 16996
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19516 15372 19572 15428
rect 20076 15484 20132 15540
rect 22764 17388 22820 17444
rect 22428 16828 22484 16884
rect 22764 16882 22820 16884
rect 22764 16830 22766 16882
rect 22766 16830 22818 16882
rect 22818 16830 22820 16882
rect 22764 16828 22820 16830
rect 22092 15932 22148 15988
rect 18284 14476 18340 14532
rect 18956 13468 19012 13524
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 17500 3612 17556 3668
rect 19628 14530 19684 14532
rect 19628 14478 19630 14530
rect 19630 14478 19682 14530
rect 19682 14478 19684 14530
rect 19628 14476 19684 14478
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 23996 18396 24052 18452
rect 24220 18284 24276 18340
rect 25228 20188 25284 20244
rect 25116 18284 25172 18340
rect 25452 18450 25508 18452
rect 25452 18398 25454 18450
rect 25454 18398 25506 18450
rect 25506 18398 25508 18450
rect 25452 18396 25508 18398
rect 25228 18172 25284 18228
rect 26572 22482 26628 22484
rect 26572 22430 26574 22482
rect 26574 22430 26626 22482
rect 26626 22430 26628 22482
rect 26572 22428 26628 22430
rect 27356 21698 27412 21700
rect 27356 21646 27358 21698
rect 27358 21646 27410 21698
rect 27410 21646 27412 21698
rect 27356 21644 27412 21646
rect 28028 22988 28084 23044
rect 28028 21586 28084 21588
rect 28028 21534 28030 21586
rect 28030 21534 28082 21586
rect 28082 21534 28084 21586
rect 28028 21532 28084 21534
rect 29372 21586 29428 21588
rect 29372 21534 29374 21586
rect 29374 21534 29426 21586
rect 29426 21534 29428 21586
rect 29372 21532 29428 21534
rect 27580 20300 27636 20356
rect 27132 20130 27188 20132
rect 27132 20078 27134 20130
rect 27134 20078 27186 20130
rect 27186 20078 27188 20130
rect 27132 20076 27188 20078
rect 29148 20524 29204 20580
rect 37660 23938 37716 23940
rect 37660 23886 37662 23938
rect 37662 23886 37714 23938
rect 37714 23886 37716 23938
rect 37660 23884 37716 23886
rect 40012 23548 40068 23604
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 30716 21532 30772 21588
rect 29820 20802 29876 20804
rect 29820 20750 29822 20802
rect 29822 20750 29874 20802
rect 29874 20750 29876 20802
rect 29820 20748 29876 20750
rect 37660 21586 37716 21588
rect 37660 21534 37662 21586
rect 37662 21534 37714 21586
rect 37714 21534 37716 21586
rect 37660 21532 37716 21534
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 30716 20748 30772 20804
rect 30268 20578 30324 20580
rect 30268 20526 30270 20578
rect 30270 20526 30322 20578
rect 30322 20526 30324 20578
rect 30268 20524 30324 20526
rect 30492 20300 30548 20356
rect 29372 20076 29428 20132
rect 27020 18508 27076 18564
rect 25676 18338 25732 18340
rect 25676 18286 25678 18338
rect 25678 18286 25730 18338
rect 25730 18286 25732 18338
rect 25676 18284 25732 18286
rect 24556 17388 24612 17444
rect 23436 15932 23492 15988
rect 25788 17612 25844 17668
rect 25452 17500 25508 17556
rect 25116 15932 25172 15988
rect 25340 15426 25396 15428
rect 25340 15374 25342 15426
rect 25342 15374 25394 15426
rect 25394 15374 25396 15426
rect 25340 15372 25396 15374
rect 26796 18396 26852 18452
rect 26908 17836 26964 17892
rect 25900 17500 25956 17556
rect 26908 17612 26964 17668
rect 26684 16882 26740 16884
rect 26684 16830 26686 16882
rect 26686 16830 26738 16882
rect 26738 16830 26740 16882
rect 26684 16828 26740 16830
rect 28028 18562 28084 18564
rect 28028 18510 28030 18562
rect 28030 18510 28082 18562
rect 28082 18510 28084 18562
rect 28028 18508 28084 18510
rect 27244 18450 27300 18452
rect 27244 18398 27246 18450
rect 27246 18398 27298 18450
rect 27298 18398 27300 18450
rect 27244 18396 27300 18398
rect 37660 20802 37716 20804
rect 37660 20750 37662 20802
rect 37662 20750 37714 20802
rect 37714 20750 37716 20802
rect 37660 20748 37716 20750
rect 40012 20860 40068 20916
rect 39788 20188 39844 20244
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 40236 19516 40292 19572
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 27804 17836 27860 17892
rect 27244 16940 27300 16996
rect 27132 16828 27188 16884
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 37660 17836 37716 17892
rect 28252 17612 28308 17668
rect 28140 17554 28196 17556
rect 28140 17502 28142 17554
rect 28142 17502 28194 17554
rect 28194 17502 28196 17554
rect 28140 17500 28196 17502
rect 29596 17612 29652 17668
rect 29260 16940 29316 16996
rect 37660 17666 37716 17668
rect 37660 17614 37662 17666
rect 37662 17614 37714 17666
rect 37714 17614 37716 17666
rect 37660 17612 37716 17614
rect 40012 17500 40068 17556
rect 30044 16994 30100 16996
rect 30044 16942 30046 16994
rect 30046 16942 30098 16994
rect 30098 16942 30100 16994
rect 30044 16940 30100 16942
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 26348 15932 26404 15988
rect 27132 15986 27188 15988
rect 27132 15934 27134 15986
rect 27134 15934 27186 15986
rect 27186 15934 27188 15986
rect 27132 15932 27188 15934
rect 29484 15874 29540 15876
rect 29484 15822 29486 15874
rect 29486 15822 29538 15874
rect 29538 15822 29540 15874
rect 29484 15820 29540 15822
rect 26348 15372 26404 15428
rect 40012 16828 40068 16884
rect 40012 16210 40068 16212
rect 40012 16158 40014 16210
rect 40014 16158 40066 16210
rect 40066 16158 40068 16210
rect 40012 16156 40068 16158
rect 37884 15820 37940 15876
rect 37660 15372 37716 15428
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 20300 13468 20356 13524
rect 21084 13468 21140 13524
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 18844 4060 18900 4116
rect 18620 3666 18676 3668
rect 18620 3614 18622 3666
rect 18622 3614 18674 3666
rect 18674 3614 18676 3666
rect 18620 3612 18676 3614
rect 20076 4114 20132 4116
rect 20076 4062 20078 4114
rect 20078 4062 20130 4114
rect 20130 4062 20132 4114
rect 20076 4060 20132 4062
rect 20860 3612 20916 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 22092 3666 22148 3668
rect 22092 3614 22094 3666
rect 22094 3614 22146 3666
rect 22146 3614 22148 3666
rect 22092 3612 22148 3614
rect 24220 3612 24276 3668
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 24882 38220 24892 38276
rect 24948 38220 26124 38276
rect 26180 38220 26190 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 20178 37436 20188 37492
rect 20244 37436 21420 37492
rect 21476 37436 21486 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 19618 27692 19628 27748
rect 19684 27692 20972 27748
rect 21028 27692 21038 27748
rect 18722 27468 18732 27524
rect 18788 27468 19516 27524
rect 19572 27468 19582 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 24098 27132 24108 27188
rect 24164 27132 25116 27188
rect 25172 27132 25182 27188
rect 15698 27020 15708 27076
rect 15764 27020 16380 27076
rect 16436 27020 17612 27076
rect 17668 27020 18956 27076
rect 19012 27020 19022 27076
rect 22306 27020 22316 27076
rect 22372 27020 25228 27076
rect 25284 27020 26124 27076
rect 26180 27020 26190 27076
rect 0 26964 800 26992
rect 0 26908 4172 26964
rect 4228 26908 4238 26964
rect 21522 26908 21532 26964
rect 21588 26908 22428 26964
rect 22484 26908 22494 26964
rect 0 26880 800 26908
rect 20178 26796 20188 26852
rect 20244 26796 21644 26852
rect 21700 26796 24220 26852
rect 24276 26796 25004 26852
rect 25060 26796 25070 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 16482 26460 16492 26516
rect 16548 26460 17388 26516
rect 17444 26460 17454 26516
rect 18498 26348 18508 26404
rect 18564 26348 19068 26404
rect 19124 26348 19134 26404
rect 41200 26292 42000 26320
rect 40002 26236 40012 26292
rect 40068 26236 42000 26292
rect 41200 26208 42000 26236
rect 28130 26124 28140 26180
rect 28196 26124 37660 26180
rect 37716 26124 37726 26180
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 4274 25452 4284 25508
rect 4340 25452 13468 25508
rect 13524 25452 15260 25508
rect 15316 25452 15326 25508
rect 24994 25452 25004 25508
rect 25060 25452 25788 25508
rect 25844 25452 25854 25508
rect 19282 25340 19292 25396
rect 19348 25340 20524 25396
rect 20580 25340 20590 25396
rect 25890 25340 25900 25396
rect 25956 25340 28140 25396
rect 28196 25340 28206 25396
rect 20850 25228 20860 25284
rect 20916 25228 23436 25284
rect 23492 25228 23502 25284
rect 26852 25116 27468 25172
rect 27524 25116 28588 25172
rect 28644 25116 29148 25172
rect 29204 25116 29214 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 26852 25060 26908 25116
rect 25890 25004 25900 25060
rect 25956 25004 26908 25060
rect 0 24948 800 24976
rect 41200 24948 42000 24976
rect 0 24892 1932 24948
rect 1988 24892 1998 24948
rect 16146 24892 16156 24948
rect 16212 24892 17052 24948
rect 17108 24892 17118 24948
rect 40002 24892 40012 24948
rect 40068 24892 42000 24948
rect 0 24864 800 24892
rect 41200 24864 42000 24892
rect 14690 24668 14700 24724
rect 14756 24668 15596 24724
rect 15652 24668 15662 24724
rect 4274 24556 4284 24612
rect 4340 24556 14364 24612
rect 14420 24556 14430 24612
rect 27906 24556 27916 24612
rect 27972 24556 28700 24612
rect 28756 24556 37660 24612
rect 37716 24556 37726 24612
rect 1922 24444 1932 24500
rect 1988 24444 1998 24500
rect 0 24276 800 24304
rect 1932 24276 1988 24444
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 0 24220 1988 24276
rect 0 24192 800 24220
rect 18050 24108 18060 24164
rect 18116 24108 21196 24164
rect 21252 24108 22204 24164
rect 22260 24108 23436 24164
rect 23492 24108 23502 24164
rect 14018 23996 14028 24052
rect 14084 23996 14476 24052
rect 14532 23996 15036 24052
rect 15092 23996 21644 24052
rect 21700 23996 21710 24052
rect 23650 23996 23660 24052
rect 23716 23996 25228 24052
rect 25284 23996 26908 24052
rect 26964 23996 26974 24052
rect 17266 23884 17276 23940
rect 17332 23884 18620 23940
rect 18676 23884 18686 23940
rect 20626 23884 20636 23940
rect 20692 23884 22876 23940
rect 22932 23884 24220 23940
rect 24276 23884 24286 23940
rect 26674 23884 26684 23940
rect 26740 23884 27692 23940
rect 27748 23884 27758 23940
rect 29250 23884 29260 23940
rect 29316 23884 30716 23940
rect 30772 23884 37660 23940
rect 37716 23884 37726 23940
rect 12898 23772 12908 23828
rect 12964 23772 14140 23828
rect 14196 23772 14206 23828
rect 17714 23772 17724 23828
rect 17780 23772 19404 23828
rect 19460 23772 26236 23828
rect 26292 23772 26302 23828
rect 27234 23772 27244 23828
rect 27300 23772 28028 23828
rect 28084 23772 29372 23828
rect 29428 23772 29438 23828
rect 18946 23660 18956 23716
rect 19012 23660 20076 23716
rect 20132 23660 20972 23716
rect 21028 23660 21038 23716
rect 41200 23604 42000 23632
rect 11554 23548 11564 23604
rect 11620 23548 13804 23604
rect 13860 23548 14924 23604
rect 14980 23548 16156 23604
rect 16212 23548 16222 23604
rect 16930 23548 16940 23604
rect 16996 23548 18060 23604
rect 18116 23548 18126 23604
rect 18610 23548 18620 23604
rect 18676 23548 19516 23604
rect 19572 23548 19582 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 41200 23520 42000 23548
rect 20514 23436 20524 23492
rect 20580 23436 25452 23492
rect 25508 23436 26012 23492
rect 26068 23436 26078 23492
rect 23762 23324 23772 23380
rect 23828 23324 24444 23380
rect 24500 23324 25564 23380
rect 25620 23324 25630 23380
rect 19842 23212 19852 23268
rect 19908 23212 21308 23268
rect 21364 23212 21374 23268
rect 4274 23100 4284 23156
rect 4340 23100 8428 23156
rect 14466 23100 14476 23156
rect 14532 23100 17500 23156
rect 17556 23100 17566 23156
rect 18722 23100 18732 23156
rect 18788 23100 19292 23156
rect 19348 23100 19358 23156
rect 21858 23100 21868 23156
rect 21924 23100 22652 23156
rect 22708 23100 24668 23156
rect 24724 23100 24734 23156
rect 8372 23044 8428 23100
rect 8372 22988 10892 23044
rect 10948 22988 10958 23044
rect 13010 22988 13020 23044
rect 13076 22988 14252 23044
rect 14308 22988 14318 23044
rect 23538 22988 23548 23044
rect 23604 22988 28028 23044
rect 28084 22988 28094 23044
rect 0 22932 800 22960
rect 0 22876 1932 22932
rect 1988 22876 1998 22932
rect 12674 22876 12684 22932
rect 12740 22876 13580 22932
rect 13636 22876 13646 22932
rect 17042 22876 17052 22932
rect 17108 22876 18172 22932
rect 18228 22876 18238 22932
rect 0 22848 800 22876
rect 16818 22764 16828 22820
rect 16884 22764 18284 22820
rect 18340 22764 20412 22820
rect 20468 22764 21084 22820
rect 21140 22764 21150 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 19618 22540 19628 22596
rect 19684 22540 20412 22596
rect 20468 22540 21420 22596
rect 21476 22540 21486 22596
rect 25554 22540 25564 22596
rect 25620 22540 26460 22596
rect 26516 22540 26526 22596
rect 13570 22428 13580 22484
rect 13636 22428 17724 22484
rect 17780 22428 18732 22484
rect 18788 22428 18798 22484
rect 19058 22428 19068 22484
rect 19124 22428 19852 22484
rect 19908 22428 19918 22484
rect 20738 22428 20748 22484
rect 20804 22428 22988 22484
rect 23044 22428 26572 22484
rect 26628 22428 26638 22484
rect 10882 22316 10892 22372
rect 10948 22316 13804 22372
rect 13860 22316 13870 22372
rect 16370 22316 16380 22372
rect 16436 22316 17612 22372
rect 17668 22316 17678 22372
rect 18498 22316 18508 22372
rect 18564 22316 20300 22372
rect 20356 22316 20366 22372
rect 22866 22316 22876 22372
rect 22932 22316 25004 22372
rect 25060 22316 25070 22372
rect 15092 22204 16044 22260
rect 16100 22204 17388 22260
rect 17444 22204 17454 22260
rect 18732 22204 21644 22260
rect 21700 22204 22652 22260
rect 22708 22204 22718 22260
rect 23874 22204 23884 22260
rect 23940 22204 25676 22260
rect 25732 22204 25742 22260
rect 15092 22148 15148 22204
rect 18732 22148 18788 22204
rect 14690 22092 14700 22148
rect 14756 22092 15148 22148
rect 16370 22092 16380 22148
rect 16436 22092 18732 22148
rect 18788 22092 18798 22148
rect 19254 22092 19292 22148
rect 19348 22092 19358 22148
rect 19618 22092 19628 22148
rect 19684 22092 20244 22148
rect 21746 22092 21756 22148
rect 21812 22092 22988 22148
rect 23044 22092 23054 22148
rect 19628 22036 19684 22092
rect 17266 21980 17276 22036
rect 17332 21980 19684 22036
rect 20188 22036 20244 22092
rect 20188 21980 22316 22036
rect 22372 21980 23660 22036
rect 23716 21980 23726 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 22530 21868 22540 21924
rect 22596 21868 23324 21924
rect 23380 21868 24108 21924
rect 24164 21868 24174 21924
rect 17490 21756 17500 21812
rect 17556 21756 22092 21812
rect 22148 21756 22876 21812
rect 22932 21756 22942 21812
rect 14914 21644 14924 21700
rect 14980 21644 17612 21700
rect 17668 21644 17678 21700
rect 24546 21644 24556 21700
rect 24612 21644 27356 21700
rect 27412 21644 27422 21700
rect 20066 21532 20076 21588
rect 20132 21532 23884 21588
rect 23940 21532 23950 21588
rect 28018 21532 28028 21588
rect 28084 21532 29372 21588
rect 29428 21532 29438 21588
rect 30706 21532 30716 21588
rect 30772 21532 37660 21588
rect 37716 21532 37726 21588
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 41200 20916 42000 20944
rect 17938 20860 17948 20916
rect 18004 20860 19740 20916
rect 19796 20860 19806 20916
rect 40002 20860 40012 20916
rect 40068 20860 42000 20916
rect 41200 20832 42000 20860
rect 16818 20748 16828 20804
rect 16884 20748 18284 20804
rect 18340 20748 20076 20804
rect 20132 20748 20142 20804
rect 22642 20748 22652 20804
rect 22708 20748 23324 20804
rect 23380 20748 23390 20804
rect 29810 20748 29820 20804
rect 29876 20748 30716 20804
rect 30772 20748 30782 20804
rect 31892 20748 37660 20804
rect 37716 20748 37726 20804
rect 31892 20580 31948 20748
rect 24434 20524 24444 20580
rect 24500 20524 25116 20580
rect 25172 20524 29148 20580
rect 29204 20524 29214 20580
rect 30258 20524 30268 20580
rect 30324 20524 31948 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 27570 20300 27580 20356
rect 27636 20300 30492 20356
rect 30548 20300 30558 20356
rect 41200 20244 42000 20272
rect 21970 20188 21980 20244
rect 22036 20188 23212 20244
rect 23268 20188 25228 20244
rect 25284 20188 25294 20244
rect 39778 20188 39788 20244
rect 39844 20188 42000 20244
rect 41200 20160 42000 20188
rect 16818 20076 16828 20132
rect 16884 20076 18732 20132
rect 18788 20076 19628 20132
rect 19684 20076 19694 20132
rect 20178 20076 20188 20132
rect 20244 20076 20748 20132
rect 20804 20076 27132 20132
rect 27188 20076 29372 20132
rect 29428 20076 29438 20132
rect 14354 19964 14364 20020
rect 14420 19964 16492 20020
rect 16548 19964 16558 20020
rect 18386 19964 18396 20020
rect 18452 19964 19404 20020
rect 19460 19964 19470 20020
rect 18396 19908 18452 19964
rect 4162 19852 4172 19908
rect 4228 19852 18452 19908
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 15092 19516 17052 19572
rect 17108 19516 18676 19572
rect 40226 19516 40236 19572
rect 40292 19516 42000 19572
rect 15092 19124 15148 19516
rect 18620 19460 18676 19516
rect 41200 19488 42000 19516
rect 17378 19404 17388 19460
rect 17444 19404 17454 19460
rect 18610 19404 18620 19460
rect 18676 19404 18686 19460
rect 19618 19404 19628 19460
rect 19684 19404 21644 19460
rect 21700 19404 21710 19460
rect 17388 19348 17444 19404
rect 16818 19292 16828 19348
rect 16884 19292 20300 19348
rect 20356 19292 21420 19348
rect 21476 19292 21486 19348
rect 18274 19180 18284 19236
rect 18340 19180 18956 19236
rect 19012 19180 19022 19236
rect 14354 19068 14364 19124
rect 14420 19068 15148 19124
rect 15932 19068 18172 19124
rect 18228 19068 18238 19124
rect 22082 19068 22092 19124
rect 22148 19068 22988 19124
rect 23044 19068 23054 19124
rect 15932 19012 15988 19068
rect 14130 18956 14140 19012
rect 14196 18956 15988 19012
rect 16146 18956 16156 19012
rect 16212 18956 17500 19012
rect 17556 18956 19404 19012
rect 19460 18956 19470 19012
rect 22306 18956 22316 19012
rect 22372 18956 23772 19012
rect 23828 18956 23838 19012
rect 18834 18844 18844 18900
rect 18900 18844 19180 18900
rect 19236 18844 19628 18900
rect 19684 18844 19694 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 18610 18620 18620 18676
rect 18676 18620 20188 18676
rect 20244 18620 20254 18676
rect 14914 18508 14924 18564
rect 14980 18508 18844 18564
rect 18900 18508 19292 18564
rect 19348 18508 19358 18564
rect 19842 18508 19852 18564
rect 19908 18508 22652 18564
rect 22708 18508 22718 18564
rect 27010 18508 27020 18564
rect 27076 18508 28028 18564
rect 28084 18508 28094 18564
rect 11554 18396 11564 18452
rect 11620 18396 12796 18452
rect 12852 18396 14028 18452
rect 14084 18396 14812 18452
rect 14868 18396 15596 18452
rect 15652 18396 16156 18452
rect 16212 18396 16222 18452
rect 17154 18396 17164 18452
rect 17220 18396 18620 18452
rect 18676 18396 18686 18452
rect 20738 18396 20748 18452
rect 20804 18396 22092 18452
rect 22148 18396 22764 18452
rect 22820 18396 22830 18452
rect 23986 18396 23996 18452
rect 24052 18396 25452 18452
rect 25508 18396 25518 18452
rect 26786 18396 26796 18452
rect 26852 18396 27244 18452
rect 27300 18396 27310 18452
rect 21410 18284 21420 18340
rect 21476 18284 22316 18340
rect 22372 18284 22382 18340
rect 24210 18284 24220 18340
rect 24276 18284 25116 18340
rect 25172 18284 25676 18340
rect 25732 18284 25742 18340
rect 41200 18228 42000 18256
rect 17938 18172 17948 18228
rect 18004 18172 25228 18228
rect 25284 18172 25294 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 19516 18116 19572 18172
rect 41200 18144 42000 18172
rect 19506 18060 19516 18116
rect 19572 18060 19582 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 18498 17948 18508 18004
rect 18564 17948 19292 18004
rect 19348 17948 21644 18004
rect 21700 17948 21710 18004
rect 26898 17836 26908 17892
rect 26964 17836 27804 17892
rect 27860 17836 37660 17892
rect 37716 17836 37726 17892
rect 4274 17612 4284 17668
rect 4340 17612 11228 17668
rect 11284 17612 14140 17668
rect 14196 17612 14206 17668
rect 25778 17612 25788 17668
rect 25844 17612 26908 17668
rect 26964 17612 26974 17668
rect 28242 17612 28252 17668
rect 28308 17612 29596 17668
rect 29652 17612 37660 17668
rect 37716 17612 37726 17668
rect 41200 17556 42000 17584
rect 13682 17500 13692 17556
rect 13748 17500 14700 17556
rect 14756 17500 17164 17556
rect 17220 17500 17230 17556
rect 25442 17500 25452 17556
rect 25508 17500 25900 17556
rect 25956 17500 28140 17556
rect 28196 17500 28206 17556
rect 40002 17500 40012 17556
rect 40068 17500 42000 17556
rect 41200 17472 42000 17500
rect 14242 17388 14252 17444
rect 14308 17388 14588 17444
rect 14644 17388 21308 17444
rect 21364 17388 21980 17444
rect 22036 17388 22046 17444
rect 22754 17388 22764 17444
rect 22820 17388 24556 17444
rect 24612 17388 24622 17444
rect 18946 17276 18956 17332
rect 19012 17276 19236 17332
rect 19180 17220 19236 17276
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 19170 17164 19180 17220
rect 19236 17164 19246 17220
rect 22764 16996 22820 17388
rect 18722 16940 18732 16996
rect 18788 16940 19068 16996
rect 19124 16940 19628 16996
rect 19684 16940 20300 16996
rect 20356 16940 20860 16996
rect 20916 16940 20926 16996
rect 22428 16940 22820 16996
rect 26684 16940 27244 16996
rect 27300 16940 29260 16996
rect 29316 16940 30044 16996
rect 30100 16940 30110 16996
rect 0 16884 800 16912
rect 22428 16884 22484 16940
rect 26684 16884 26740 16940
rect 41200 16884 42000 16912
rect 0 16828 1932 16884
rect 1988 16828 1998 16884
rect 13458 16828 13468 16884
rect 13524 16828 14700 16884
rect 14756 16828 14766 16884
rect 20402 16828 20412 16884
rect 20468 16828 22260 16884
rect 22418 16828 22428 16884
rect 22484 16828 22494 16884
rect 22652 16828 22764 16884
rect 22820 16828 26516 16884
rect 26674 16828 26684 16884
rect 26740 16828 26750 16884
rect 26852 16828 27132 16884
rect 27188 16828 27198 16884
rect 40002 16828 40012 16884
rect 40068 16828 42000 16884
rect 0 16800 800 16828
rect 22204 16772 22260 16828
rect 22652 16772 22708 16828
rect 4274 16716 4284 16772
rect 4340 16716 11340 16772
rect 11396 16716 11406 16772
rect 22204 16716 22708 16772
rect 26460 16772 26516 16828
rect 26852 16772 26908 16828
rect 41200 16800 42000 16828
rect 26460 16716 26908 16772
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 0 16212 800 16240
rect 41200 16212 42000 16240
rect 0 16156 1932 16212
rect 1988 16156 1998 16212
rect 40002 16156 40012 16212
rect 40068 16156 42000 16212
rect 0 16128 800 16156
rect 41200 16128 42000 16156
rect 14354 16044 14364 16100
rect 14420 16044 15148 16100
rect 15204 16044 15214 16100
rect 19170 16044 19180 16100
rect 19236 16044 26908 16100
rect 11330 15932 11340 15988
rect 11396 15932 14812 15988
rect 14868 15932 14878 15988
rect 22082 15932 22092 15988
rect 22148 15932 23436 15988
rect 23492 15932 25116 15988
rect 25172 15932 26348 15988
rect 26404 15932 26414 15988
rect 26852 15876 26908 16044
rect 27122 15932 27132 15988
rect 27188 15932 27198 15988
rect 27132 15876 27188 15932
rect 17714 15820 17724 15876
rect 17780 15820 18284 15876
rect 18340 15820 19180 15876
rect 19236 15820 19246 15876
rect 26852 15820 27188 15876
rect 29474 15820 29484 15876
rect 29540 15820 37884 15876
rect 37940 15820 37950 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 18274 15484 18284 15540
rect 18340 15484 18508 15540
rect 18564 15484 18956 15540
rect 19012 15484 20076 15540
rect 20132 15484 20142 15540
rect 16268 15372 17500 15428
rect 17556 15372 18396 15428
rect 18452 15372 18462 15428
rect 18834 15372 18844 15428
rect 18900 15372 19516 15428
rect 19572 15372 19582 15428
rect 25330 15372 25340 15428
rect 25396 15372 26348 15428
rect 26404 15372 37660 15428
rect 37716 15372 37726 15428
rect 16268 15316 16324 15372
rect 15138 15260 15148 15316
rect 15204 15260 16268 15316
rect 16324 15260 16334 15316
rect 16594 15260 16604 15316
rect 16660 15260 17612 15316
rect 17668 15260 17678 15316
rect 18162 15260 18172 15316
rect 18228 15260 18732 15316
rect 18788 15260 18798 15316
rect 14690 15036 14700 15092
rect 14756 15036 16268 15092
rect 16324 15036 16334 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 16258 14476 16268 14532
rect 16324 14476 18284 14532
rect 18340 14476 19628 14532
rect 19684 14476 19694 14532
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 18946 13468 18956 13524
rect 19012 13468 20300 13524
rect 20356 13468 21084 13524
rect 21140 13468 21150 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 18834 4060 18844 4116
rect 18900 4060 20076 4116
rect 20132 4060 20142 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 17490 3612 17500 3668
rect 17556 3612 18620 3668
rect 18676 3612 18686 3668
rect 20850 3612 20860 3668
rect 20916 3612 22092 3668
rect 22148 3612 22158 3668
rect 24210 3612 24220 3668
rect 24276 3612 25564 3668
rect 25620 3612 25630 3668
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19292 22092 19348 22148
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 19292 18508 19348 18564
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 19292 22148 19348 22158
rect 19292 18564 19348 22092
rect 19292 18498 19348 18508
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_
timestamp 1698175906
transform -1 0 21840 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24192 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16352 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _109_
timestamp 1698175906
transform 1 0 16352 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21280 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23632 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _112_
timestamp 1698175906
transform -1 0 24416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_
timestamp 1698175906
transform -1 0 23520 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21840 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _115_
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _116_
timestamp 1698175906
transform -1 0 19824 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _117_
timestamp 1698175906
transform 1 0 22512 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _118_
timestamp 1698175906
transform 1 0 18592 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform -1 0 19152 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698175906
transform -1 0 20944 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _121_
timestamp 1698175906
transform 1 0 19936 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21840 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _123_
timestamp 1698175906
transform -1 0 23296 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _124_
timestamp 1698175906
transform -1 0 14448 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform -1 0 17696 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform -1 0 23520 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _127_
timestamp 1698175906
transform -1 0 21952 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _128_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_
timestamp 1698175906
transform -1 0 16576 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14896 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _131_
timestamp 1698175906
transform -1 0 18928 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _132_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13664 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _134_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14672 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _135_
timestamp 1698175906
transform -1 0 13104 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _136_
timestamp 1698175906
transform -1 0 26768 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _138_
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _139_
timestamp 1698175906
transform -1 0 20944 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _140_
timestamp 1698175906
transform -1 0 20048 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _141_
timestamp 1698175906
transform 1 0 20384 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _142_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24864 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _143_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23968 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _144_
timestamp 1698175906
transform -1 0 22064 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _145_
timestamp 1698175906
transform -1 0 16688 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _146_
timestamp 1698175906
transform 1 0 16128 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _147_
timestamp 1698175906
transform 1 0 22288 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _148_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17360 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _149_
timestamp 1698175906
transform -1 0 23968 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _150_
timestamp 1698175906
transform -1 0 25536 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _151_
timestamp 1698175906
transform -1 0 20384 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _152_
timestamp 1698175906
transform -1 0 19376 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _153_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24864 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _154_
timestamp 1698175906
transform -1 0 25648 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _155_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21952 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _156_
timestamp 1698175906
transform -1 0 24864 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _157_
timestamp 1698175906
transform -1 0 24416 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698175906
transform -1 0 23744 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _159_
timestamp 1698175906
transform 1 0 14560 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform -1 0 15008 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _161_
timestamp 1698175906
transform 1 0 14448 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _162_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23184 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _163_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19152 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _164_
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _165_
timestamp 1698175906
transform -1 0 20160 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _166_
timestamp 1698175906
transform -1 0 20048 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _167_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21840 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _168_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19376 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _169_
timestamp 1698175906
transform -1 0 21616 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _170_
timestamp 1698175906
transform -1 0 17472 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _171_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16912 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _172_
timestamp 1698175906
transform -1 0 17920 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _173_
timestamp 1698175906
transform -1 0 21840 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _174_
timestamp 1698175906
transform -1 0 20944 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _175_
timestamp 1698175906
transform -1 0 19488 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _176_
timestamp 1698175906
transform -1 0 19264 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _177_
timestamp 1698175906
transform -1 0 18256 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _178_
timestamp 1698175906
transform -1 0 18480 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _179_
timestamp 1698175906
transform 1 0 19376 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _180_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 -1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _181_
timestamp 1698175906
transform 1 0 20496 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _182_
timestamp 1698175906
transform -1 0 18928 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _183_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18928 0 -1 23520
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _184_
timestamp 1698175906
transform 1 0 26768 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _185_
timestamp 1698175906
transform -1 0 28224 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _186_
timestamp 1698175906
transform 1 0 25872 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _187_
timestamp 1698175906
transform 1 0 25648 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _188_
timestamp 1698175906
transform -1 0 25872 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _189_
timestamp 1698175906
transform -1 0 18144 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _190_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18928 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _191_
timestamp 1698175906
transform -1 0 17024 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _192_
timestamp 1698175906
transform -1 0 15792 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _193_
timestamp 1698175906
transform 1 0 15792 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _194_
timestamp 1698175906
transform -1 0 14336 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _195_
timestamp 1698175906
transform 1 0 14000 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _196_
timestamp 1698175906
transform 1 0 13888 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _197_
timestamp 1698175906
transform -1 0 13104 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _198_
timestamp 1698175906
transform 1 0 30016 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _199_
timestamp 1698175906
transform 1 0 26768 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _200_
timestamp 1698175906
transform -1 0 30016 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _201_
timestamp 1698175906
transform -1 0 29120 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _202_
timestamp 1698175906
transform 1 0 18480 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _203_
timestamp 1698175906
transform 1 0 28000 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _204_
timestamp 1698175906
transform -1 0 27664 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _205_
timestamp 1698175906
transform -1 0 27104 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _206_
timestamp 1698175906
transform 1 0 23520 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _207_
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _208_
timestamp 1698175906
transform -1 0 29568 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _209_
timestamp 1698175906
transform -1 0 28784 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21840 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform -1 0 14448 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 12656 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 11312 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform -1 0 28336 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 19824 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 17472 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 23296 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 22064 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform -1 0 14448 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 15568 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 19376 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 16128 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform -1 0 22064 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 25648 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 14672 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform -1 0 16576 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform -1 0 14000 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 11312 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 27104 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 27664 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 26544 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform 1 0 24752 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 27664 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _238_
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _239_
timestamp 1698175906
transform -1 0 18928 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__144__B dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__164__B
timestamp 1698175906
transform -1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__A1
timestamp 1698175906
transform 1 0 19152 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__A1
timestamp 1698175906
transform 1 0 28000 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 25312 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 14672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 16128 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 14784 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 29344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 19600 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 20944 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 26544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 26096 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 15568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 19600 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 19152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 19600 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 22288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 29120 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 28560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform -1 0 18368 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 16800 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 14896 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 15008 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 26880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 27440 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 30016 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 29232 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 27440 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 18368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 22848 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 23184 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698175906
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698175906
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_150
timestamp 1698175906
transform 1 0 18144 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_155
timestamp 1698175906
transform 1 0 18704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_183 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21840 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_199
timestamp 1698175906
transform 1 0 23632 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_115
timestamp 1698175906
transform 1 0 14224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_148
timestamp 1698175906
transform 1 0 17920 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_152
timestamp 1698175906
transform 1 0 18368 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_168
timestamp 1698175906
transform 1 0 20160 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_172
timestamp 1698175906
transform 1 0 20608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_150
timestamp 1698175906
transform 1 0 18144 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_154
timestamp 1698175906
transform 1 0 18592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_185
timestamp 1698175906
transform 1 0 22064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_189
timestamp 1698175906
transform 1 0 22512 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_205
timestamp 1698175906
transform 1 0 24304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_131
timestamp 1698175906
transform 1 0 16016 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_161
timestamp 1698175906
transform 1 0 19376 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_165
timestamp 1698175906
transform 1 0 19824 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698175906
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_181
timestamp 1698175906
transform 1 0 21616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_212
timestamp 1698175906
transform 1 0 25088 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_216
timestamp 1698175906
transform 1 0 25536 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_232
timestamp 1698175906
transform 1 0 27328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_240
timestamp 1698175906
transform 1 0 28224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_117
timestamp 1698175906
transform 1 0 14448 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_121
timestamp 1698175906
transform 1 0 14896 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_129
timestamp 1698175906
transform 1 0 15792 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_131
timestamp 1698175906
transform 1 0 16016 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_177
timestamp 1698175906
transform 1 0 21168 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_185
timestamp 1698175906
transform 1 0 22064 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_189
timestamp 1698175906
transform 1 0 22512 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_196
timestamp 1698175906
transform 1 0 23296 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_204
timestamp 1698175906
transform 1 0 24192 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698175906
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_217
timestamp 1698175906
transform 1 0 25648 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_227
timestamp 1698175906
transform 1 0 26768 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_259
timestamp 1698175906
transform 1 0 30352 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_275
timestamp 1698175906
transform 1 0 32144 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_109
timestamp 1698175906
transform 1 0 13552 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_123
timestamp 1698175906
transform 1 0 15120 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_139
timestamp 1698175906
transform 1 0 16912 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_143
timestamp 1698175906
transform 1 0 17360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_150
timestamp 1698175906
transform 1 0 18144 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_157
timestamp 1698175906
transform 1 0 18928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_167
timestamp 1698175906
transform 1 0 20048 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_193
timestamp 1698175906
transform 1 0 22960 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_195
timestamp 1698175906
transform 1 0 23184 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_225
timestamp 1698175906
transform 1 0 26544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_235
timestamp 1698175906
transform 1 0 27664 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_253
timestamp 1698175906
transform 1 0 29680 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_285
timestamp 1698175906
transform 1 0 33264 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_301
timestamp 1698175906
transform 1 0 35056 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_309
timestamp 1698175906
transform 1 0 35952 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_313
timestamp 1698175906
transform 1 0 36400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 37296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 4480 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_125
timestamp 1698175906
transform 1 0 15344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_129
timestamp 1698175906
transform 1 0 15792 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698175906
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_150
timestamp 1698175906
transform 1 0 18144 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_154
timestamp 1698175906
transform 1 0 18592 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_162
timestamp 1698175906
transform 1 0 19488 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_178
timestamp 1698175906
transform 1 0 21280 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_182
timestamp 1698175906
transform 1 0 21728 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_199
timestamp 1698175906
transform 1 0 23632 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_201
timestamp 1698175906
transform 1 0 23856 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_220
timestamp 1698175906
transform 1 0 25984 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_224
timestamp 1698175906
transform 1 0 26432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_254
timestamp 1698175906
transform 1 0 29792 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_258
timestamp 1698175906
transform 1 0 30240 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_274
timestamp 1698175906
transform 1 0 32032 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698175906
transform 1 0 32480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 36512 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 37408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_111
timestamp 1698175906
transform 1 0 13776 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_122
timestamp 1698175906
transform 1 0 15008 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_154
timestamp 1698175906
transform 1 0 18592 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_162
timestamp 1698175906
transform 1 0 19488 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698175906
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_183
timestamp 1698175906
transform 1 0 21840 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_199
timestamp 1698175906
transform 1 0 23632 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_207
timestamp 1698175906
transform 1 0 24528 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698175906
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_251
timestamp 1698175906
transform 1 0 29456 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_88
timestamp 1698175906
transform 1 0 11200 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_96
timestamp 1698175906
transform 1 0 12096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_100
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_130
timestamp 1698175906
transform 1 0 15904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_134
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698175906
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_150
timestamp 1698175906
transform 1 0 18144 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_152
timestamp 1698175906
transform 1 0 18368 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_168
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_194
timestamp 1698175906
transform 1 0 23072 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_223
timestamp 1698175906
transform 1 0 26320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_225
timestamp 1698175906
transform 1 0 26544 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_259
timestamp 1698175906
transform 1 0 30352 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_275
timestamp 1698175906
transform 1 0 32144 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_69
timestamp 1698175906
transform 1 0 9072 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_85
timestamp 1698175906
transform 1 0 10864 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_93
timestamp 1698175906
transform 1 0 11760 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_97
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_119
timestamp 1698175906
transform 1 0 14672 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_127
timestamp 1698175906
transform 1 0 15568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_129
timestamp 1698175906
transform 1 0 15792 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_146
timestamp 1698175906
transform 1 0 17696 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_165
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_188
timestamp 1698175906
transform 1 0 22400 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_203
timestamp 1698175906
transform 1 0 24080 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_219
timestamp 1698175906
transform 1 0 25872 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_227
timestamp 1698175906
transform 1 0 26768 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_230
timestamp 1698175906
transform 1 0 27104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_232
timestamp 1698175906
transform 1 0 27328 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_235
timestamp 1698175906
transform 1 0 27664 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698175906
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_88
timestamp 1698175906
transform 1 0 11200 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_118
timestamp 1698175906
transform 1 0 14560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_122
timestamp 1698175906
transform 1 0 15008 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_130
timestamp 1698175906
transform 1 0 15904 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_150
timestamp 1698175906
transform 1 0 18144 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_220
timestamp 1698175906
transform 1 0 25984 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_224
timestamp 1698175906
transform 1 0 26432 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_226
timestamp 1698175906
transform 1 0 26656 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_264
timestamp 1698175906
transform 1 0 30912 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_330
timestamp 1698175906
transform 1 0 38304 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_338
timestamp 1698175906
transform 1 0 39200 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_342
timestamp 1698175906
transform 1 0 39648 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_344
timestamp 1698175906
transform 1 0 39872 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_111
timestamp 1698175906
transform 1 0 13776 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_121
timestamp 1698175906
transform 1 0 14896 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_129
timestamp 1698175906
transform 1 0 15792 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_137
timestamp 1698175906
transform 1 0 16688 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_141
timestamp 1698175906
transform 1 0 17136 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698175906
transform 1 0 20720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_185
timestamp 1698175906
transform 1 0 22064 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_261
timestamp 1698175906
transform 1 0 30576 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_293
timestamp 1698175906
transform 1 0 34160 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_309
timestamp 1698175906
transform 1 0 35952 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_313
timestamp 1698175906
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_104
timestamp 1698175906
transform 1 0 12992 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_120
timestamp 1698175906
transform 1 0 14784 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_128
timestamp 1698175906
transform 1 0 15680 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_198
timestamp 1698175906
transform 1 0 23520 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698175906
transform 1 0 24416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_241
timestamp 1698175906
transform 1 0 28336 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_243
timestamp 1698175906
transform 1 0 28560 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_248
timestamp 1698175906
transform 1 0 29120 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_252
timestamp 1698175906
transform 1 0 29568 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_268
timestamp 1698175906
transform 1 0 31360 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698175906
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_116
timestamp 1698175906
transform 1 0 14336 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_124
timestamp 1698175906
transform 1 0 15232 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_128
timestamp 1698175906
transform 1 0 15680 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_157
timestamp 1698175906
transform 1 0 18928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_167
timestamp 1698175906
transform 1 0 20048 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_177
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_227
timestamp 1698175906
transform 1 0 26768 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_235
timestamp 1698175906
transform 1 0 27664 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_237
timestamp 1698175906
transform 1 0 27888 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 4480 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_80
timestamp 1698175906
transform 1 0 10304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_119
timestamp 1698175906
transform 1 0 14672 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_123
timestamp 1698175906
transform 1 0 15120 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_131
timestamp 1698175906
transform 1 0 16016 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_135
timestamp 1698175906
transform 1 0 16464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_137
timestamp 1698175906
transform 1 0 16688 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_228
timestamp 1698175906
transform 1 0 26880 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_232
timestamp 1698175906
transform 1 0 27328 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_264
timestamp 1698175906
transform 1 0 30912 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 40320 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_69
timestamp 1698175906
transform 1 0 9072 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_85
timestamp 1698175906
transform 1 0 10864 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_93
timestamp 1698175906
transform 1 0 11760 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_97
timestamp 1698175906
transform 1 0 12208 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_111
timestamp 1698175906
transform 1 0 13776 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_120
timestamp 1698175906
transform 1 0 14784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_124
timestamp 1698175906
transform 1 0 15232 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_132
timestamp 1698175906
transform 1 0 16128 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_136
timestamp 1698175906
transform 1 0 16576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_138
timestamp 1698175906
transform 1 0 16800 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_149
timestamp 1698175906
transform 1 0 18032 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_151
timestamp 1698175906
transform 1 0 18256 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_167
timestamp 1698175906
transform 1 0 20048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_185
timestamp 1698175906
transform 1 0 22064 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_195
timestamp 1698175906
transform 1 0 23184 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_206
timestamp 1698175906
transform 1 0 24416 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_214
timestamp 1698175906
transform 1 0 25312 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_218
timestamp 1698175906
transform 1 0 25760 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_233
timestamp 1698175906
transform 1 0 27440 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_240
timestamp 1698175906
transform 1 0 28224 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_252
timestamp 1698175906
transform 1 0 29568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_284
timestamp 1698175906
transform 1 0 33152 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_300
timestamp 1698175906
transform 1 0 34944 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_308
timestamp 1698175906
transform 1 0 35840 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_312
timestamp 1698175906
transform 1 0 36288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698175906
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 4480 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 8064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_88
timestamp 1698175906
transform 1 0 11200 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_118
timestamp 1698175906
transform 1 0 14560 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_120
timestamp 1698175906
transform 1 0 14784 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_135
timestamp 1698175906
transform 1 0 16464 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_158
timestamp 1698175906
transform 1 0 19040 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_162
timestamp 1698175906
transform 1 0 19488 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_194
timestamp 1698175906
transform 1 0 23072 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_216
timestamp 1698175906
transform 1 0 25536 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_246
timestamp 1698175906
transform 1 0 28896 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_250
timestamp 1698175906
transform 1 0 29344 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_266
timestamp 1698175906
transform 1 0 31136 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_274
timestamp 1698175906
transform 1 0 32032 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698175906
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_136
timestamp 1698175906
transform 1 0 16576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_140
timestamp 1698175906
transform 1 0 17024 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_156
timestamp 1698175906
transform 1 0 18816 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_164
timestamp 1698175906
transform 1 0 19712 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_168
timestamp 1698175906
transform 1 0 20160 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_187
timestamp 1698175906
transform 1 0 22288 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_203
timestamp 1698175906
transform 1 0 24080 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_207
timestamp 1698175906
transform 1 0 24528 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_209
timestamp 1698175906
transform 1 0 24752 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_216
timestamp 1698175906
transform 1 0 25536 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_222
timestamp 1698175906
transform 1 0 26208 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_238
timestamp 1698175906
transform 1 0 28000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698175906
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698175906
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_148
timestamp 1698175906
transform 1 0 17920 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_150
timestamp 1698175906
transform 1 0 18144 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_157
timestamp 1698175906
transform 1 0 18928 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_190
timestamp 1698175906
transform 1 0 22624 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_194
timestamp 1698175906
transform 1 0 23072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_200
timestamp 1698175906
transform 1 0 23744 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698175906
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_241
timestamp 1698175906
transform 1 0 28336 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_245
timestamp 1698175906
transform 1 0 28784 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 32368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_123
timestamp 1698175906
transform 1 0 15120 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_161
timestamp 1698175906
transform 1 0 19376 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_183
timestamp 1698175906
transform 1 0 21840 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_219
timestamp 1698175906
transform 1 0 25872 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_223
timestamp 1698175906
transform 1 0 26320 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_239
timestamp 1698175906
transform 1 0 28112 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698175906
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_173
timestamp 1698175906
transform 1 0 20720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_177
timestamp 1698175906
transform 1 0 21168 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_195
timestamp 1698175906
transform 1 0 23184 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698175906
transform 1 0 24080 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 25536 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_221
timestamp 1698175906
transform 1 0 26096 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_253
timestamp 1698175906
transform 1 0 29680 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_269
timestamp 1698175906
transform 1 0 31472 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_277
timestamp 1698175906
transform 1 0 32368 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_206
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_210
timestamp 1698175906
transform 1 0 24864 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_237
timestamp 1698175906
transform 1 0 27888 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita60_24 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 39984 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita60_25
timestamp 1698175906
transform -1 0 18704 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita60_26
timestamp 1698175906
transform -1 0 26096 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 4480 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 17472 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 37520 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 20272 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18928 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 20944 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 37520 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 37520 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 21280 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 4480 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 24976 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 20272 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 4480 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform -1 0 4480 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 37520 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 41200 16800 42000 16912 0 FreeSans 448 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 18144 41200 18256 42000 0 FreeSans 448 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 41200 17472 42000 17584 0 FreeSans 448 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 25536 41200 25648 42000 0 FreeSans 448 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 41200 24864 42000 24976 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 41200 26208 42000 26320 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 41200 20160 42000 20272 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 18816 41200 18928 42000 0 FreeSans 448 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 24864 41200 24976 42000 0 FreeSans 448 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 20160 41200 20272 42000 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 41200 16128 42000 16240 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 24248 16632 24248 16632 0 _000_
rlabel metal2 23128 26936 23128 26936 0 _001_
rlabel metal3 14112 16856 14112 16856 0 _002_
rlabel metal3 16968 26488 16968 26488 0 _003_
rlabel metal2 20440 26600 20440 26600 0 _004_
rlabel metal2 17080 14728 17080 14728 0 _005_
rlabel metal2 21056 13832 21056 13832 0 _006_
rlabel metal2 26152 24304 26152 24304 0 _007_
rlabel metal2 25816 27272 25816 27272 0 _008_
rlabel metal2 16128 15512 16128 15512 0 _009_
rlabel metal2 16072 25144 16072 25144 0 _010_
rlabel metal3 13664 23016 13664 23016 0 _011_
rlabel metal2 12600 24360 12600 24360 0 _012_
rlabel metal3 27552 18536 27552 18536 0 _013_
rlabel metal2 28840 20748 28840 20748 0 _014_
rlabel metal2 27440 16184 27440 16184 0 _015_
rlabel metal2 25648 17752 25648 17752 0 _016_
rlabel metal2 28560 22568 28560 22568 0 _017_
rlabel metal2 22792 15008 22792 15008 0 _018_
rlabel metal2 13496 15456 13496 15456 0 _019_
rlabel metal2 13888 20776 13888 20776 0 _020_
rlabel metal2 12600 19488 12600 19488 0 _021_
rlabel metal2 24584 22344 24584 22344 0 _022_
rlabel metal2 21784 24304 21784 24304 0 _023_
rlabel metal2 18872 27384 18872 27384 0 _024_
rlabel metal2 25088 15512 25088 15512 0 _025_
rlabel metal2 29176 20664 29176 20664 0 _026_
rlabel metal2 23744 26264 23744 26264 0 _027_
rlabel metal2 14840 16576 14840 16576 0 _028_
rlabel metal2 14504 17136 14504 17136 0 _029_
rlabel metal2 19656 21504 19656 21504 0 _030_
rlabel metal2 17752 23856 17752 23856 0 _031_
rlabel metal2 17528 23520 17528 23520 0 _032_
rlabel metal2 18816 23688 18816 23688 0 _033_
rlabel metal2 19208 15288 19208 15288 0 _034_
rlabel metal3 19992 23688 19992 23688 0 _035_
rlabel metal2 18648 23968 18648 23968 0 _036_
rlabel metal2 18312 23016 18312 23016 0 _037_
rlabel metal2 17080 24416 17080 24416 0 _038_
rlabel metal2 17808 24136 17808 24136 0 _039_
rlabel metal2 21056 26936 21056 26936 0 _040_
rlabel metal2 19880 15960 19880 15960 0 _041_
rlabel metal3 18480 15288 18480 15288 0 _042_
rlabel metal2 17976 18592 17976 18592 0 _043_
rlabel metal2 19880 15400 19880 15400 0 _044_
rlabel metal2 20664 15456 20664 15456 0 _045_
rlabel metal2 13608 22624 13608 22624 0 _046_
rlabel metal2 25536 26936 25536 26936 0 _047_
rlabel metal2 29904 20552 29904 20552 0 _048_
rlabel metal3 27216 23912 27216 23912 0 _049_
rlabel metal2 25816 26936 25816 26936 0 _050_
rlabel metal3 17136 15288 17136 15288 0 _051_
rlabel metal2 16968 19096 16968 19096 0 _052_
rlabel metal2 15736 24472 15736 24472 0 _053_
rlabel metal2 14112 22456 14112 22456 0 _054_
rlabel metal3 13552 23800 13552 23800 0 _055_
rlabel metal3 29064 20328 29064 20328 0 _056_
rlabel metal2 29288 21168 29288 21168 0 _057_
rlabel metal3 27160 15904 27160 15904 0 _058_
rlabel metal2 27608 16352 27608 16352 0 _059_
rlabel metal2 26152 18312 26152 18312 0 _060_
rlabel metal3 24752 18424 24752 18424 0 _061_
rlabel metal2 28672 22344 28672 22344 0 _062_
rlabel metal2 20384 23688 20384 23688 0 _063_
rlabel metal2 14168 21196 14168 21196 0 _064_
rlabel metal2 23912 15904 23912 15904 0 _065_
rlabel metal2 21448 20048 21448 20048 0 _066_
rlabel metal3 17808 20104 17808 20104 0 _067_
rlabel metal2 23800 18760 23800 18760 0 _068_
rlabel metal2 23128 17136 23128 17136 0 _069_
rlabel metal2 23352 21840 23352 21840 0 _070_
rlabel metal2 23016 22848 23016 22848 0 _071_
rlabel metal3 21448 18424 21448 18424 0 _072_
rlabel metal3 18480 18984 18480 18984 0 _073_
rlabel metal2 19880 18368 19880 18368 0 _074_
rlabel metal2 22792 17808 22792 17808 0 _075_
rlabel metal2 19880 22848 19880 22848 0 _076_
rlabel metal2 14392 19152 14392 19152 0 _077_
rlabel metal2 18760 16520 18760 16520 0 _078_
rlabel metal2 27160 18144 27160 18144 0 _079_
rlabel metal2 23016 15960 23016 15960 0 _080_
rlabel metal2 14000 16072 14000 16072 0 _081_
rlabel metal2 23016 21952 23016 21952 0 _082_
rlabel metal2 15064 24360 15064 24360 0 _083_
rlabel metal2 18760 21448 18760 21448 0 _084_
rlabel metal2 14728 21448 14728 21448 0 _085_
rlabel metal2 13944 20356 13944 20356 0 _086_
rlabel metal2 15176 16464 15176 16464 0 _087_
rlabel metal2 14168 19096 14168 19096 0 _088_
rlabel metal2 13216 19096 13216 19096 0 _089_
rlabel metal3 24136 23352 24136 23352 0 _090_
rlabel metal2 21896 22344 21896 22344 0 _091_
rlabel metal3 28280 20104 28280 20104 0 _092_
rlabel metal2 19656 23240 19656 23240 0 _093_
rlabel metal2 19264 25368 19264 25368 0 _094_
rlabel metal2 23464 25816 23464 25816 0 _095_
rlabel metal2 28280 22232 28280 22232 0 _096_
rlabel metal2 16296 22064 16296 22064 0 _097_
rlabel metal2 23912 22288 23912 22288 0 _098_
rlabel metal2 17640 21056 17640 21056 0 _099_
rlabel metal2 18592 23128 18592 23128 0 _100_
rlabel metal2 26936 23968 26936 23968 0 _101_
rlabel metal3 20944 26824 20944 26824 0 _102_
rlabel metal2 19208 27160 19208 27160 0 _103_
rlabel metal2 25928 20440 25928 20440 0 _104_
rlabel metal3 2478 26936 2478 26936 0 clk
rlabel metal2 23352 20440 23352 20440 0 clknet_0_clk
rlabel metal2 15008 23688 15008 23688 0 clknet_1_0__leaf_clk
rlabel metal3 23800 27048 23800 27048 0 clknet_1_1__leaf_clk
rlabel metal2 16072 18704 16072 18704 0 dut60.count\[0\]
rlabel metal2 14392 19936 14392 19936 0 dut60.count\[1\]
rlabel metal2 21952 19432 21952 19432 0 dut60.count\[2\]
rlabel metal2 20664 23072 20664 23072 0 dut60.count\[3\]
rlabel metal3 6356 23128 6356 23128 0 net1
rlabel metal2 27944 24192 27944 24192 0 net10
rlabel metal2 28168 25760 28168 25760 0 net11
rlabel metal3 22008 26936 22008 26936 0 net12
rlabel metal2 30296 20356 30296 20356 0 net13
rlabel metal3 30296 20776 30296 20776 0 net14
rlabel metal2 18088 34972 18088 34972 0 net15
rlabel metal2 4312 16800 4312 16800 0 net16
rlabel metal2 25144 27832 25144 27832 0 net17
rlabel metal2 20552 32480 20552 32480 0 net18
rlabel metal2 4312 24640 4312 24640 0 net19
rlabel metal2 17696 13048 17696 13048 0 net2
rlabel metal2 11312 15176 11312 15176 0 net20
rlabel metal2 30744 23464 30744 23464 0 net21
rlabel metal2 24584 5964 24584 5964 0 net22
rlabel metal2 37688 15736 37688 15736 0 net23
rlabel metal3 40754 19544 40754 19544 0 net24
rlabel metal2 18200 2590 18200 2590 0 net25
rlabel metal2 25704 37464 25704 37464 0 net26
rlabel metal2 13496 25536 13496 25536 0 net3
rlabel metal2 27832 17808 27832 17808 0 net4
rlabel metal2 37912 16352 37912 16352 0 net5
rlabel metal2 18648 27328 18648 27328 0 net6
rlabel metal2 29624 17192 29624 17192 0 net7
rlabel metal2 19152 14616 19152 14616 0 net8
rlabel metal2 21112 8512 21112 8512 0 net9
rlabel metal3 1358 22904 1358 22904 0 segm[10]
rlabel metal2 17528 2198 17528 2198 0 segm[11]
rlabel metal3 1358 24920 1358 24920 0 segm[12]
rlabel metal3 40642 18200 40642 18200 0 segm[13]
rlabel metal2 40040 16800 40040 16800 0 segm[1]
rlabel metal2 18200 39298 18200 39298 0 segm[2]
rlabel metal2 40040 17640 40040 17640 0 segm[4]
rlabel metal2 18872 2422 18872 2422 0 segm[6]
rlabel metal2 20888 2198 20888 2198 0 segm[7]
rlabel metal2 40040 25256 40040 25256 0 segm[8]
rlabel metal2 40040 26712 40040 26712 0 segm[9]
rlabel metal2 22232 39746 22232 39746 0 sel[0]
rlabel metal2 39816 20552 39816 20552 0 sel[10]
rlabel metal2 40040 21112 40040 21112 0 sel[11]
rlabel metal2 18872 39690 18872 39690 0 sel[1]
rlabel metal3 1358 16184 1358 16184 0 sel[2]
rlabel metal2 24920 39746 24920 39746 0 sel[3]
rlabel metal2 20216 39354 20216 39354 0 sel[4]
rlabel metal3 1358 24248 1358 24248 0 sel[5]
rlabel metal3 1358 16856 1358 16856 0 sel[6]
rlabel metal2 40040 23800 40040 23800 0 sel[7]
rlabel metal2 24248 2198 24248 2198 0 sel[8]
rlabel metal3 40642 16184 40642 16184 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
