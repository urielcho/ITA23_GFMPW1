magic
tech gf180mcuD
magscale 1 10
timestamp 1699643243
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 18062 38274 18114 38286
rect 18062 38210 18114 38222
rect 22430 38274 22482 38286
rect 22430 38210 22482 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 17042 37998 17054 38050
rect 17106 37998 17118 38050
rect 21746 37998 21758 38050
rect 21810 37998 21822 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 19854 37490 19906 37502
rect 19854 37426 19906 37438
rect 22766 37490 22818 37502
rect 22766 37426 22818 37438
rect 26798 37490 26850 37502
rect 26798 37426 26850 37438
rect 18834 37214 18846 37266
rect 18898 37214 18910 37266
rect 22082 37214 22094 37266
rect 22146 37214 22158 37266
rect 25778 37214 25790 37266
rect 25842 37214 25854 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 19170 29374 19182 29426
rect 19234 29374 19246 29426
rect 22542 29314 22594 29326
rect 19842 29262 19854 29314
rect 19906 29262 19918 29314
rect 21970 29262 21982 29314
rect 22034 29262 22046 29314
rect 22542 29250 22594 29262
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 15150 28642 15202 28654
rect 15150 28578 15202 28590
rect 18510 28642 18562 28654
rect 21970 28590 21982 28642
rect 22034 28590 22046 28642
rect 18510 28578 18562 28590
rect 15262 28530 15314 28542
rect 15262 28466 15314 28478
rect 18734 28530 18786 28542
rect 18734 28466 18786 28478
rect 18846 28530 18898 28542
rect 21746 28478 21758 28530
rect 21810 28478 21822 28530
rect 18846 28466 18898 28478
rect 17166 28418 17218 28430
rect 17166 28354 17218 28366
rect 17614 28418 17666 28430
rect 17614 28354 17666 28366
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 14354 27918 14366 27970
rect 14418 27918 14430 27970
rect 25342 27858 25394 27870
rect 13682 27806 13694 27858
rect 13746 27806 13758 27858
rect 17378 27806 17390 27858
rect 17442 27806 17454 27858
rect 21634 27806 21646 27858
rect 21698 27806 21710 27858
rect 25342 27794 25394 27806
rect 16482 27694 16494 27746
rect 16546 27694 16558 27746
rect 18162 27694 18174 27746
rect 18226 27694 18238 27746
rect 20290 27694 20302 27746
rect 20354 27694 20366 27746
rect 22418 27694 22430 27746
rect 22482 27694 22494 27746
rect 24546 27694 24558 27746
rect 24610 27694 24622 27746
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 15486 27298 15538 27310
rect 15486 27234 15538 27246
rect 19966 27298 20018 27310
rect 19966 27234 20018 27246
rect 15822 27186 15874 27198
rect 15822 27122 15874 27134
rect 16494 27186 16546 27198
rect 19630 27186 19682 27198
rect 17378 27134 17390 27186
rect 17442 27134 17454 27186
rect 16494 27122 16546 27134
rect 19630 27122 19682 27134
rect 22094 27186 22146 27198
rect 26126 27186 26178 27198
rect 25666 27134 25678 27186
rect 25730 27134 25742 27186
rect 22094 27122 22146 27134
rect 26126 27122 26178 27134
rect 40014 27186 40066 27198
rect 40014 27122 40066 27134
rect 16606 27074 16658 27086
rect 16606 27010 16658 27022
rect 17054 27074 17106 27086
rect 18398 27074 18450 27086
rect 17490 27022 17502 27074
rect 17554 27022 17566 27074
rect 17054 27010 17106 27022
rect 18398 27010 18450 27022
rect 18734 27074 18786 27086
rect 18734 27010 18786 27022
rect 18846 27074 18898 27086
rect 19518 27074 19570 27086
rect 19170 27022 19182 27074
rect 19234 27022 19246 27074
rect 20290 27022 20302 27074
rect 20354 27022 20366 27074
rect 22754 27022 22766 27074
rect 22818 27022 22830 27074
rect 37650 27022 37662 27074
rect 37714 27022 37726 27074
rect 18846 27010 18898 27022
rect 19518 27010 19570 27022
rect 16046 26962 16098 26974
rect 16046 26898 16098 26910
rect 16382 26962 16434 26974
rect 16382 26898 16434 26910
rect 18062 26962 18114 26974
rect 21982 26962 22034 26974
rect 19730 26910 19742 26962
rect 19794 26910 19806 26962
rect 18062 26898 18114 26910
rect 21982 26898 22034 26910
rect 22206 26962 22258 26974
rect 22206 26898 22258 26910
rect 22430 26962 22482 26974
rect 23538 26910 23550 26962
rect 23602 26910 23614 26962
rect 22430 26898 22482 26910
rect 18510 26850 18562 26862
rect 18510 26786 18562 26798
rect 21870 26850 21922 26862
rect 21870 26786 21922 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 18174 26514 18226 26526
rect 18174 26450 18226 26462
rect 21422 26514 21474 26526
rect 21422 26450 21474 26462
rect 23550 26514 23602 26526
rect 23550 26450 23602 26462
rect 24446 26514 24498 26526
rect 24446 26450 24498 26462
rect 19070 26290 19122 26302
rect 4274 26238 4286 26290
rect 4338 26238 4350 26290
rect 14578 26238 14590 26290
rect 14642 26238 14654 26290
rect 18834 26238 18846 26290
rect 18898 26238 18910 26290
rect 19070 26226 19122 26238
rect 19294 26290 19346 26302
rect 19294 26226 19346 26238
rect 23438 26290 23490 26302
rect 23438 26226 23490 26238
rect 23662 26290 23714 26302
rect 23662 26226 23714 26238
rect 23998 26290 24050 26302
rect 23998 26226 24050 26238
rect 24334 26290 24386 26302
rect 25554 26238 25566 26290
rect 25618 26238 25630 26290
rect 24334 26226 24386 26238
rect 15150 26178 15202 26190
rect 11778 26126 11790 26178
rect 11842 26126 11854 26178
rect 13906 26126 13918 26178
rect 13970 26126 13982 26178
rect 15150 26114 15202 26126
rect 18062 26178 18114 26190
rect 28926 26178 28978 26190
rect 21298 26126 21310 26178
rect 21362 26126 21374 26178
rect 26338 26126 26350 26178
rect 26402 26126 26414 26178
rect 28466 26126 28478 26178
rect 28530 26126 28542 26178
rect 18062 26114 18114 26126
rect 28926 26114 28978 26126
rect 1934 26066 1986 26078
rect 1934 26002 1986 26014
rect 17950 26066 18002 26078
rect 17950 26002 18002 26014
rect 19406 26066 19458 26078
rect 19406 26002 19458 26014
rect 21646 26066 21698 26078
rect 21646 26002 21698 26014
rect 24446 26066 24498 26078
rect 24446 26002 24498 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 15822 25730 15874 25742
rect 15822 25666 15874 25678
rect 24446 25618 24498 25630
rect 24446 25554 24498 25566
rect 25790 25618 25842 25630
rect 25790 25554 25842 25566
rect 40014 25618 40066 25630
rect 40014 25554 40066 25566
rect 14814 25506 14866 25518
rect 15486 25506 15538 25518
rect 15250 25454 15262 25506
rect 15314 25454 15326 25506
rect 14814 25442 14866 25454
rect 15486 25442 15538 25454
rect 15710 25506 15762 25518
rect 21310 25506 21362 25518
rect 18274 25454 18286 25506
rect 18338 25454 18350 25506
rect 15710 25442 15762 25454
rect 21310 25442 21362 25454
rect 24670 25506 24722 25518
rect 24670 25442 24722 25454
rect 25902 25506 25954 25518
rect 37650 25454 37662 25506
rect 37714 25454 37726 25506
rect 25902 25442 25954 25454
rect 14702 25394 14754 25406
rect 14702 25330 14754 25342
rect 14926 25394 14978 25406
rect 14926 25330 14978 25342
rect 17502 25394 17554 25406
rect 17502 25330 17554 25342
rect 17838 25394 17890 25406
rect 24334 25394 24386 25406
rect 18498 25342 18510 25394
rect 18562 25342 18574 25394
rect 17838 25330 17890 25342
rect 24334 25330 24386 25342
rect 24894 25394 24946 25406
rect 24894 25330 24946 25342
rect 26126 25394 26178 25406
rect 26126 25330 26178 25342
rect 27246 25394 27298 25406
rect 27246 25330 27298 25342
rect 27470 25394 27522 25406
rect 27470 25330 27522 25342
rect 27582 25394 27634 25406
rect 27582 25330 27634 25342
rect 21422 25282 21474 25294
rect 21422 25218 21474 25230
rect 21646 25282 21698 25294
rect 21646 25218 21698 25230
rect 25566 25282 25618 25294
rect 25566 25218 25618 25230
rect 25678 25282 25730 25294
rect 25678 25218 25730 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 18286 24946 18338 24958
rect 16482 24894 16494 24946
rect 16546 24894 16558 24946
rect 18286 24882 18338 24894
rect 26462 24946 26514 24958
rect 26462 24882 26514 24894
rect 23998 24834 24050 24846
rect 18610 24782 18622 24834
rect 18674 24782 18686 24834
rect 23998 24770 24050 24782
rect 26910 24834 26962 24846
rect 26910 24770 26962 24782
rect 30942 24834 30994 24846
rect 30942 24770 30994 24782
rect 17838 24722 17890 24734
rect 16706 24670 16718 24722
rect 16770 24670 16782 24722
rect 17378 24670 17390 24722
rect 17442 24670 17454 24722
rect 17838 24658 17890 24670
rect 24334 24722 24386 24734
rect 24334 24658 24386 24670
rect 24558 24722 24610 24734
rect 24558 24658 24610 24670
rect 27022 24722 27074 24734
rect 27346 24670 27358 24722
rect 27410 24670 27422 24722
rect 30706 24670 30718 24722
rect 30770 24670 30782 24722
rect 37650 24670 37662 24722
rect 37714 24670 37726 24722
rect 27022 24658 27074 24670
rect 24110 24610 24162 24622
rect 28130 24558 28142 24610
rect 28194 24558 28206 24610
rect 30258 24558 30270 24610
rect 30322 24558 30334 24610
rect 24110 24546 24162 24558
rect 17614 24498 17666 24510
rect 17614 24434 17666 24446
rect 17950 24498 18002 24510
rect 17950 24434 18002 24446
rect 26910 24498 26962 24510
rect 26910 24434 26962 24446
rect 40014 24498 40066 24510
rect 40014 24434 40066 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 28030 24162 28082 24174
rect 28030 24098 28082 24110
rect 16942 24050 16994 24062
rect 26126 24050 26178 24062
rect 25666 23998 25678 24050
rect 25730 23998 25742 24050
rect 16942 23986 16994 23998
rect 26126 23986 26178 23998
rect 26686 24050 26738 24062
rect 26686 23986 26738 23998
rect 29262 24050 29314 24062
rect 29262 23986 29314 23998
rect 40014 24050 40066 24062
rect 40014 23986 40066 23998
rect 16158 23938 16210 23950
rect 16158 23874 16210 23886
rect 16606 23938 16658 23950
rect 16606 23874 16658 23886
rect 21982 23938 22034 23950
rect 28142 23938 28194 23950
rect 22754 23886 22766 23938
rect 22818 23886 22830 23938
rect 21982 23874 22034 23886
rect 28142 23874 28194 23886
rect 29038 23938 29090 23950
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 29038 23874 29090 23886
rect 17278 23826 17330 23838
rect 17278 23762 17330 23774
rect 21310 23826 21362 23838
rect 28030 23826 28082 23838
rect 23538 23774 23550 23826
rect 23602 23774 23614 23826
rect 21310 23762 21362 23774
rect 28030 23762 28082 23774
rect 29598 23826 29650 23838
rect 29598 23762 29650 23774
rect 17614 23714 17666 23726
rect 17614 23650 17666 23662
rect 21422 23714 21474 23726
rect 21422 23650 21474 23662
rect 21534 23714 21586 23726
rect 21534 23650 21586 23662
rect 29374 23714 29426 23726
rect 29374 23650 29426 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 21086 23378 21138 23390
rect 16482 23326 16494 23378
rect 16546 23326 16558 23378
rect 21086 23314 21138 23326
rect 21982 23378 22034 23390
rect 21982 23314 22034 23326
rect 23662 23378 23714 23390
rect 23662 23314 23714 23326
rect 23886 23378 23938 23390
rect 23886 23314 23938 23326
rect 23998 23378 24050 23390
rect 23998 23314 24050 23326
rect 24110 23378 24162 23390
rect 26450 23326 26462 23378
rect 26514 23326 26526 23378
rect 24110 23314 24162 23326
rect 15934 23266 15986 23278
rect 19742 23266 19794 23278
rect 21646 23266 21698 23278
rect 12562 23214 12574 23266
rect 12626 23214 12638 23266
rect 17378 23214 17390 23266
rect 17442 23214 17454 23266
rect 17714 23214 17726 23266
rect 17778 23214 17790 23266
rect 20402 23214 20414 23266
rect 20466 23214 20478 23266
rect 15934 23202 15986 23214
rect 19742 23202 19794 23214
rect 21646 23202 21698 23214
rect 22094 23266 22146 23278
rect 27794 23214 27806 23266
rect 27858 23214 27870 23266
rect 22094 23202 22146 23214
rect 15598 23154 15650 23166
rect 11890 23102 11902 23154
rect 11954 23102 11966 23154
rect 15598 23090 15650 23102
rect 16046 23154 16098 23166
rect 16046 23090 16098 23102
rect 16830 23154 16882 23166
rect 19406 23154 19458 23166
rect 18050 23102 18062 23154
rect 18114 23102 18126 23154
rect 16830 23090 16882 23102
rect 19406 23090 19458 23102
rect 20078 23154 20130 23166
rect 20078 23090 20130 23102
rect 21870 23154 21922 23166
rect 21870 23090 21922 23102
rect 26126 23154 26178 23166
rect 27010 23102 27022 23154
rect 27074 23102 27086 23154
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 26126 23090 26178 23102
rect 15150 23042 15202 23054
rect 14690 22990 14702 23042
rect 14754 22990 14766 23042
rect 15150 22978 15202 22990
rect 15710 23042 15762 23054
rect 15710 22978 15762 22990
rect 18398 23042 18450 23054
rect 21186 22990 21198 23042
rect 21250 22990 21262 23042
rect 29922 22990 29934 23042
rect 29986 22990 29998 23042
rect 18398 22978 18450 22990
rect 18622 22930 18674 22942
rect 18622 22866 18674 22878
rect 18958 22930 19010 22942
rect 18958 22866 19010 22878
rect 20862 22930 20914 22942
rect 20862 22866 20914 22878
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 18286 22594 18338 22606
rect 18286 22530 18338 22542
rect 19966 22594 20018 22606
rect 19966 22530 20018 22542
rect 28254 22594 28306 22606
rect 28254 22530 28306 22542
rect 16158 22482 16210 22494
rect 40014 22482 40066 22494
rect 24882 22430 24894 22482
rect 24946 22430 24958 22482
rect 16158 22418 16210 22430
rect 40014 22418 40066 22430
rect 20414 22370 20466 22382
rect 14802 22318 14814 22370
rect 14866 22318 14878 22370
rect 16370 22318 16382 22370
rect 16434 22318 16446 22370
rect 17714 22318 17726 22370
rect 17778 22318 17790 22370
rect 19618 22318 19630 22370
rect 19682 22318 19694 22370
rect 20414 22306 20466 22318
rect 21534 22370 21586 22382
rect 23874 22318 23886 22370
rect 23938 22318 23950 22370
rect 24210 22318 24222 22370
rect 24274 22318 24286 22370
rect 25218 22318 25230 22370
rect 25282 22318 25294 22370
rect 28354 22318 28366 22370
rect 28418 22318 28430 22370
rect 37874 22318 37886 22370
rect 37938 22318 37950 22370
rect 21534 22306 21586 22318
rect 16046 22258 16098 22270
rect 21310 22258 21362 22270
rect 23214 22258 23266 22270
rect 17042 22206 17054 22258
rect 17106 22206 17118 22258
rect 17490 22206 17502 22258
rect 17554 22206 17566 22258
rect 22194 22206 22206 22258
rect 22258 22206 22270 22258
rect 16046 22194 16098 22206
rect 21310 22194 21362 22206
rect 23214 22194 23266 22206
rect 26686 22258 26738 22270
rect 28142 22258 28194 22270
rect 27010 22206 27022 22258
rect 27074 22206 27086 22258
rect 26686 22194 26738 22206
rect 28142 22194 28194 22206
rect 28590 22258 28642 22270
rect 28590 22194 28642 22206
rect 15374 22146 15426 22158
rect 16718 22146 16770 22158
rect 15026 22094 15038 22146
rect 15090 22094 15102 22146
rect 15698 22094 15710 22146
rect 15762 22094 15774 22146
rect 15374 22082 15426 22094
rect 16718 22082 16770 22094
rect 18622 22146 18674 22158
rect 18622 22082 18674 22094
rect 19294 22146 19346 22158
rect 19294 22082 19346 22094
rect 19406 22146 19458 22158
rect 19406 22082 19458 22094
rect 19518 22146 19570 22158
rect 22542 22146 22594 22158
rect 20738 22094 20750 22146
rect 20802 22094 20814 22146
rect 21858 22094 21870 22146
rect 21922 22094 21934 22146
rect 22866 22094 22878 22146
rect 22930 22094 22942 22146
rect 19518 22082 19570 22094
rect 22542 22082 22594 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 17390 21810 17442 21822
rect 16370 21758 16382 21810
rect 16434 21758 16446 21810
rect 17390 21746 17442 21758
rect 17950 21810 18002 21822
rect 17950 21746 18002 21758
rect 25342 21810 25394 21822
rect 25342 21746 25394 21758
rect 25454 21810 25506 21822
rect 25454 21746 25506 21758
rect 26910 21810 26962 21822
rect 26910 21746 26962 21758
rect 15934 21698 15986 21710
rect 12562 21646 12574 21698
rect 12626 21646 12638 21698
rect 15934 21634 15986 21646
rect 16718 21698 16770 21710
rect 16718 21634 16770 21646
rect 16830 21698 16882 21710
rect 16830 21634 16882 21646
rect 17502 21698 17554 21710
rect 17502 21634 17554 21646
rect 15710 21586 15762 21598
rect 11890 21534 11902 21586
rect 11954 21534 11966 21586
rect 15710 21522 15762 21534
rect 15822 21586 15874 21598
rect 15822 21522 15874 21534
rect 17838 21586 17890 21598
rect 17838 21522 17890 21534
rect 18174 21586 18226 21598
rect 18174 21522 18226 21534
rect 18622 21586 18674 21598
rect 18946 21534 18958 21586
rect 19010 21534 19022 21586
rect 27234 21534 27246 21586
rect 27298 21534 27310 21586
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 18622 21522 18674 21534
rect 15150 21474 15202 21486
rect 37438 21474 37490 21486
rect 14690 21422 14702 21474
rect 14754 21422 14766 21474
rect 22642 21422 22654 21474
rect 22706 21422 22718 21474
rect 28018 21422 28030 21474
rect 28082 21422 28094 21474
rect 30146 21422 30158 21474
rect 30210 21422 30222 21474
rect 39890 21422 39902 21474
rect 39954 21422 39966 21474
rect 15150 21410 15202 21422
rect 37438 21410 37490 21422
rect 25230 21362 25282 21374
rect 25230 21298 25282 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 1934 20914 1986 20926
rect 13582 20914 13634 20926
rect 29262 20914 29314 20926
rect 9986 20862 9998 20914
rect 10050 20862 10062 20914
rect 15362 20862 15374 20914
rect 15426 20862 15438 20914
rect 22306 20862 22318 20914
rect 22370 20862 22382 20914
rect 1934 20850 1986 20862
rect 13582 20850 13634 20862
rect 29262 20850 29314 20862
rect 40014 20914 40066 20926
rect 40014 20850 40066 20862
rect 28142 20802 28194 20814
rect 4274 20750 4286 20802
rect 4338 20750 4350 20802
rect 12898 20750 12910 20802
rect 12962 20750 12974 20802
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 21970 20750 21982 20802
rect 22034 20750 22046 20802
rect 22642 20750 22654 20802
rect 22706 20750 22718 20802
rect 28142 20738 28194 20750
rect 28478 20802 28530 20814
rect 28478 20738 28530 20750
rect 29038 20802 29090 20814
rect 29362 20750 29374 20802
rect 29426 20750 29438 20802
rect 37874 20750 37886 20802
rect 37938 20750 37950 20802
rect 29038 20738 29090 20750
rect 21758 20690 21810 20702
rect 29598 20690 29650 20702
rect 12114 20638 12126 20690
rect 12178 20638 12190 20690
rect 22082 20638 22094 20690
rect 22146 20638 22158 20690
rect 26786 20638 26798 20690
rect 26850 20638 26862 20690
rect 21758 20626 21810 20638
rect 29598 20626 29650 20638
rect 21534 20578 21586 20590
rect 21534 20514 21586 20526
rect 28366 20578 28418 20590
rect 28366 20514 28418 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 11902 20242 11954 20254
rect 11902 20178 11954 20190
rect 17614 20242 17666 20254
rect 17614 20178 17666 20190
rect 22878 20242 22930 20254
rect 22878 20178 22930 20190
rect 15822 20130 15874 20142
rect 15822 20066 15874 20078
rect 17726 20130 17778 20142
rect 21534 20130 21586 20142
rect 19506 20078 19518 20130
rect 19570 20078 19582 20130
rect 20962 20078 20974 20130
rect 21026 20078 21038 20130
rect 17726 20066 17778 20078
rect 21534 20066 21586 20078
rect 22206 20130 22258 20142
rect 22206 20066 22258 20078
rect 23438 20130 23490 20142
rect 23438 20066 23490 20078
rect 27134 20130 27186 20142
rect 27134 20066 27186 20078
rect 28366 20130 28418 20142
rect 28366 20066 28418 20078
rect 28478 20130 28530 20142
rect 29698 20078 29710 20130
rect 29762 20078 29774 20130
rect 28478 20066 28530 20078
rect 12238 20018 12290 20030
rect 20302 20018 20354 20030
rect 22766 20018 22818 20030
rect 17378 19966 17390 20018
rect 17442 19966 17454 20018
rect 20066 19966 20078 20018
rect 20130 19966 20142 20018
rect 20402 19966 20414 20018
rect 20466 19966 20478 20018
rect 12238 19954 12290 19966
rect 20302 19954 20354 19966
rect 22766 19954 22818 19966
rect 23102 20018 23154 20030
rect 23102 19954 23154 19966
rect 27358 20018 27410 20030
rect 27358 19954 27410 19966
rect 27806 20018 27858 20030
rect 27806 19954 27858 19966
rect 28142 20018 28194 20030
rect 28142 19954 28194 19966
rect 29374 20018 29426 20030
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 29374 19954 29426 19966
rect 22430 19906 22482 19918
rect 21410 19854 21422 19906
rect 21474 19854 21486 19906
rect 22082 19854 22094 19906
rect 22146 19854 22158 19906
rect 22430 19842 22482 19854
rect 27582 19906 27634 19918
rect 27582 19842 27634 19854
rect 15710 19794 15762 19806
rect 15710 19730 15762 19742
rect 16046 19794 16098 19806
rect 16046 19730 16098 19742
rect 21758 19794 21810 19806
rect 21758 19730 21810 19742
rect 40014 19794 40066 19806
rect 40014 19730 40066 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 15822 19458 15874 19470
rect 14690 19406 14702 19458
rect 14754 19406 14766 19458
rect 15822 19394 15874 19406
rect 15598 19346 15650 19358
rect 15598 19282 15650 19294
rect 16158 19346 16210 19358
rect 16158 19282 16210 19294
rect 16606 19346 16658 19358
rect 22430 19346 22482 19358
rect 40014 19346 40066 19358
rect 19618 19294 19630 19346
rect 19682 19294 19694 19346
rect 23986 19294 23998 19346
rect 24050 19294 24062 19346
rect 26114 19294 26126 19346
rect 26178 19294 26190 19346
rect 16606 19282 16658 19294
rect 22430 19282 22482 19294
rect 40014 19282 40066 19294
rect 14142 19234 14194 19246
rect 14142 19170 14194 19182
rect 14366 19234 14418 19246
rect 14366 19170 14418 19182
rect 17278 19234 17330 19246
rect 17278 19170 17330 19182
rect 18622 19234 18674 19246
rect 22318 19234 22370 19246
rect 19282 19182 19294 19234
rect 19346 19182 19358 19234
rect 20178 19182 20190 19234
rect 20242 19182 20254 19234
rect 18622 19170 18674 19182
rect 22318 19170 22370 19182
rect 22542 19234 22594 19246
rect 22542 19170 22594 19182
rect 22766 19234 22818 19246
rect 23314 19182 23326 19234
rect 23378 19182 23390 19234
rect 27906 19182 27918 19234
rect 27970 19182 27982 19234
rect 37650 19182 37662 19234
rect 37714 19182 37726 19234
rect 22766 19170 22818 19182
rect 19058 19070 19070 19122
rect 19122 19070 19134 19122
rect 16494 19010 16546 19022
rect 18510 19010 18562 19022
rect 16930 18958 16942 19010
rect 16994 18958 17006 19010
rect 16494 18946 16546 18958
rect 18510 18946 18562 18958
rect 26574 19010 26626 19022
rect 28130 18958 28142 19010
rect 28194 18958 28206 19010
rect 26574 18946 26626 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 14590 18674 14642 18686
rect 15822 18674 15874 18686
rect 14914 18622 14926 18674
rect 14978 18622 14990 18674
rect 14590 18610 14642 18622
rect 15822 18610 15874 18622
rect 16046 18674 16098 18686
rect 16046 18610 16098 18622
rect 22094 18674 22146 18686
rect 25230 18674 25282 18686
rect 23538 18622 23550 18674
rect 23602 18622 23614 18674
rect 22094 18610 22146 18622
rect 25230 18610 25282 18622
rect 25454 18674 25506 18686
rect 25454 18610 25506 18622
rect 21870 18562 21922 18574
rect 11666 18510 11678 18562
rect 11730 18510 11742 18562
rect 19170 18510 19182 18562
rect 19234 18510 19246 18562
rect 19618 18510 19630 18562
rect 19682 18510 19694 18562
rect 21186 18510 21198 18562
rect 21250 18510 21262 18562
rect 23090 18510 23102 18562
rect 23154 18510 23166 18562
rect 23314 18510 23326 18562
rect 23378 18510 23390 18562
rect 27794 18510 27806 18562
rect 27858 18510 27870 18562
rect 21870 18498 21922 18510
rect 17950 18450 18002 18462
rect 10994 18398 11006 18450
rect 11058 18398 11070 18450
rect 15586 18398 15598 18450
rect 15650 18398 15662 18450
rect 16258 18398 16270 18450
rect 16322 18398 16334 18450
rect 17950 18386 18002 18398
rect 18510 18450 18562 18462
rect 21534 18450 21586 18462
rect 25902 18450 25954 18462
rect 18946 18398 18958 18450
rect 19010 18398 19022 18450
rect 19506 18398 19518 18450
rect 19570 18398 19582 18450
rect 20626 18398 20638 18450
rect 20690 18398 20702 18450
rect 22866 18398 22878 18450
rect 22930 18398 22942 18450
rect 27010 18398 27022 18450
rect 27074 18398 27086 18450
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 18510 18386 18562 18398
rect 21534 18386 21586 18398
rect 25902 18386 25954 18398
rect 14254 18338 14306 18350
rect 13794 18286 13806 18338
rect 13858 18286 13870 18338
rect 14254 18274 14306 18286
rect 15934 18338 15986 18350
rect 25342 18338 25394 18350
rect 17490 18286 17502 18338
rect 17554 18286 17566 18338
rect 20290 18286 20302 18338
rect 20354 18286 20366 18338
rect 15934 18274 15986 18286
rect 25342 18274 25394 18286
rect 26686 18338 26738 18350
rect 29922 18286 29934 18338
rect 29986 18286 29998 18338
rect 26686 18274 26738 18286
rect 18398 18226 18450 18238
rect 18398 18162 18450 18174
rect 22206 18226 22258 18238
rect 22206 18162 22258 18174
rect 40014 18226 40066 18238
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 18062 17890 18114 17902
rect 18062 17826 18114 17838
rect 22878 17890 22930 17902
rect 22878 17826 22930 17838
rect 17054 17778 17106 17790
rect 22654 17778 22706 17790
rect 40014 17778 40066 17790
rect 10770 17726 10782 17778
rect 10834 17726 10846 17778
rect 12898 17726 12910 17778
rect 12962 17726 12974 17778
rect 21858 17726 21870 17778
rect 21922 17726 21934 17778
rect 28242 17726 28254 17778
rect 28306 17726 28318 17778
rect 17054 17714 17106 17726
rect 22654 17714 22706 17726
rect 40014 17714 40066 17726
rect 14478 17666 14530 17678
rect 20862 17666 20914 17678
rect 10098 17614 10110 17666
rect 10162 17614 10174 17666
rect 16258 17614 16270 17666
rect 16322 17614 16334 17666
rect 17154 17614 17166 17666
rect 17218 17614 17230 17666
rect 18274 17614 18286 17666
rect 18338 17614 18350 17666
rect 18498 17614 18510 17666
rect 18562 17614 18574 17666
rect 19506 17614 19518 17666
rect 19570 17614 19582 17666
rect 14478 17602 14530 17614
rect 20862 17602 20914 17614
rect 21534 17666 21586 17678
rect 23886 17666 23938 17678
rect 22082 17614 22094 17666
rect 22146 17614 22158 17666
rect 23762 17614 23774 17666
rect 23826 17614 23838 17666
rect 21534 17602 21586 17614
rect 23886 17602 23938 17614
rect 23998 17666 24050 17678
rect 23998 17602 24050 17614
rect 24334 17666 24386 17678
rect 25330 17614 25342 17666
rect 25394 17614 25406 17666
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 24334 17602 24386 17614
rect 14814 17554 14866 17566
rect 19406 17554 19458 17566
rect 20526 17554 20578 17566
rect 16482 17502 16494 17554
rect 16546 17502 16558 17554
rect 18610 17502 18622 17554
rect 18674 17502 18686 17554
rect 20066 17502 20078 17554
rect 20130 17502 20142 17554
rect 14814 17490 14866 17502
rect 19406 17490 19458 17502
rect 20526 17490 20578 17502
rect 21646 17554 21698 17566
rect 21646 17490 21698 17502
rect 24222 17554 24274 17566
rect 26114 17502 26126 17554
rect 26178 17502 26190 17554
rect 24222 17490 24274 17502
rect 13582 17442 13634 17454
rect 15822 17442 15874 17454
rect 15474 17390 15486 17442
rect 15538 17390 15550 17442
rect 13582 17378 13634 17390
rect 15822 17378 15874 17390
rect 20638 17442 20690 17454
rect 20638 17378 20690 17390
rect 21870 17442 21922 17454
rect 29262 17442 29314 17454
rect 23202 17390 23214 17442
rect 23266 17390 23278 17442
rect 21870 17378 21922 17390
rect 29262 17378 29314 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 19294 17106 19346 17118
rect 20190 17106 20242 17118
rect 21758 17106 21810 17118
rect 19618 17054 19630 17106
rect 19682 17054 19694 17106
rect 21186 17054 21198 17106
rect 21250 17054 21262 17106
rect 19294 17042 19346 17054
rect 20190 17042 20242 17054
rect 21758 17042 21810 17054
rect 21982 17106 22034 17118
rect 21982 17042 22034 17054
rect 22094 17106 22146 17118
rect 22094 17042 22146 17054
rect 22990 17106 23042 17118
rect 22990 17042 23042 17054
rect 15486 16994 15538 17006
rect 15486 16930 15538 16942
rect 15710 16994 15762 17006
rect 15710 16930 15762 16942
rect 15934 16994 15986 17006
rect 15934 16930 15986 16942
rect 19966 16994 20018 17006
rect 19966 16930 20018 16942
rect 22766 16994 22818 17006
rect 24334 16994 24386 17006
rect 24098 16942 24110 16994
rect 24162 16942 24174 16994
rect 22766 16930 22818 16942
rect 24334 16930 24386 16942
rect 15262 16882 15314 16894
rect 15262 16818 15314 16830
rect 20638 16882 20690 16894
rect 20638 16818 20690 16830
rect 20862 16882 20914 16894
rect 23102 16882 23154 16894
rect 21522 16830 21534 16882
rect 21586 16830 21598 16882
rect 22530 16830 22542 16882
rect 22594 16830 22606 16882
rect 23538 16830 23550 16882
rect 23602 16830 23614 16882
rect 20862 16818 20914 16830
rect 23102 16818 23154 16830
rect 22878 16770 22930 16782
rect 20290 16718 20302 16770
rect 20354 16718 20366 16770
rect 22878 16706 22930 16718
rect 24222 16770 24274 16782
rect 24222 16706 24274 16718
rect 23762 16606 23774 16658
rect 23826 16606 23838 16658
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 15262 16322 15314 16334
rect 15262 16258 15314 16270
rect 1934 16210 1986 16222
rect 27358 16210 27410 16222
rect 24770 16158 24782 16210
rect 24834 16158 24846 16210
rect 26898 16158 26910 16210
rect 26962 16158 26974 16210
rect 1934 16146 1986 16158
rect 27358 16146 27410 16158
rect 16382 16098 16434 16110
rect 19966 16098 20018 16110
rect 4274 16046 4286 16098
rect 4338 16046 4350 16098
rect 16594 16046 16606 16098
rect 16658 16046 16670 16098
rect 16382 16034 16434 16046
rect 19966 16034 20018 16046
rect 21646 16098 21698 16110
rect 21646 16034 21698 16046
rect 21982 16098 22034 16110
rect 23986 16046 23998 16098
rect 24050 16046 24062 16098
rect 21982 16034 22034 16046
rect 15374 15986 15426 15998
rect 21758 15986 21810 15998
rect 19618 15934 19630 15986
rect 19682 15934 19694 15986
rect 15374 15922 15426 15934
rect 21758 15922 21810 15934
rect 14814 15874 14866 15886
rect 14814 15810 14866 15822
rect 15262 15874 15314 15886
rect 15262 15810 15314 15822
rect 16494 15874 16546 15886
rect 16494 15810 16546 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 15486 15538 15538 15550
rect 15486 15474 15538 15486
rect 16718 15538 16770 15550
rect 16718 15474 16770 15486
rect 17390 15538 17442 15550
rect 17390 15474 17442 15486
rect 15150 15426 15202 15438
rect 13794 15374 13806 15426
rect 13858 15374 13870 15426
rect 15150 15362 15202 15374
rect 16606 15426 16658 15438
rect 17714 15374 17726 15426
rect 17778 15374 17790 15426
rect 16606 15362 16658 15374
rect 15262 15314 15314 15326
rect 14578 15262 14590 15314
rect 14642 15262 14654 15314
rect 15262 15250 15314 15262
rect 15598 15314 15650 15326
rect 15598 15250 15650 15262
rect 16942 15314 16994 15326
rect 16942 15250 16994 15262
rect 11666 15150 11678 15202
rect 11730 15150 11742 15202
rect 15138 15150 15150 15202
rect 15202 15150 15214 15202
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 14926 14754 14978 14766
rect 14926 14690 14978 14702
rect 18398 14754 18450 14766
rect 18398 14690 18450 14702
rect 19182 14754 19234 14766
rect 19182 14690 19234 14702
rect 19630 14754 19682 14766
rect 19630 14690 19682 14702
rect 19742 14754 19794 14766
rect 19742 14690 19794 14702
rect 21534 14754 21586 14766
rect 21534 14690 21586 14702
rect 21758 14754 21810 14766
rect 21758 14690 21810 14702
rect 23998 14754 24050 14766
rect 23998 14690 24050 14702
rect 24334 14754 24386 14766
rect 24334 14690 24386 14702
rect 17054 14642 17106 14654
rect 17054 14578 17106 14590
rect 21422 14642 21474 14654
rect 21422 14578 21474 14590
rect 17166 14530 17218 14542
rect 16818 14478 16830 14530
rect 16882 14478 16894 14530
rect 17166 14466 17218 14478
rect 17726 14530 17778 14542
rect 18622 14530 18674 14542
rect 18274 14478 18286 14530
rect 18338 14478 18350 14530
rect 17726 14466 17778 14478
rect 18622 14466 18674 14478
rect 18958 14530 19010 14542
rect 18958 14466 19010 14478
rect 19518 14530 19570 14542
rect 19518 14466 19570 14478
rect 20414 14530 20466 14542
rect 20414 14466 20466 14478
rect 14702 14418 14754 14430
rect 14702 14354 14754 14366
rect 21870 14418 21922 14430
rect 21870 14354 21922 14366
rect 14814 14306 14866 14318
rect 14814 14242 14866 14254
rect 17390 14306 17442 14318
rect 17390 14242 17442 14254
rect 17614 14306 17666 14318
rect 17614 14242 17666 14254
rect 18062 14306 18114 14318
rect 18062 14242 18114 14254
rect 20750 14306 20802 14318
rect 20750 14242 20802 14254
rect 24110 14306 24162 14318
rect 24110 14242 24162 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 25342 13970 25394 13982
rect 25342 13906 25394 13918
rect 16270 13858 16322 13870
rect 13122 13806 13134 13858
rect 13186 13806 13198 13858
rect 16270 13794 16322 13806
rect 16830 13858 16882 13870
rect 19618 13806 19630 13858
rect 19682 13806 19694 13858
rect 22418 13806 22430 13858
rect 22482 13806 22494 13858
rect 16830 13794 16882 13806
rect 16494 13746 16546 13758
rect 12450 13694 12462 13746
rect 12514 13694 12526 13746
rect 20402 13694 20414 13746
rect 20466 13694 20478 13746
rect 21746 13694 21758 13746
rect 21810 13694 21822 13746
rect 16494 13682 16546 13694
rect 15710 13634 15762 13646
rect 15250 13582 15262 13634
rect 15314 13582 15326 13634
rect 15710 13570 15762 13582
rect 16382 13634 16434 13646
rect 20862 13634 20914 13646
rect 17490 13582 17502 13634
rect 17554 13582 17566 13634
rect 24546 13582 24558 13634
rect 24610 13582 24622 13634
rect 16382 13570 16434 13582
rect 20862 13570 20914 13582
rect 15474 13470 15486 13522
rect 15538 13519 15550 13522
rect 16034 13519 16046 13522
rect 15538 13473 16046 13519
rect 15538 13470 15550 13473
rect 16034 13470 16046 13473
rect 16098 13470 16110 13522
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 18062 13074 18114 13086
rect 15362 13022 15374 13074
rect 15426 13022 15438 13074
rect 17490 13022 17502 13074
rect 17554 13022 17566 13074
rect 18062 13010 18114 13022
rect 14690 12910 14702 12962
rect 14754 12910 14766 12962
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 23550 12402 23602 12414
rect 23550 12338 23602 12350
rect 20962 12238 20974 12290
rect 21026 12238 21038 12290
rect 20290 12126 20302 12178
rect 20354 12126 20366 12178
rect 23090 12014 23102 12066
rect 23154 12014 23166 12066
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 16718 5234 16770 5246
rect 16718 5170 16770 5182
rect 15698 5070 15710 5122
rect 15762 5070 15774 5122
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 19730 4286 19742 4338
rect 19794 4286 19806 4338
rect 20750 4114 20802 4126
rect 20750 4050 20802 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 18622 3666 18674 3678
rect 18622 3602 18674 3614
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 17602 3502 17614 3554
rect 17666 3502 17678 3554
rect 23538 3502 23550 3554
rect 23602 3502 23614 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 22194 3390 22206 3442
rect 22258 3390 22270 3442
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 18062 38222 18114 38274
rect 22430 38222 22482 38274
rect 25566 38222 25618 38274
rect 17054 37998 17106 38050
rect 21758 37998 21810 38050
rect 24558 37998 24610 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 19854 37438 19906 37490
rect 22766 37438 22818 37490
rect 26798 37438 26850 37490
rect 18846 37214 18898 37266
rect 22094 37214 22146 37266
rect 25790 37214 25842 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 19182 29374 19234 29426
rect 19854 29262 19906 29314
rect 21982 29262 22034 29314
rect 22542 29262 22594 29314
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 15150 28590 15202 28642
rect 18510 28590 18562 28642
rect 21982 28590 22034 28642
rect 15262 28478 15314 28530
rect 18734 28478 18786 28530
rect 18846 28478 18898 28530
rect 21758 28478 21810 28530
rect 17166 28366 17218 28418
rect 17614 28366 17666 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 14366 27918 14418 27970
rect 13694 27806 13746 27858
rect 17390 27806 17442 27858
rect 21646 27806 21698 27858
rect 25342 27806 25394 27858
rect 16494 27694 16546 27746
rect 18174 27694 18226 27746
rect 20302 27694 20354 27746
rect 22430 27694 22482 27746
rect 24558 27694 24610 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 15486 27246 15538 27298
rect 19966 27246 20018 27298
rect 15822 27134 15874 27186
rect 16494 27134 16546 27186
rect 17390 27134 17442 27186
rect 19630 27134 19682 27186
rect 22094 27134 22146 27186
rect 25678 27134 25730 27186
rect 26126 27134 26178 27186
rect 40014 27134 40066 27186
rect 16606 27022 16658 27074
rect 17054 27022 17106 27074
rect 17502 27022 17554 27074
rect 18398 27022 18450 27074
rect 18734 27022 18786 27074
rect 18846 27022 18898 27074
rect 19182 27022 19234 27074
rect 19518 27022 19570 27074
rect 20302 27022 20354 27074
rect 22766 27022 22818 27074
rect 37662 27022 37714 27074
rect 16046 26910 16098 26962
rect 16382 26910 16434 26962
rect 18062 26910 18114 26962
rect 19742 26910 19794 26962
rect 21982 26910 22034 26962
rect 22206 26910 22258 26962
rect 22430 26910 22482 26962
rect 23550 26910 23602 26962
rect 18510 26798 18562 26850
rect 21870 26798 21922 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 18174 26462 18226 26514
rect 21422 26462 21474 26514
rect 23550 26462 23602 26514
rect 24446 26462 24498 26514
rect 4286 26238 4338 26290
rect 14590 26238 14642 26290
rect 18846 26238 18898 26290
rect 19070 26238 19122 26290
rect 19294 26238 19346 26290
rect 23438 26238 23490 26290
rect 23662 26238 23714 26290
rect 23998 26238 24050 26290
rect 24334 26238 24386 26290
rect 25566 26238 25618 26290
rect 11790 26126 11842 26178
rect 13918 26126 13970 26178
rect 15150 26126 15202 26178
rect 18062 26126 18114 26178
rect 21310 26126 21362 26178
rect 26350 26126 26402 26178
rect 28478 26126 28530 26178
rect 28926 26126 28978 26178
rect 1934 26014 1986 26066
rect 17950 26014 18002 26066
rect 19406 26014 19458 26066
rect 21646 26014 21698 26066
rect 24446 26014 24498 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 15822 25678 15874 25730
rect 24446 25566 24498 25618
rect 25790 25566 25842 25618
rect 40014 25566 40066 25618
rect 14814 25454 14866 25506
rect 15262 25454 15314 25506
rect 15486 25454 15538 25506
rect 15710 25454 15762 25506
rect 18286 25454 18338 25506
rect 21310 25454 21362 25506
rect 24670 25454 24722 25506
rect 25902 25454 25954 25506
rect 37662 25454 37714 25506
rect 14702 25342 14754 25394
rect 14926 25342 14978 25394
rect 17502 25342 17554 25394
rect 17838 25342 17890 25394
rect 18510 25342 18562 25394
rect 24334 25342 24386 25394
rect 24894 25342 24946 25394
rect 26126 25342 26178 25394
rect 27246 25342 27298 25394
rect 27470 25342 27522 25394
rect 27582 25342 27634 25394
rect 21422 25230 21474 25282
rect 21646 25230 21698 25282
rect 25566 25230 25618 25282
rect 25678 25230 25730 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 16494 24894 16546 24946
rect 18286 24894 18338 24946
rect 26462 24894 26514 24946
rect 18622 24782 18674 24834
rect 23998 24782 24050 24834
rect 26910 24782 26962 24834
rect 30942 24782 30994 24834
rect 16718 24670 16770 24722
rect 17390 24670 17442 24722
rect 17838 24670 17890 24722
rect 24334 24670 24386 24722
rect 24558 24670 24610 24722
rect 27022 24670 27074 24722
rect 27358 24670 27410 24722
rect 30718 24670 30770 24722
rect 37662 24670 37714 24722
rect 24110 24558 24162 24610
rect 28142 24558 28194 24610
rect 30270 24558 30322 24610
rect 17614 24446 17666 24498
rect 17950 24446 18002 24498
rect 26910 24446 26962 24498
rect 40014 24446 40066 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 28030 24110 28082 24162
rect 16942 23998 16994 24050
rect 25678 23998 25730 24050
rect 26126 23998 26178 24050
rect 26686 23998 26738 24050
rect 29262 23998 29314 24050
rect 40014 23998 40066 24050
rect 16158 23886 16210 23938
rect 16606 23886 16658 23938
rect 21982 23886 22034 23938
rect 22766 23886 22818 23938
rect 28142 23886 28194 23938
rect 29038 23886 29090 23938
rect 37662 23886 37714 23938
rect 17278 23774 17330 23826
rect 21310 23774 21362 23826
rect 23550 23774 23602 23826
rect 28030 23774 28082 23826
rect 29598 23774 29650 23826
rect 17614 23662 17666 23714
rect 21422 23662 21474 23714
rect 21534 23662 21586 23714
rect 29374 23662 29426 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 16494 23326 16546 23378
rect 21086 23326 21138 23378
rect 21982 23326 22034 23378
rect 23662 23326 23714 23378
rect 23886 23326 23938 23378
rect 23998 23326 24050 23378
rect 24110 23326 24162 23378
rect 26462 23326 26514 23378
rect 12574 23214 12626 23266
rect 15934 23214 15986 23266
rect 17390 23214 17442 23266
rect 17726 23214 17778 23266
rect 19742 23214 19794 23266
rect 20414 23214 20466 23266
rect 21646 23214 21698 23266
rect 22094 23214 22146 23266
rect 27806 23214 27858 23266
rect 11902 23102 11954 23154
rect 15598 23102 15650 23154
rect 16046 23102 16098 23154
rect 16830 23102 16882 23154
rect 18062 23102 18114 23154
rect 19406 23102 19458 23154
rect 20078 23102 20130 23154
rect 21870 23102 21922 23154
rect 26126 23102 26178 23154
rect 27022 23102 27074 23154
rect 37662 23102 37714 23154
rect 14702 22990 14754 23042
rect 15150 22990 15202 23042
rect 15710 22990 15762 23042
rect 18398 22990 18450 23042
rect 21198 22990 21250 23042
rect 29934 22990 29986 23042
rect 18622 22878 18674 22930
rect 18958 22878 19010 22930
rect 20862 22878 20914 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 18286 22542 18338 22594
rect 19966 22542 20018 22594
rect 28254 22542 28306 22594
rect 16158 22430 16210 22482
rect 24894 22430 24946 22482
rect 40014 22430 40066 22482
rect 14814 22318 14866 22370
rect 16382 22318 16434 22370
rect 17726 22318 17778 22370
rect 19630 22318 19682 22370
rect 20414 22318 20466 22370
rect 21534 22318 21586 22370
rect 23886 22318 23938 22370
rect 24222 22318 24274 22370
rect 25230 22318 25282 22370
rect 28366 22318 28418 22370
rect 37886 22318 37938 22370
rect 16046 22206 16098 22258
rect 17054 22206 17106 22258
rect 17502 22206 17554 22258
rect 21310 22206 21362 22258
rect 22206 22206 22258 22258
rect 23214 22206 23266 22258
rect 26686 22206 26738 22258
rect 27022 22206 27074 22258
rect 28142 22206 28194 22258
rect 28590 22206 28642 22258
rect 15038 22094 15090 22146
rect 15374 22094 15426 22146
rect 15710 22094 15762 22146
rect 16718 22094 16770 22146
rect 18622 22094 18674 22146
rect 19294 22094 19346 22146
rect 19406 22094 19458 22146
rect 19518 22094 19570 22146
rect 20750 22094 20802 22146
rect 21870 22094 21922 22146
rect 22542 22094 22594 22146
rect 22878 22094 22930 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 16382 21758 16434 21810
rect 17390 21758 17442 21810
rect 17950 21758 18002 21810
rect 25342 21758 25394 21810
rect 25454 21758 25506 21810
rect 26910 21758 26962 21810
rect 12574 21646 12626 21698
rect 15934 21646 15986 21698
rect 16718 21646 16770 21698
rect 16830 21646 16882 21698
rect 17502 21646 17554 21698
rect 11902 21534 11954 21586
rect 15710 21534 15762 21586
rect 15822 21534 15874 21586
rect 17838 21534 17890 21586
rect 18174 21534 18226 21586
rect 18622 21534 18674 21586
rect 18958 21534 19010 21586
rect 27246 21534 27298 21586
rect 37662 21534 37714 21586
rect 14702 21422 14754 21474
rect 15150 21422 15202 21474
rect 22654 21422 22706 21474
rect 28030 21422 28082 21474
rect 30158 21422 30210 21474
rect 37438 21422 37490 21474
rect 39902 21422 39954 21474
rect 25230 21310 25282 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 1934 20862 1986 20914
rect 9998 20862 10050 20914
rect 13582 20862 13634 20914
rect 15374 20862 15426 20914
rect 22318 20862 22370 20914
rect 29262 20862 29314 20914
rect 40014 20862 40066 20914
rect 4286 20750 4338 20802
rect 12910 20750 12962 20802
rect 20078 20750 20130 20802
rect 21982 20750 22034 20802
rect 22654 20750 22706 20802
rect 28142 20750 28194 20802
rect 28478 20750 28530 20802
rect 29038 20750 29090 20802
rect 29374 20750 29426 20802
rect 37886 20750 37938 20802
rect 12126 20638 12178 20690
rect 21758 20638 21810 20690
rect 22094 20638 22146 20690
rect 26798 20638 26850 20690
rect 29598 20638 29650 20690
rect 21534 20526 21586 20578
rect 28366 20526 28418 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 11902 20190 11954 20242
rect 17614 20190 17666 20242
rect 22878 20190 22930 20242
rect 15822 20078 15874 20130
rect 17726 20078 17778 20130
rect 19518 20078 19570 20130
rect 20974 20078 21026 20130
rect 21534 20078 21586 20130
rect 22206 20078 22258 20130
rect 23438 20078 23490 20130
rect 27134 20078 27186 20130
rect 28366 20078 28418 20130
rect 28478 20078 28530 20130
rect 29710 20078 29762 20130
rect 12238 19966 12290 20018
rect 17390 19966 17442 20018
rect 20078 19966 20130 20018
rect 20302 19966 20354 20018
rect 20414 19966 20466 20018
rect 22766 19966 22818 20018
rect 23102 19966 23154 20018
rect 27358 19966 27410 20018
rect 27806 19966 27858 20018
rect 28142 19966 28194 20018
rect 29374 19966 29426 20018
rect 37662 19966 37714 20018
rect 21422 19854 21474 19906
rect 22094 19854 22146 19906
rect 22430 19854 22482 19906
rect 27582 19854 27634 19906
rect 15710 19742 15762 19794
rect 16046 19742 16098 19794
rect 21758 19742 21810 19794
rect 40014 19742 40066 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 14702 19406 14754 19458
rect 15822 19406 15874 19458
rect 15598 19294 15650 19346
rect 16158 19294 16210 19346
rect 16606 19294 16658 19346
rect 19630 19294 19682 19346
rect 22430 19294 22482 19346
rect 23998 19294 24050 19346
rect 26126 19294 26178 19346
rect 40014 19294 40066 19346
rect 14142 19182 14194 19234
rect 14366 19182 14418 19234
rect 17278 19182 17330 19234
rect 18622 19182 18674 19234
rect 19294 19182 19346 19234
rect 20190 19182 20242 19234
rect 22318 19182 22370 19234
rect 22542 19182 22594 19234
rect 22766 19182 22818 19234
rect 23326 19182 23378 19234
rect 27918 19182 27970 19234
rect 37662 19182 37714 19234
rect 19070 19070 19122 19122
rect 16494 18958 16546 19010
rect 16942 18958 16994 19010
rect 18510 18958 18562 19010
rect 26574 18958 26626 19010
rect 28142 18958 28194 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 14590 18622 14642 18674
rect 14926 18622 14978 18674
rect 15822 18622 15874 18674
rect 16046 18622 16098 18674
rect 22094 18622 22146 18674
rect 23550 18622 23602 18674
rect 25230 18622 25282 18674
rect 25454 18622 25506 18674
rect 11678 18510 11730 18562
rect 19182 18510 19234 18562
rect 19630 18510 19682 18562
rect 21198 18510 21250 18562
rect 21870 18510 21922 18562
rect 23102 18510 23154 18562
rect 23326 18510 23378 18562
rect 27806 18510 27858 18562
rect 11006 18398 11058 18450
rect 15598 18398 15650 18450
rect 16270 18398 16322 18450
rect 17950 18398 18002 18450
rect 18510 18398 18562 18450
rect 18958 18398 19010 18450
rect 19518 18398 19570 18450
rect 20638 18398 20690 18450
rect 21534 18398 21586 18450
rect 22878 18398 22930 18450
rect 25902 18398 25954 18450
rect 27022 18398 27074 18450
rect 37662 18398 37714 18450
rect 13806 18286 13858 18338
rect 14254 18286 14306 18338
rect 15934 18286 15986 18338
rect 17502 18286 17554 18338
rect 20302 18286 20354 18338
rect 25342 18286 25394 18338
rect 26686 18286 26738 18338
rect 29934 18286 29986 18338
rect 18398 18174 18450 18226
rect 22206 18174 22258 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 18062 17838 18114 17890
rect 22878 17838 22930 17890
rect 10782 17726 10834 17778
rect 12910 17726 12962 17778
rect 17054 17726 17106 17778
rect 21870 17726 21922 17778
rect 22654 17726 22706 17778
rect 28254 17726 28306 17778
rect 40014 17726 40066 17778
rect 10110 17614 10162 17666
rect 14478 17614 14530 17666
rect 16270 17614 16322 17666
rect 17166 17614 17218 17666
rect 18286 17614 18338 17666
rect 18510 17614 18562 17666
rect 19518 17614 19570 17666
rect 20862 17614 20914 17666
rect 21534 17614 21586 17666
rect 22094 17614 22146 17666
rect 23774 17614 23826 17666
rect 23886 17614 23938 17666
rect 23998 17614 24050 17666
rect 24334 17614 24386 17666
rect 25342 17614 25394 17666
rect 37662 17614 37714 17666
rect 14814 17502 14866 17554
rect 16494 17502 16546 17554
rect 18622 17502 18674 17554
rect 19406 17502 19458 17554
rect 20078 17502 20130 17554
rect 20526 17502 20578 17554
rect 21646 17502 21698 17554
rect 24222 17502 24274 17554
rect 26126 17502 26178 17554
rect 13582 17390 13634 17442
rect 15486 17390 15538 17442
rect 15822 17390 15874 17442
rect 20638 17390 20690 17442
rect 21870 17390 21922 17442
rect 23214 17390 23266 17442
rect 29262 17390 29314 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 19294 17054 19346 17106
rect 19630 17054 19682 17106
rect 20190 17054 20242 17106
rect 21198 17054 21250 17106
rect 21758 17054 21810 17106
rect 21982 17054 22034 17106
rect 22094 17054 22146 17106
rect 22990 17054 23042 17106
rect 15486 16942 15538 16994
rect 15710 16942 15762 16994
rect 15934 16942 15986 16994
rect 19966 16942 20018 16994
rect 22766 16942 22818 16994
rect 24110 16942 24162 16994
rect 24334 16942 24386 16994
rect 15262 16830 15314 16882
rect 20638 16830 20690 16882
rect 20862 16830 20914 16882
rect 21534 16830 21586 16882
rect 22542 16830 22594 16882
rect 23102 16830 23154 16882
rect 23550 16830 23602 16882
rect 20302 16718 20354 16770
rect 22878 16718 22930 16770
rect 24222 16718 24274 16770
rect 23774 16606 23826 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 15262 16270 15314 16322
rect 1934 16158 1986 16210
rect 24782 16158 24834 16210
rect 26910 16158 26962 16210
rect 27358 16158 27410 16210
rect 4286 16046 4338 16098
rect 16382 16046 16434 16098
rect 16606 16046 16658 16098
rect 19966 16046 20018 16098
rect 21646 16046 21698 16098
rect 21982 16046 22034 16098
rect 23998 16046 24050 16098
rect 15374 15934 15426 15986
rect 19630 15934 19682 15986
rect 21758 15934 21810 15986
rect 14814 15822 14866 15874
rect 15262 15822 15314 15874
rect 16494 15822 16546 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 15486 15486 15538 15538
rect 16718 15486 16770 15538
rect 17390 15486 17442 15538
rect 13806 15374 13858 15426
rect 15150 15374 15202 15426
rect 16606 15374 16658 15426
rect 17726 15374 17778 15426
rect 14590 15262 14642 15314
rect 15262 15262 15314 15314
rect 15598 15262 15650 15314
rect 16942 15262 16994 15314
rect 11678 15150 11730 15202
rect 15150 15150 15202 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 14926 14702 14978 14754
rect 18398 14702 18450 14754
rect 19182 14702 19234 14754
rect 19630 14702 19682 14754
rect 19742 14702 19794 14754
rect 21534 14702 21586 14754
rect 21758 14702 21810 14754
rect 23998 14702 24050 14754
rect 24334 14702 24386 14754
rect 17054 14590 17106 14642
rect 21422 14590 21474 14642
rect 16830 14478 16882 14530
rect 17166 14478 17218 14530
rect 17726 14478 17778 14530
rect 18286 14478 18338 14530
rect 18622 14478 18674 14530
rect 18958 14478 19010 14530
rect 19518 14478 19570 14530
rect 20414 14478 20466 14530
rect 14702 14366 14754 14418
rect 21870 14366 21922 14418
rect 14814 14254 14866 14306
rect 17390 14254 17442 14306
rect 17614 14254 17666 14306
rect 18062 14254 18114 14306
rect 20750 14254 20802 14306
rect 24110 14254 24162 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 25342 13918 25394 13970
rect 13134 13806 13186 13858
rect 16270 13806 16322 13858
rect 16830 13806 16882 13858
rect 19630 13806 19682 13858
rect 22430 13806 22482 13858
rect 12462 13694 12514 13746
rect 16494 13694 16546 13746
rect 20414 13694 20466 13746
rect 21758 13694 21810 13746
rect 15262 13582 15314 13634
rect 15710 13582 15762 13634
rect 16382 13582 16434 13634
rect 17502 13582 17554 13634
rect 20862 13582 20914 13634
rect 24558 13582 24610 13634
rect 15486 13470 15538 13522
rect 16046 13470 16098 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 15374 13022 15426 13074
rect 17502 13022 17554 13074
rect 18062 13022 18114 13074
rect 14702 12910 14754 12962
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 23550 12350 23602 12402
rect 20974 12238 21026 12290
rect 20302 12126 20354 12178
rect 23102 12014 23154 12066
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 16718 5182 16770 5234
rect 15710 5070 15762 5122
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 19742 4286 19794 4338
rect 20750 4062 20802 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18622 3614 18674 3666
rect 25566 3614 25618 3666
rect 17614 3502 17666 3554
rect 23550 3502 23602 3554
rect 24558 3502 24610 3554
rect 22206 3390 22258 3442
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 16800 41200 16912 42000
rect 18816 41200 18928 42000
rect 21504 41200 21616 42000
rect 22176 41200 22288 42000
rect 24192 41200 24304 42000
rect 25536 41200 25648 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 16828 38276 16884 41200
rect 16828 38210 16884 38220
rect 18060 38276 18116 38286
rect 18060 38182 18116 38220
rect 17052 38050 17108 38062
rect 17052 37998 17054 38050
rect 17106 37998 17108 38050
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 17052 31948 17108 37998
rect 18844 37492 18900 41200
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 18844 37426 18900 37436
rect 19852 37492 19908 37502
rect 19852 37398 19908 37436
rect 21532 37492 21588 41200
rect 22204 38276 22260 41200
rect 22428 38276 22484 38286
rect 22204 38274 22484 38276
rect 22204 38222 22430 38274
rect 22482 38222 22484 38274
rect 22204 38220 22484 38222
rect 22428 38210 22484 38220
rect 24220 38276 24276 41200
rect 25564 38612 25620 41200
rect 25564 38546 25620 38556
rect 26796 38612 26852 38622
rect 24220 38210 24276 38220
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 21532 37426 21588 37436
rect 21756 38050 21812 38062
rect 21756 37998 21758 38050
rect 21810 37998 21812 38050
rect 18844 37266 18900 37278
rect 18844 37214 18846 37266
rect 18898 37214 18900 37266
rect 18844 31948 18900 37214
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 16828 31892 17108 31948
rect 18732 31892 18900 31948
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 14364 28644 14420 28654
rect 14364 27970 14420 28588
rect 15148 28644 15204 28654
rect 15148 28550 15204 28588
rect 15260 28532 15316 28542
rect 16828 28532 16884 31892
rect 18508 28644 18564 28654
rect 15260 28530 15540 28532
rect 15260 28478 15262 28530
rect 15314 28478 15540 28530
rect 15260 28476 15540 28478
rect 15260 28466 15316 28476
rect 14364 27918 14366 27970
rect 14418 27918 14420 27970
rect 14364 27906 14420 27918
rect 13692 27858 13748 27870
rect 13692 27806 13694 27858
rect 13746 27806 13748 27858
rect 4172 27636 4228 27646
rect 1932 26066 1988 26078
rect 1932 26014 1934 26066
rect 1986 26014 1988 26066
rect 1932 25620 1988 26014
rect 1932 25554 1988 25564
rect 4172 21476 4228 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 13692 26516 13748 27806
rect 15484 27298 15540 28476
rect 16492 28476 16884 28532
rect 18396 28642 18564 28644
rect 18396 28590 18510 28642
rect 18562 28590 18564 28642
rect 18396 28588 18564 28590
rect 16492 27748 16548 28476
rect 17164 28420 17220 28430
rect 17612 28420 17668 28430
rect 17164 28418 17668 28420
rect 17164 28366 17166 28418
rect 17218 28366 17614 28418
rect 17666 28366 17668 28418
rect 17164 28364 17668 28366
rect 17164 28354 17220 28364
rect 17388 27860 17444 28364
rect 17612 28354 17668 28364
rect 17276 27858 17444 27860
rect 17276 27806 17390 27858
rect 17442 27806 17444 27858
rect 17276 27804 17444 27806
rect 16492 27746 16660 27748
rect 16492 27694 16494 27746
rect 16546 27694 16660 27746
rect 16492 27692 16660 27694
rect 16492 27682 16548 27692
rect 15484 27246 15486 27298
rect 15538 27246 15540 27298
rect 15484 27234 15540 27246
rect 15820 27188 15876 27198
rect 16492 27188 16548 27198
rect 15820 27186 16548 27188
rect 15820 27134 15822 27186
rect 15874 27134 16494 27186
rect 16546 27134 16548 27186
rect 15820 27132 16548 27134
rect 15820 27122 15876 27132
rect 16492 27122 16548 27132
rect 16604 27074 16660 27692
rect 16604 27022 16606 27074
rect 16658 27022 16660 27074
rect 16604 27010 16660 27022
rect 17052 27074 17108 27086
rect 17052 27022 17054 27074
rect 17106 27022 17108 27074
rect 16044 26962 16100 26974
rect 16044 26910 16046 26962
rect 16098 26910 16100 26962
rect 13692 26450 13748 26460
rect 14588 26516 14644 26526
rect 4284 26292 4340 26302
rect 4284 26198 4340 26236
rect 11788 26292 11844 26302
rect 11788 26178 11844 26236
rect 14588 26290 14644 26460
rect 15148 26516 15204 26526
rect 14588 26238 14590 26290
rect 14642 26238 14644 26290
rect 14588 26226 14644 26238
rect 14700 26292 14756 26302
rect 11788 26126 11790 26178
rect 11842 26126 11844 26178
rect 11788 26114 11844 26126
rect 13916 26178 13972 26190
rect 13916 26126 13918 26178
rect 13970 26126 13972 26178
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 13916 25732 13972 26126
rect 13916 25666 13972 25676
rect 14700 25394 14756 26236
rect 15148 26178 15204 26460
rect 15148 26126 15150 26178
rect 15202 26126 15204 26178
rect 14812 25508 14868 25518
rect 14812 25414 14868 25452
rect 14700 25342 14702 25394
rect 14754 25342 14756 25394
rect 14700 25330 14756 25342
rect 14924 25394 14980 25406
rect 14924 25342 14926 25394
rect 14978 25342 14980 25394
rect 12572 24500 12628 24510
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 12572 23266 12628 24444
rect 12572 23214 12574 23266
rect 12626 23214 12628 23266
rect 12572 23202 12628 23214
rect 14812 23940 14868 23950
rect 11900 23154 11956 23166
rect 11900 23102 11902 23154
rect 11954 23102 11956 23154
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4172 21410 4228 21420
rect 11900 21586 11956 23102
rect 12684 23044 12740 23054
rect 12572 21700 12628 21710
rect 12684 21700 12740 22988
rect 14700 23042 14756 23054
rect 14700 22990 14702 23042
rect 14754 22990 14756 23042
rect 14700 22596 14756 22990
rect 14700 22530 14756 22540
rect 14812 22370 14868 23884
rect 14924 23604 14980 25342
rect 14924 23538 14980 23548
rect 14812 22318 14814 22370
rect 14866 22318 14868 22370
rect 12572 21698 12740 21700
rect 12572 21646 12574 21698
rect 12626 21646 12740 21698
rect 12572 21644 12740 21646
rect 14700 21812 14756 21822
rect 12572 21634 12628 21644
rect 11900 21534 11902 21586
rect 11954 21534 11956 21586
rect 9996 21252 10052 21262
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 1932 20914 1988 20926
rect 1932 20862 1934 20914
rect 1986 20862 1988 20914
rect 1932 20244 1988 20862
rect 9996 20916 10052 21196
rect 9996 20822 10052 20860
rect 11900 20916 11956 21534
rect 14700 21474 14756 21756
rect 14700 21422 14702 21474
rect 14754 21422 14756 21474
rect 14700 21410 14756 21422
rect 11900 20850 11956 20860
rect 12908 20916 12964 20926
rect 4284 20804 4340 20814
rect 4284 20710 4340 20748
rect 12908 20802 12964 20860
rect 12908 20750 12910 20802
rect 12962 20750 12964 20802
rect 12908 20738 12964 20750
rect 13580 20916 13636 20926
rect 12124 20692 12180 20702
rect 1932 20178 1988 20188
rect 11900 20690 12180 20692
rect 11900 20638 12126 20690
rect 12178 20638 12180 20690
rect 11900 20636 12180 20638
rect 11900 20242 11956 20636
rect 12124 20626 12180 20636
rect 11900 20190 11902 20242
rect 11954 20190 11956 20242
rect 11900 20178 11956 20190
rect 12236 20020 12292 20030
rect 12236 19926 12292 19964
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 11676 18564 11732 18574
rect 11676 18470 11732 18508
rect 11004 18450 11060 18462
rect 11004 18398 11006 18450
rect 11058 18398 11060 18450
rect 10108 18340 10164 18350
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 10108 17666 10164 18284
rect 11004 18340 11060 18398
rect 11004 18274 11060 18284
rect 10780 18228 10836 18238
rect 10780 17778 10836 18172
rect 10780 17726 10782 17778
rect 10834 17726 10836 17778
rect 10780 17714 10836 17726
rect 12908 17780 12964 17790
rect 12908 17686 12964 17724
rect 10108 17614 10110 17666
rect 10162 17614 10164 17666
rect 10108 17602 10164 17614
rect 13580 17442 13636 20860
rect 14812 20188 14868 22318
rect 15148 23042 15204 26126
rect 15820 25732 15876 25742
rect 15820 25638 15876 25676
rect 15260 25508 15316 25518
rect 15260 25414 15316 25452
rect 15484 25506 15540 25518
rect 15484 25454 15486 25506
rect 15538 25454 15540 25506
rect 15484 25172 15540 25454
rect 15484 25106 15540 25116
rect 15708 25506 15764 25518
rect 15708 25454 15710 25506
rect 15762 25454 15764 25506
rect 15708 24948 15764 25454
rect 15708 24882 15764 24892
rect 15148 22990 15150 23042
rect 15202 22990 15204 23042
rect 15036 22148 15092 22158
rect 15036 22054 15092 22092
rect 15148 21474 15204 22990
rect 15484 23604 15540 23614
rect 15372 22146 15428 22158
rect 15372 22094 15374 22146
rect 15426 22094 15428 22146
rect 15372 21924 15428 22094
rect 15372 21858 15428 21868
rect 15148 21422 15150 21474
rect 15202 21422 15204 21474
rect 15148 20916 15204 21422
rect 15372 20916 15428 20926
rect 15204 20914 15428 20916
rect 15204 20862 15374 20914
rect 15426 20862 15428 20914
rect 15204 20860 15428 20862
rect 15148 20822 15204 20860
rect 15372 20850 15428 20860
rect 14700 20132 14868 20188
rect 14700 19460 14756 20132
rect 13804 19404 14308 19460
rect 13804 18338 13860 19404
rect 14140 19234 14196 19246
rect 14140 19182 14142 19234
rect 14194 19182 14196 19234
rect 14140 18564 14196 19182
rect 14252 19236 14308 19404
rect 14700 19366 14756 19404
rect 14924 19572 14980 19582
rect 14364 19236 14420 19246
rect 14252 19234 14644 19236
rect 14252 19182 14366 19234
rect 14418 19182 14644 19234
rect 14252 19180 14644 19182
rect 14364 19170 14420 19180
rect 14588 18674 14644 19180
rect 14588 18622 14590 18674
rect 14642 18622 14644 18674
rect 14588 18610 14644 18622
rect 14924 18674 14980 19516
rect 15484 19460 15540 23548
rect 15932 23268 15988 23278
rect 15932 23174 15988 23212
rect 15596 23154 15652 23166
rect 15596 23102 15598 23154
rect 15650 23102 15652 23154
rect 15596 22260 15652 23102
rect 16044 23154 16100 26910
rect 16380 26964 16436 26974
rect 16380 26870 16436 26908
rect 17052 26404 17108 27022
rect 17276 26516 17332 27804
rect 17388 27794 17444 27804
rect 18172 27746 18228 27758
rect 18172 27694 18174 27746
rect 18226 27694 18228 27746
rect 17276 26450 17332 26460
rect 17388 27186 17444 27198
rect 17388 27134 17390 27186
rect 17442 27134 17444 27186
rect 17052 26338 17108 26348
rect 17388 25172 17444 27134
rect 17500 27074 17556 27086
rect 17500 27022 17502 27074
rect 17554 27022 17556 27074
rect 17500 26964 17556 27022
rect 17500 26516 17556 26908
rect 17500 26450 17556 26460
rect 17948 27076 18004 27086
rect 17836 26404 17892 26414
rect 17836 26068 17892 26348
rect 17948 26292 18004 27020
rect 18060 26964 18116 26974
rect 18060 26870 18116 26908
rect 18172 26908 18228 27694
rect 18396 27074 18452 28588
rect 18508 28578 18564 28588
rect 18732 28530 18788 31892
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19180 29426 19236 29438
rect 19180 29374 19182 29426
rect 19234 29374 19236 29426
rect 18732 28478 18734 28530
rect 18786 28478 18788 28530
rect 18732 27748 18788 28478
rect 18844 28532 18900 28542
rect 19180 28532 19236 29374
rect 19852 29316 19908 29326
rect 18844 28530 19012 28532
rect 18844 28478 18846 28530
rect 18898 28478 19012 28530
rect 18844 28476 19012 28478
rect 18844 28466 18900 28476
rect 18732 27682 18788 27692
rect 18844 27300 18900 27310
rect 18396 27022 18398 27074
rect 18450 27022 18452 27074
rect 18396 27010 18452 27022
rect 18732 27074 18788 27086
rect 18732 27022 18734 27074
rect 18786 27022 18788 27074
rect 18732 26964 18788 27022
rect 18172 26852 18564 26908
rect 18732 26898 18788 26908
rect 18844 27074 18900 27244
rect 18844 27022 18846 27074
rect 18898 27022 18900 27074
rect 18508 26850 18564 26852
rect 18508 26798 18510 26850
rect 18562 26798 18564 26850
rect 18508 26786 18564 26798
rect 18844 26628 18900 27022
rect 18732 26572 18900 26628
rect 18172 26516 18228 26526
rect 18172 26422 18228 26460
rect 18508 26516 18564 26526
rect 17948 26236 18116 26292
rect 18060 26178 18116 26236
rect 18060 26126 18062 26178
rect 18114 26126 18116 26178
rect 17948 26068 18004 26078
rect 17500 26066 18004 26068
rect 17500 26014 17950 26066
rect 18002 26014 18004 26066
rect 17500 26012 18004 26014
rect 17500 25394 17556 26012
rect 17948 26002 18004 26012
rect 18060 25844 18116 26126
rect 17500 25342 17502 25394
rect 17554 25342 17556 25394
rect 17500 25330 17556 25342
rect 17724 25788 18116 25844
rect 17724 25172 17780 25788
rect 18284 25508 18340 25518
rect 18284 25506 18452 25508
rect 18284 25454 18286 25506
rect 18338 25454 18452 25506
rect 18284 25452 18452 25454
rect 18284 25442 18340 25452
rect 17836 25396 17892 25406
rect 17836 25394 18004 25396
rect 17836 25342 17838 25394
rect 17890 25342 18004 25394
rect 17836 25340 18004 25342
rect 17836 25330 17892 25340
rect 17724 25116 17892 25172
rect 16492 24948 16548 24958
rect 16492 24854 16548 24892
rect 16716 24724 16772 24734
rect 17388 24724 17444 25116
rect 16716 24630 16772 24668
rect 16940 24722 17444 24724
rect 16940 24670 17390 24722
rect 17442 24670 17444 24722
rect 16940 24668 17444 24670
rect 16940 24050 16996 24668
rect 17388 24658 17444 24668
rect 17724 24724 17780 24734
rect 16940 23998 16942 24050
rect 16994 23998 16996 24050
rect 16940 23986 16996 23998
rect 17612 24498 17668 24510
rect 17612 24446 17614 24498
rect 17666 24446 17668 24498
rect 16156 23940 16212 23950
rect 16156 23846 16212 23884
rect 16604 23938 16660 23950
rect 16604 23886 16606 23938
rect 16658 23886 16660 23938
rect 16604 23492 16660 23886
rect 17612 23940 17668 24446
rect 17612 23874 17668 23884
rect 17276 23828 17332 23838
rect 16492 23436 16604 23492
rect 16492 23378 16548 23436
rect 16604 23426 16660 23436
rect 16940 23826 17332 23828
rect 16940 23774 17278 23826
rect 17330 23774 17332 23826
rect 16940 23772 17332 23774
rect 16492 23326 16494 23378
rect 16546 23326 16548 23378
rect 16492 23314 16548 23326
rect 16044 23102 16046 23154
rect 16098 23102 16100 23154
rect 15708 23044 15764 23054
rect 15708 22950 15764 22988
rect 15596 22194 15652 22204
rect 15932 22596 15988 22606
rect 15708 22146 15764 22158
rect 15708 22094 15710 22146
rect 15762 22094 15764 22146
rect 15708 22036 15764 22094
rect 15708 21970 15764 21980
rect 15932 21924 15988 22540
rect 16044 22484 16100 23102
rect 16828 23156 16884 23166
rect 16828 23062 16884 23100
rect 16156 22484 16212 22494
rect 16044 22482 16212 22484
rect 16044 22430 16158 22482
rect 16210 22430 16212 22482
rect 16044 22428 16212 22430
rect 16156 22418 16212 22428
rect 16380 22484 16436 22494
rect 16380 22370 16436 22428
rect 16380 22318 16382 22370
rect 16434 22318 16436 22370
rect 16380 22306 16436 22318
rect 16044 22260 16100 22270
rect 16100 22204 16324 22260
rect 16044 22166 16100 22204
rect 15932 21698 15988 21868
rect 15932 21646 15934 21698
rect 15986 21646 15988 21698
rect 15932 21634 15988 21646
rect 15708 21586 15764 21598
rect 15708 21534 15710 21586
rect 15762 21534 15764 21586
rect 15708 20132 15764 21534
rect 15820 21586 15876 21598
rect 15820 21534 15822 21586
rect 15874 21534 15876 21586
rect 15820 20692 15876 21534
rect 16268 21588 16324 22204
rect 16380 22148 16436 22158
rect 16716 22148 16772 22158
rect 16940 22148 16996 23772
rect 17276 23762 17332 23772
rect 17612 23714 17668 23726
rect 17612 23662 17614 23714
rect 17666 23662 17668 23714
rect 17388 23268 17444 23278
rect 17388 23174 17444 23212
rect 17612 23156 17668 23662
rect 17612 22596 17668 23100
rect 17612 22530 17668 22540
rect 17724 23266 17780 24668
rect 17836 24722 17892 25116
rect 17948 25060 18004 25340
rect 17948 25004 18340 25060
rect 17836 24670 17838 24722
rect 17890 24670 17892 24722
rect 17836 24658 17892 24670
rect 17948 24500 18004 24510
rect 17948 24406 18004 24444
rect 18172 23492 18228 25004
rect 18284 24946 18340 25004
rect 18284 24894 18286 24946
rect 18338 24894 18340 24946
rect 18284 24882 18340 24894
rect 18396 24724 18452 25452
rect 18508 25394 18564 26460
rect 18508 25342 18510 25394
rect 18562 25342 18564 25394
rect 18508 25330 18564 25342
rect 18732 25060 18788 26572
rect 18844 26404 18900 26414
rect 18956 26404 19012 28476
rect 19180 28466 19236 28476
rect 19628 29314 19908 29316
rect 19628 29262 19854 29314
rect 19906 29262 19908 29314
rect 19628 29260 19908 29262
rect 19628 27186 19684 29260
rect 19852 29250 19908 29260
rect 21644 28532 21700 28542
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 21644 27858 21700 28476
rect 21756 28530 21812 37998
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 22764 37492 22820 37502
rect 22764 37398 22820 37436
rect 22092 37266 22148 37278
rect 22092 37214 22094 37266
rect 22146 37214 22148 37266
rect 21980 29316 22036 29326
rect 22092 29316 22148 37214
rect 21980 29314 22148 29316
rect 21980 29262 21982 29314
rect 22034 29262 22148 29314
rect 21980 29260 22148 29262
rect 22540 29314 22596 29326
rect 22540 29262 22542 29314
rect 22594 29262 22596 29314
rect 21980 28644 22036 29260
rect 21756 28478 21758 28530
rect 21810 28478 21812 28530
rect 21756 28466 21812 28478
rect 21868 28642 22036 28644
rect 21868 28590 21982 28642
rect 22034 28590 22036 28642
rect 21868 28588 22036 28590
rect 21644 27806 21646 27858
rect 21698 27806 21700 27858
rect 21644 27794 21700 27806
rect 20300 27748 20356 27758
rect 20300 27654 20356 27692
rect 19964 27300 20020 27310
rect 19964 27206 20020 27244
rect 19628 27134 19630 27186
rect 19682 27134 19684 27186
rect 19628 27122 19684 27134
rect 19180 27074 19236 27086
rect 19180 27022 19182 27074
rect 19234 27022 19236 27074
rect 18900 26348 19012 26404
rect 19068 26516 19124 26526
rect 18844 26290 18900 26348
rect 18844 26238 18846 26290
rect 18898 26238 18900 26290
rect 18844 26226 18900 26238
rect 19068 26290 19124 26460
rect 19068 26238 19070 26290
rect 19122 26238 19124 26290
rect 19068 26226 19124 26238
rect 19180 26068 19236 27022
rect 19516 27076 19572 27086
rect 19516 26982 19572 27020
rect 20300 27074 20356 27086
rect 21868 27076 21924 28588
rect 21980 28578 22036 28588
rect 22540 28532 22596 29262
rect 22596 28476 22820 28532
rect 22540 28466 22596 28476
rect 22428 27748 22484 27758
rect 22092 27746 22484 27748
rect 22092 27694 22430 27746
rect 22482 27694 22484 27746
rect 22092 27692 22484 27694
rect 22092 27186 22148 27692
rect 22428 27682 22484 27692
rect 22764 27748 22820 28476
rect 24556 27748 24612 37998
rect 26796 37490 26852 38556
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 26796 37438 26798 37490
rect 26850 37438 26852 37490
rect 26796 37426 26852 37438
rect 25788 37266 25844 37278
rect 25788 37214 25790 37266
rect 25842 37214 25844 37266
rect 25788 31948 25844 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 25676 31892 25844 31948
rect 25340 27858 25396 27870
rect 25340 27806 25342 27858
rect 25394 27806 25396 27858
rect 22092 27134 22094 27186
rect 22146 27134 22148 27186
rect 22092 27122 22148 27134
rect 20300 27022 20302 27074
rect 20354 27022 20356 27074
rect 19740 26962 19796 26974
rect 19740 26910 19742 26962
rect 19794 26910 19796 26962
rect 19740 26908 19796 26910
rect 19516 26852 19796 26908
rect 20300 26908 20356 27022
rect 21756 27020 21924 27076
rect 22764 27074 22820 27692
rect 22764 27022 22766 27074
rect 22818 27022 22820 27074
rect 21756 26908 21812 27020
rect 20300 26852 21364 26908
rect 19292 26292 19348 26302
rect 19516 26292 19572 26852
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19292 26290 19572 26292
rect 19292 26238 19294 26290
rect 19346 26238 19572 26290
rect 19292 26236 19572 26238
rect 19292 26226 19348 26236
rect 19404 26068 19460 26078
rect 19180 26066 19460 26068
rect 19180 26014 19406 26066
rect 19458 26014 19460 26066
rect 19180 26012 19460 26014
rect 19404 25508 19460 26012
rect 19404 25442 19460 25452
rect 18732 25004 19124 25060
rect 18620 24836 18676 24846
rect 18620 24742 18676 24780
rect 18844 24836 18900 24846
rect 18396 24658 18452 24668
rect 17724 23214 17726 23266
rect 17778 23214 17780 23266
rect 17052 22484 17108 22494
rect 17052 22258 17108 22428
rect 17724 22372 17780 23214
rect 17948 23268 18004 23278
rect 17948 22820 18004 23212
rect 18060 23156 18116 23166
rect 18172 23156 18228 23436
rect 18060 23154 18228 23156
rect 18060 23102 18062 23154
rect 18114 23102 18228 23154
rect 18060 23100 18228 23102
rect 18284 23828 18340 23838
rect 18060 23090 18116 23100
rect 17948 22764 18228 22820
rect 17612 22370 17780 22372
rect 17612 22318 17726 22370
rect 17778 22318 17780 22370
rect 17612 22316 17780 22318
rect 17500 22260 17556 22270
rect 17052 22206 17054 22258
rect 17106 22206 17108 22258
rect 17052 22194 17108 22206
rect 17164 22258 17556 22260
rect 17164 22206 17502 22258
rect 17554 22206 17556 22258
rect 17164 22204 17556 22206
rect 16380 21810 16436 22092
rect 16604 22146 16772 22148
rect 16604 22094 16718 22146
rect 16770 22094 16772 22146
rect 16604 22092 16772 22094
rect 16604 22036 16660 22092
rect 16716 22082 16772 22092
rect 16828 22092 16996 22148
rect 16604 21970 16660 21980
rect 16380 21758 16382 21810
rect 16434 21758 16436 21810
rect 16380 21746 16436 21758
rect 16716 21924 16772 21934
rect 16828 21924 16884 22092
rect 16772 21868 16884 21924
rect 16716 21698 16772 21868
rect 16716 21646 16718 21698
rect 16770 21646 16772 21698
rect 16716 21634 16772 21646
rect 16828 21700 16884 21710
rect 17164 21700 17220 22204
rect 17500 22194 17556 22204
rect 16828 21698 17220 21700
rect 16828 21646 16830 21698
rect 16882 21646 17220 21698
rect 16828 21644 17220 21646
rect 17276 22036 17332 22046
rect 17612 22036 17668 22316
rect 17724 22306 17780 22316
rect 18060 22596 18116 22606
rect 16828 21634 16884 21644
rect 15820 20636 15988 20692
rect 15820 20132 15876 20142
rect 15708 20130 15876 20132
rect 15708 20078 15822 20130
rect 15874 20078 15876 20130
rect 15708 20076 15876 20078
rect 14924 18622 14926 18674
rect 14978 18622 14980 18674
rect 14924 18610 14980 18622
rect 15372 19404 15540 19460
rect 15708 19794 15764 19806
rect 15708 19742 15710 19794
rect 15762 19742 15764 19794
rect 14140 18508 14532 18564
rect 13804 18286 13806 18338
rect 13858 18286 13860 18338
rect 13804 18274 13860 18286
rect 14252 18340 14308 18350
rect 13580 17390 13582 17442
rect 13634 17390 13636 17442
rect 13580 16884 13636 17390
rect 13580 16818 13636 16828
rect 13804 16996 13860 17006
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 1932 16210 1988 16222
rect 1932 16158 1934 16210
rect 1986 16158 1988 16210
rect 1932 15540 1988 16158
rect 1932 15474 1988 15484
rect 4284 16098 4340 16110
rect 4284 16046 4286 16098
rect 4338 16046 4340 16098
rect 4284 15316 4340 16046
rect 4284 15250 4340 15260
rect 11676 15876 11732 15886
rect 11676 15316 11732 15820
rect 13804 15426 13860 16940
rect 14252 16884 14308 18284
rect 14476 17780 14532 18508
rect 14476 17666 14532 17724
rect 14476 17614 14478 17666
rect 14530 17614 14532 17666
rect 14476 17602 14532 17614
rect 14812 18116 14868 18126
rect 14812 17554 14868 18060
rect 15372 17556 15428 19404
rect 15596 19348 15652 19358
rect 15708 19348 15764 19742
rect 15820 19684 15876 20076
rect 15932 19796 15988 20636
rect 16044 19796 16100 19806
rect 15932 19794 16100 19796
rect 15932 19742 16046 19794
rect 16098 19742 16100 19794
rect 15932 19740 16100 19742
rect 15820 19628 15988 19684
rect 15820 19460 15876 19470
rect 15820 19366 15876 19404
rect 15484 19346 15764 19348
rect 15484 19294 15598 19346
rect 15650 19294 15764 19346
rect 15484 19292 15764 19294
rect 15484 17668 15540 19292
rect 15596 19282 15652 19292
rect 15932 19236 15988 19628
rect 15708 19180 15988 19236
rect 16044 19572 16100 19740
rect 16044 19236 16100 19516
rect 16156 19348 16212 19358
rect 16156 19254 16212 19292
rect 15596 18450 15652 18462
rect 15596 18398 15598 18450
rect 15650 18398 15652 18450
rect 15596 17892 15652 18398
rect 15708 18116 15764 19180
rect 16044 19170 16100 19180
rect 15820 19012 15876 19022
rect 15820 18676 15876 18956
rect 15820 18582 15876 18620
rect 16044 18676 16100 18686
rect 16044 18582 16100 18620
rect 16268 18450 16324 21532
rect 16604 19348 16660 19358
rect 16604 19254 16660 19292
rect 16492 19012 16548 19022
rect 16492 18918 16548 18956
rect 16940 19010 16996 19022
rect 16940 18958 16942 19010
rect 16994 18958 16996 19010
rect 16940 18676 16996 18958
rect 16940 18610 16996 18620
rect 16268 18398 16270 18450
rect 16322 18398 16324 18450
rect 16268 18386 16324 18398
rect 15708 18050 15764 18060
rect 15932 18338 15988 18350
rect 15932 18286 15934 18338
rect 15986 18286 15988 18338
rect 15596 17826 15652 17836
rect 15932 17668 15988 18286
rect 16156 17780 16212 17790
rect 15484 17612 15652 17668
rect 14812 17502 14814 17554
rect 14866 17502 14868 17554
rect 14812 17490 14868 17502
rect 15148 17500 15540 17556
rect 14252 16818 14308 16828
rect 14812 16884 14868 16894
rect 13804 15374 13806 15426
rect 13858 15374 13860 15426
rect 13804 15362 13860 15374
rect 14812 15874 14868 16828
rect 15036 16212 15092 16222
rect 14812 15822 14814 15874
rect 14866 15822 14868 15874
rect 11676 15202 11732 15260
rect 11676 15150 11678 15202
rect 11730 15150 11732 15202
rect 11676 15138 11732 15150
rect 14588 15316 14644 15326
rect 14812 15316 14868 15822
rect 14588 15314 14868 15316
rect 14588 15262 14590 15314
rect 14642 15262 14868 15314
rect 14588 15260 14868 15262
rect 14924 16156 15036 16212
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 13132 14308 13188 14318
rect 13132 13858 13188 14252
rect 13132 13806 13134 13858
rect 13186 13806 13188 13858
rect 13132 13794 13188 13806
rect 12460 13748 12516 13758
rect 12460 13654 12516 13692
rect 14588 13748 14644 15260
rect 14924 15204 14980 16156
rect 15036 16146 15092 16156
rect 15148 16212 15204 17500
rect 15484 17442 15540 17500
rect 15484 17390 15486 17442
rect 15538 17390 15540 17442
rect 15484 17378 15540 17390
rect 15484 17220 15540 17230
rect 15372 17164 15484 17220
rect 15260 16882 15316 16894
rect 15260 16830 15262 16882
rect 15314 16830 15316 16882
rect 15260 16322 15316 16830
rect 15372 16772 15428 17164
rect 15484 17154 15540 17164
rect 15484 16996 15540 17006
rect 15484 16902 15540 16940
rect 15372 16716 15540 16772
rect 15260 16270 15262 16322
rect 15314 16270 15316 16322
rect 15260 16258 15316 16270
rect 15148 16146 15204 16156
rect 15372 15986 15428 15998
rect 15372 15934 15374 15986
rect 15426 15934 15428 15986
rect 15260 15876 15316 15886
rect 15260 15782 15316 15820
rect 15372 15540 15428 15934
rect 15148 15484 15428 15540
rect 15484 15876 15540 16716
rect 15484 15538 15540 15820
rect 15484 15486 15486 15538
rect 15538 15486 15540 15538
rect 15148 15428 15204 15484
rect 15484 15474 15540 15486
rect 15148 15334 15204 15372
rect 15260 15314 15316 15326
rect 15260 15262 15262 15314
rect 15314 15262 15316 15314
rect 15148 15204 15204 15214
rect 14700 15148 14980 15204
rect 15036 15202 15204 15204
rect 15036 15150 15150 15202
rect 15202 15150 15204 15202
rect 15036 15148 15204 15150
rect 14700 14418 14756 15148
rect 14924 14756 14980 14766
rect 15036 14756 15092 15148
rect 15148 15138 15204 15148
rect 14924 14754 15092 14756
rect 14924 14702 14926 14754
rect 14978 14702 15092 14754
rect 14924 14700 15092 14702
rect 14924 14690 14980 14700
rect 14700 14366 14702 14418
rect 14754 14366 14756 14418
rect 14700 14354 14756 14366
rect 14812 14308 14868 14318
rect 14812 14214 14868 14252
rect 14588 13412 14644 13692
rect 15260 13634 15316 15262
rect 15596 15314 15652 17612
rect 15708 17612 15988 17668
rect 16044 17724 16156 17780
rect 15708 16994 15764 17612
rect 15820 17444 15876 17454
rect 16044 17444 16100 17724
rect 16156 17714 16212 17724
rect 17052 17780 17108 21644
rect 17276 19908 17332 21980
rect 17388 21980 17668 22036
rect 17388 21810 17444 21980
rect 17948 21812 18004 21822
rect 17388 21758 17390 21810
rect 17442 21758 17444 21810
rect 17388 21746 17444 21758
rect 17612 21810 18004 21812
rect 17612 21758 17950 21810
rect 18002 21758 18004 21810
rect 17612 21756 18004 21758
rect 17500 21700 17556 21710
rect 17500 21606 17556 21644
rect 17612 20242 17668 21756
rect 17948 21746 18004 21756
rect 17836 21588 17892 21598
rect 17836 21494 17892 21532
rect 17612 20190 17614 20242
rect 17666 20190 17668 20242
rect 17388 20018 17444 20030
rect 17388 19966 17390 20018
rect 17442 19966 17444 20018
rect 17388 19908 17444 19966
rect 17164 19852 17444 19908
rect 17164 19012 17220 19852
rect 17276 19236 17332 19246
rect 17612 19236 17668 20190
rect 17724 20132 17780 20142
rect 18060 20132 18116 22540
rect 18172 21812 18228 22764
rect 18284 22594 18340 23772
rect 18284 22542 18286 22594
rect 18338 22542 18340 22594
rect 18284 22148 18340 22542
rect 18284 22082 18340 22092
rect 18396 23042 18452 23054
rect 18396 22990 18398 23042
rect 18450 22990 18452 23042
rect 18172 21756 18340 21812
rect 18172 21586 18228 21598
rect 18172 21534 18174 21586
rect 18226 21534 18228 21586
rect 18172 20580 18228 21534
rect 18172 20514 18228 20524
rect 17724 20130 18116 20132
rect 17724 20078 17726 20130
rect 17778 20078 18116 20130
rect 17724 20076 18116 20078
rect 17724 20066 17780 20076
rect 18284 19908 18340 21756
rect 18396 21700 18452 22990
rect 18620 22930 18676 22942
rect 18620 22878 18622 22930
rect 18674 22878 18676 22930
rect 18620 22596 18676 22878
rect 18620 22530 18676 22540
rect 18620 22148 18676 22158
rect 18396 21634 18452 21644
rect 18508 22146 18676 22148
rect 18508 22094 18622 22146
rect 18674 22094 18676 22146
rect 18508 22092 18676 22094
rect 18284 19842 18340 19852
rect 18508 19236 18564 22092
rect 18620 22082 18676 22092
rect 18620 21588 18676 21598
rect 18620 21494 18676 21532
rect 17276 19234 17668 19236
rect 17276 19182 17278 19234
rect 17330 19182 17668 19234
rect 17276 19180 17668 19182
rect 18172 19180 18564 19236
rect 18620 19236 18676 19246
rect 17276 19170 17332 19180
rect 17164 18956 17332 19012
rect 17052 17686 17108 17724
rect 16268 17666 16324 17678
rect 16268 17614 16270 17666
rect 16322 17614 16324 17666
rect 16268 17556 16324 17614
rect 16268 17490 16324 17500
rect 16492 17668 16548 17678
rect 16492 17554 16548 17612
rect 17164 17668 17220 17678
rect 17164 17574 17220 17612
rect 16492 17502 16494 17554
rect 16546 17502 16548 17554
rect 15820 17442 16100 17444
rect 15820 17390 15822 17442
rect 15874 17390 16100 17442
rect 15820 17388 16100 17390
rect 15820 17378 15876 17388
rect 15708 16942 15710 16994
rect 15762 16942 15764 16994
rect 15708 16930 15764 16942
rect 15932 16996 15988 17006
rect 15932 16902 15988 16940
rect 16380 16212 16436 16222
rect 16380 16098 16436 16156
rect 16380 16046 16382 16098
rect 16434 16046 16436 16098
rect 16380 15428 16436 16046
rect 16492 16100 16548 17502
rect 17276 17556 17332 18956
rect 17500 18452 17556 18462
rect 17500 18338 17556 18396
rect 17500 18286 17502 18338
rect 17554 18286 17556 18338
rect 17388 17556 17444 17566
rect 17276 17500 17388 17556
rect 17388 17490 17444 17500
rect 17500 16996 17556 18286
rect 17948 18452 18004 18462
rect 18172 18452 18228 19180
rect 18620 19142 18676 19180
rect 18508 19010 18564 19022
rect 18508 18958 18510 19010
rect 18562 18958 18564 19010
rect 18508 18676 18564 18958
rect 18396 18620 18564 18676
rect 18396 18452 18452 18620
rect 17948 18450 18228 18452
rect 17948 18398 17950 18450
rect 18002 18398 18228 18450
rect 17948 18396 18228 18398
rect 18284 18396 18452 18452
rect 18508 18452 18564 18462
rect 17948 17108 18004 18396
rect 18060 17892 18116 17902
rect 18060 17798 18116 17836
rect 18284 17668 18340 18396
rect 18508 18358 18564 18396
rect 18396 18228 18452 18238
rect 18396 18134 18452 18172
rect 18620 17780 18676 17790
rect 18284 17574 18340 17612
rect 18508 17666 18564 17678
rect 18508 17614 18510 17666
rect 18562 17614 18564 17666
rect 18508 17556 18564 17614
rect 18508 17490 18564 17500
rect 18620 17554 18676 17724
rect 18620 17502 18622 17554
rect 18674 17502 18676 17554
rect 18620 17490 18676 17502
rect 17948 17042 18004 17052
rect 17500 16930 17556 16940
rect 16604 16100 16660 16110
rect 16492 16098 16772 16100
rect 16492 16046 16606 16098
rect 16658 16046 16772 16098
rect 16492 16044 16772 16046
rect 16604 16034 16660 16044
rect 16492 15876 16548 15886
rect 16492 15782 16548 15820
rect 16716 15540 16772 16044
rect 17388 15540 17444 15550
rect 16716 15538 17444 15540
rect 16716 15486 16718 15538
rect 16770 15486 17390 15538
rect 17442 15486 17444 15538
rect 16716 15484 17444 15486
rect 16716 15474 16772 15484
rect 17388 15474 17444 15484
rect 16604 15428 16660 15438
rect 16380 15426 16660 15428
rect 16380 15374 16606 15426
rect 16658 15374 16660 15426
rect 16380 15372 16660 15374
rect 16604 15362 16660 15372
rect 17724 15428 17780 15438
rect 15596 15262 15598 15314
rect 15650 15262 15652 15314
rect 15596 14532 15652 15262
rect 16940 15314 16996 15326
rect 16940 15262 16942 15314
rect 16994 15262 16996 15314
rect 16940 15148 16996 15262
rect 16940 15092 17220 15148
rect 17052 14644 17108 14654
rect 16940 14588 17052 14644
rect 15596 14466 15652 14476
rect 16828 14532 16884 14542
rect 16828 14438 16884 14476
rect 16492 14420 16548 14430
rect 16268 14308 16324 14318
rect 16268 13858 16324 14252
rect 16268 13806 16270 13858
rect 16322 13806 16324 13858
rect 16268 13794 16324 13806
rect 16492 13746 16548 14364
rect 16828 13860 16884 13870
rect 16940 13860 16996 14588
rect 17052 14550 17108 14588
rect 17164 14532 17220 15092
rect 17164 14438 17220 14476
rect 17724 14532 17780 15372
rect 18844 15148 18900 24780
rect 18956 22932 19012 22942
rect 18956 22838 19012 22876
rect 18956 21588 19012 21598
rect 18956 21494 19012 21532
rect 19068 19796 19124 25004
rect 19516 23380 19572 26236
rect 21308 26178 21364 26852
rect 21420 26852 21812 26908
rect 21980 26962 22036 26974
rect 21980 26910 21982 26962
rect 22034 26910 22036 26962
rect 21868 26852 21924 26862
rect 21420 26514 21476 26852
rect 21868 26758 21924 26796
rect 21420 26462 21422 26514
rect 21474 26462 21476 26514
rect 21420 26450 21476 26462
rect 21308 26126 21310 26178
rect 21362 26126 21364 26178
rect 21308 26114 21364 26126
rect 21644 26068 21700 26078
rect 21980 26068 22036 26910
rect 22204 26964 22260 26974
rect 22204 26870 22260 26908
rect 22428 26962 22484 26974
rect 22428 26910 22430 26962
rect 22482 26910 22484 26962
rect 22428 26292 22484 26910
rect 22428 26226 22484 26236
rect 21644 26066 22036 26068
rect 21644 26014 21646 26066
rect 21698 26014 22036 26066
rect 21644 26012 22036 26014
rect 21644 26002 21700 26012
rect 21308 25508 21364 25518
rect 21308 25414 21364 25452
rect 21420 25282 21476 25294
rect 21420 25230 21422 25282
rect 21474 25230 21476 25282
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 21420 24388 21476 25230
rect 21420 24322 21476 24332
rect 21644 25282 21700 25294
rect 21644 25230 21646 25282
rect 21698 25230 21700 25282
rect 21308 23828 21364 23838
rect 21308 23734 21364 23772
rect 21644 23828 21700 25230
rect 21644 23762 21700 23772
rect 21420 23716 21476 23726
rect 21420 23622 21476 23660
rect 21532 23714 21588 23726
rect 21532 23662 21534 23714
rect 21586 23662 21588 23714
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 21532 23492 21588 23662
rect 19836 23482 20100 23492
rect 21196 23436 21588 23492
rect 19516 23314 19572 23324
rect 21084 23380 21140 23390
rect 21084 23286 21140 23324
rect 19740 23266 19796 23278
rect 19740 23214 19742 23266
rect 19794 23214 19796 23266
rect 19404 23156 19460 23166
rect 19068 19122 19124 19740
rect 19180 23154 19460 23156
rect 19180 23102 19406 23154
rect 19458 23102 19460 23154
rect 19180 23100 19460 23102
rect 19180 19236 19236 23100
rect 19404 23090 19460 23100
rect 19740 23156 19796 23214
rect 20412 23268 20468 23278
rect 20412 23174 20468 23212
rect 19740 23090 19796 23100
rect 20076 23154 20132 23166
rect 20076 23102 20078 23154
rect 20130 23102 20132 23154
rect 19964 22708 20020 22718
rect 19964 22594 20020 22652
rect 19964 22542 19966 22594
rect 20018 22542 20020 22594
rect 19964 22530 20020 22542
rect 20076 22596 20132 23102
rect 21196 23042 21252 23436
rect 21868 23380 21924 26012
rect 21980 24948 22036 24958
rect 21980 23938 22036 24892
rect 22316 24388 22372 24398
rect 22372 24332 22484 24388
rect 22316 24322 22372 24332
rect 21980 23886 21982 23938
rect 22034 23886 22036 23938
rect 21980 23874 22036 23886
rect 21980 23380 22036 23390
rect 21868 23378 22036 23380
rect 21868 23326 21982 23378
rect 22034 23326 22036 23378
rect 21868 23324 22036 23326
rect 21980 23314 22036 23324
rect 22204 23380 22260 23390
rect 21196 22990 21198 23042
rect 21250 22990 21252 23042
rect 21196 22978 21252 22990
rect 21644 23266 21700 23278
rect 21644 23214 21646 23266
rect 21698 23214 21700 23266
rect 20076 22530 20132 22540
rect 20412 22932 20468 22942
rect 19628 22370 19684 22382
rect 19628 22318 19630 22370
rect 19682 22318 19684 22370
rect 19292 22146 19348 22158
rect 19292 22094 19294 22146
rect 19346 22094 19348 22146
rect 19292 20244 19348 22094
rect 19404 22146 19460 22158
rect 19404 22094 19406 22146
rect 19458 22094 19460 22146
rect 19404 21140 19460 22094
rect 19516 22146 19572 22158
rect 19516 22094 19518 22146
rect 19570 22094 19572 22146
rect 19516 21476 19572 22094
rect 19516 21410 19572 21420
rect 19404 21084 19572 21140
rect 19292 20178 19348 20188
rect 19516 20130 19572 21084
rect 19516 20078 19518 20130
rect 19570 20078 19572 20130
rect 19516 20066 19572 20078
rect 19180 19170 19236 19180
rect 19292 19908 19348 19918
rect 19292 19684 19348 19852
rect 19292 19234 19348 19628
rect 19628 19348 19684 22318
rect 20412 22372 20468 22876
rect 20860 22930 20916 22942
rect 20860 22878 20862 22930
rect 20914 22878 20916 22930
rect 20860 22708 20916 22878
rect 20412 22370 20580 22372
rect 20412 22318 20414 22370
rect 20466 22318 20580 22370
rect 20412 22316 20580 22318
rect 20412 22306 20468 22316
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20076 20804 20132 20814
rect 20076 20710 20132 20748
rect 20188 20580 20244 20590
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20076 20018 20132 20030
rect 20076 19966 20078 20018
rect 20130 19966 20132 20018
rect 20076 19908 20132 19966
rect 20076 19842 20132 19852
rect 19628 19254 19684 19292
rect 19852 19572 19908 19582
rect 19292 19182 19294 19234
rect 19346 19182 19348 19234
rect 19292 19170 19348 19182
rect 19068 19070 19070 19122
rect 19122 19070 19124 19122
rect 19068 19012 19124 19070
rect 19852 19012 19908 19516
rect 20188 19234 20244 20524
rect 20524 20132 20580 22316
rect 20748 22148 20804 22158
rect 20860 22148 20916 22652
rect 21644 22596 21700 23214
rect 22092 23268 22148 23278
rect 22092 23174 22148 23212
rect 21644 22530 21700 22540
rect 21756 23156 21812 23166
rect 21868 23156 21924 23166
rect 21812 23154 21924 23156
rect 21812 23102 21870 23154
rect 21922 23102 21924 23154
rect 21812 23100 21924 23102
rect 21532 22372 21588 22382
rect 21756 22372 21812 23100
rect 21868 23090 21924 23100
rect 21532 22370 21812 22372
rect 21532 22318 21534 22370
rect 21586 22318 21812 22370
rect 21532 22316 21812 22318
rect 20748 22146 20916 22148
rect 20748 22094 20750 22146
rect 20802 22094 20916 22146
rect 20748 22092 20916 22094
rect 21308 22258 21364 22270
rect 21308 22206 21310 22258
rect 21362 22206 21364 22258
rect 20748 21924 20804 22092
rect 20748 21858 20804 21868
rect 20524 20066 20580 20076
rect 20972 20130 21028 20142
rect 20972 20078 20974 20130
rect 21026 20078 21028 20130
rect 20300 20020 20356 20030
rect 20300 19926 20356 19964
rect 20412 20018 20468 20030
rect 20412 19966 20414 20018
rect 20466 19966 20468 20018
rect 20412 19796 20468 19966
rect 20412 19730 20468 19740
rect 20636 19908 20692 19918
rect 20188 19182 20190 19234
rect 20242 19182 20244 19234
rect 20188 19170 20244 19182
rect 19068 18956 19572 19012
rect 19180 18562 19236 18574
rect 19180 18510 19182 18562
rect 19234 18510 19236 18562
rect 18956 18450 19012 18462
rect 18956 18398 18958 18450
rect 19010 18398 19012 18450
rect 18956 18228 19012 18398
rect 18956 18162 19012 18172
rect 19180 18452 19236 18510
rect 19180 17556 19236 18396
rect 19516 18450 19572 18956
rect 19628 18956 19908 19012
rect 19628 18564 19684 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 18470 19684 18508
rect 19516 18398 19518 18450
rect 19570 18398 19572 18450
rect 19516 18386 19572 18398
rect 20636 18450 20692 19852
rect 20972 19572 21028 20078
rect 20972 19506 21028 19516
rect 20636 18398 20638 18450
rect 20690 18398 20692 18450
rect 20636 18386 20692 18398
rect 21196 18562 21252 18574
rect 21196 18510 21198 18562
rect 21250 18510 21252 18562
rect 20300 18340 20356 18350
rect 20300 18338 20468 18340
rect 20300 18286 20302 18338
rect 20354 18286 20468 18338
rect 20300 18284 20468 18286
rect 20300 18274 20356 18284
rect 19516 17668 19572 17678
rect 19180 17108 19236 17500
rect 19404 17554 19460 17566
rect 19404 17502 19406 17554
rect 19458 17502 19460 17554
rect 19292 17108 19348 17118
rect 19180 17106 19348 17108
rect 19180 17054 19294 17106
rect 19346 17054 19348 17106
rect 19180 17052 19348 17054
rect 19292 17042 19348 17052
rect 19404 16884 19460 17502
rect 19516 16996 19572 17612
rect 20076 17556 20132 17566
rect 20300 17556 20356 17566
rect 20132 17500 20244 17556
rect 20076 17462 20132 17500
rect 19516 16930 19572 16940
rect 19628 17444 19684 17454
rect 19628 17106 19684 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 17054 19630 17106
rect 19682 17054 19684 17106
rect 19404 16818 19460 16828
rect 19628 16660 19684 17054
rect 20188 17106 20244 17500
rect 20188 17054 20190 17106
rect 20242 17054 20244 17106
rect 20188 17042 20244 17054
rect 19404 16604 19684 16660
rect 19964 16996 20020 17006
rect 18620 15092 18900 15148
rect 19180 15988 19236 15998
rect 18396 14756 18452 14766
rect 18396 14662 18452 14700
rect 18284 14532 18340 14542
rect 17724 14530 18340 14532
rect 17724 14478 17726 14530
rect 17778 14478 18286 14530
rect 18338 14478 18340 14530
rect 17724 14476 18340 14478
rect 17724 14466 17780 14476
rect 18284 14466 18340 14476
rect 18620 14530 18676 15092
rect 19180 14754 19236 15932
rect 19404 15148 19460 16604
rect 19964 16098 20020 16940
rect 20300 16770 20356 17500
rect 20300 16718 20302 16770
rect 20354 16718 20356 16770
rect 20300 16706 20356 16718
rect 19964 16046 19966 16098
rect 20018 16046 20020 16098
rect 19964 16034 20020 16046
rect 19628 15988 19684 15998
rect 19628 15894 19684 15932
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19404 15092 19572 15148
rect 19180 14702 19182 14754
rect 19234 14702 19236 14754
rect 19180 14690 19236 14702
rect 18620 14478 18622 14530
rect 18674 14478 18676 14530
rect 18620 14466 18676 14478
rect 18956 14532 19012 14542
rect 18956 14438 19012 14476
rect 19516 14530 19572 15092
rect 19516 14478 19518 14530
rect 19570 14478 19572 14530
rect 19516 14466 19572 14478
rect 19628 14754 19684 14766
rect 19628 14702 19630 14754
rect 19682 14702 19684 14754
rect 17388 14308 17444 14318
rect 17388 14214 17444 14252
rect 17612 14308 17668 14318
rect 17612 14306 17892 14308
rect 17612 14254 17614 14306
rect 17666 14254 17892 14306
rect 17612 14252 17892 14254
rect 17612 14242 17668 14252
rect 16828 13858 16996 13860
rect 16828 13806 16830 13858
rect 16882 13806 16996 13858
rect 16828 13804 16996 13806
rect 16828 13794 16884 13804
rect 16492 13694 16494 13746
rect 16546 13694 16548 13746
rect 16492 13682 16548 13694
rect 15260 13582 15262 13634
rect 15314 13582 15316 13634
rect 14700 13412 14756 13422
rect 4476 13356 4740 13366
rect 14588 13356 14700 13412
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 14700 12962 14756 13356
rect 14700 12910 14702 12962
rect 14754 12910 14756 12962
rect 14700 12898 14756 12910
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 15260 11284 15316 13582
rect 15708 13634 15764 13646
rect 15708 13582 15710 13634
rect 15762 13582 15764 13634
rect 15484 13522 15540 13534
rect 15484 13470 15486 13522
rect 15538 13470 15540 13522
rect 15372 13076 15428 13086
rect 15484 13076 15540 13470
rect 15708 13524 15764 13582
rect 16380 13634 16436 13646
rect 17500 13636 17556 13646
rect 16380 13582 16382 13634
rect 16434 13582 16436 13634
rect 15708 13458 15764 13468
rect 16044 13524 16100 13534
rect 16380 13524 16436 13582
rect 16044 13522 16436 13524
rect 16044 13470 16046 13522
rect 16098 13470 16436 13522
rect 16044 13468 16436 13470
rect 17388 13580 17500 13636
rect 16044 13458 16100 13468
rect 15372 13074 15540 13076
rect 15372 13022 15374 13074
rect 15426 13022 15540 13074
rect 15372 13020 15540 13022
rect 15372 13010 15428 13020
rect 15260 11228 15652 11284
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 15484 5236 15540 5246
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 15484 800 15540 5180
rect 15596 5124 15652 11228
rect 16716 5236 16772 5246
rect 16716 5142 16772 5180
rect 15708 5124 15764 5134
rect 15596 5122 15764 5124
rect 15596 5070 15710 5122
rect 15762 5070 15764 5122
rect 15596 5068 15764 5070
rect 15708 5058 15764 5068
rect 17388 4340 17444 13580
rect 17500 13542 17556 13580
rect 17500 13076 17556 13086
rect 17836 13076 17892 14252
rect 18060 14306 18116 14318
rect 18060 14254 18062 14306
rect 18114 14254 18116 14306
rect 18060 13636 18116 14254
rect 19628 13858 19684 14702
rect 19740 14756 19796 14766
rect 19740 14662 19796 14700
rect 20412 14530 20468 18284
rect 20860 18116 20916 18126
rect 20860 17666 20916 18060
rect 21196 17780 21252 18510
rect 21308 18228 21364 22206
rect 21532 22148 21588 22316
rect 21532 22082 21588 22092
rect 21868 22260 21924 22270
rect 22204 22260 22260 23324
rect 21868 22146 21924 22204
rect 21868 22094 21870 22146
rect 21922 22094 21924 22146
rect 21868 22082 21924 22094
rect 21980 22258 22260 22260
rect 21980 22206 22206 22258
rect 22258 22206 22260 22258
rect 21980 22204 22260 22206
rect 21980 21924 22036 22204
rect 22204 22194 22260 22204
rect 21756 21868 22036 21924
rect 22092 21924 22148 21934
rect 21756 20690 21812 21868
rect 22092 21812 22148 21868
rect 21756 20638 21758 20690
rect 21810 20638 21812 20690
rect 21756 20626 21812 20638
rect 21980 21756 22148 21812
rect 21980 20802 22036 21756
rect 21980 20750 21982 20802
rect 22034 20750 22036 20802
rect 21532 20580 21588 20590
rect 21532 20578 21700 20580
rect 21532 20526 21534 20578
rect 21586 20526 21700 20578
rect 21532 20524 21700 20526
rect 21532 20514 21588 20524
rect 21420 20244 21476 20254
rect 21420 19906 21476 20188
rect 21532 20132 21588 20142
rect 21532 20038 21588 20076
rect 21420 19854 21422 19906
rect 21474 19854 21476 19906
rect 21420 19842 21476 19854
rect 21532 19684 21588 19694
rect 21644 19684 21700 20524
rect 21756 19796 21812 19806
rect 21756 19702 21812 19740
rect 21588 19628 21700 19684
rect 21532 19618 21588 19628
rect 21308 18162 21364 18172
rect 21532 18676 21588 18686
rect 21532 18450 21588 18620
rect 21980 18676 22036 20750
rect 22316 20914 22372 20926
rect 22316 20862 22318 20914
rect 22370 20862 22372 20914
rect 22092 20690 22148 20702
rect 22092 20638 22094 20690
rect 22146 20638 22148 20690
rect 22092 20132 22148 20638
rect 22092 20066 22148 20076
rect 22204 20130 22260 20142
rect 22204 20078 22206 20130
rect 22258 20078 22260 20130
rect 22092 19908 22148 19918
rect 22092 19814 22148 19852
rect 22092 19684 22148 19694
rect 22204 19684 22260 20078
rect 22148 19628 22260 19684
rect 22092 19618 22148 19628
rect 22204 19460 22260 19470
rect 21980 18610 22036 18620
rect 22092 19404 22204 19460
rect 22092 18674 22148 19404
rect 22204 19394 22260 19404
rect 22316 19234 22372 20862
rect 22428 20132 22484 24332
rect 22764 23938 22820 27022
rect 24444 27746 24612 27748
rect 24444 27694 24558 27746
rect 24610 27694 24612 27746
rect 24444 27692 24612 27694
rect 23548 26962 23604 26974
rect 23548 26910 23550 26962
rect 23602 26910 23604 26962
rect 23436 26852 23492 26862
rect 23436 26292 23492 26796
rect 23548 26514 23604 26910
rect 23548 26462 23550 26514
rect 23602 26462 23604 26514
rect 23548 26450 23604 26462
rect 24444 26514 24500 27692
rect 24556 27682 24612 27692
rect 25228 27748 25284 27758
rect 25340 27748 25396 27806
rect 25284 27692 25620 27748
rect 25228 27682 25284 27692
rect 24444 26462 24446 26514
rect 24498 26462 24500 26514
rect 24444 26450 24500 26462
rect 25452 26964 25508 26974
rect 23436 26290 23604 26292
rect 23436 26238 23438 26290
rect 23490 26238 23604 26290
rect 23436 26236 23604 26238
rect 23436 26226 23492 26236
rect 23548 24052 23604 26236
rect 23660 26290 23716 26302
rect 23660 26238 23662 26290
rect 23714 26238 23716 26290
rect 23660 24948 23716 26238
rect 23996 26292 24052 26302
rect 23996 26290 24276 26292
rect 23996 26238 23998 26290
rect 24050 26238 24276 26290
rect 23996 26236 24276 26238
rect 23996 26226 24052 26236
rect 24220 25620 24276 26236
rect 24332 26290 24388 26302
rect 24332 26238 24334 26290
rect 24386 26238 24388 26290
rect 24332 25844 24388 26238
rect 24444 26292 24500 26302
rect 24444 26066 24500 26236
rect 24444 26014 24446 26066
rect 24498 26014 24500 26066
rect 24444 26002 24500 26014
rect 25452 25956 25508 26908
rect 25564 26290 25620 27692
rect 25564 26238 25566 26290
rect 25618 26238 25620 26290
rect 25564 26226 25620 26238
rect 25676 27186 25732 31892
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 25788 27748 25844 27758
rect 25844 27692 26180 27748
rect 25788 27682 25844 27692
rect 25676 27134 25678 27186
rect 25730 27134 25732 27186
rect 25452 25890 25508 25900
rect 24332 25788 24612 25844
rect 24444 25620 24500 25630
rect 24220 25618 24500 25620
rect 24220 25566 24446 25618
rect 24498 25566 24500 25618
rect 24220 25564 24500 25566
rect 24444 25554 24500 25564
rect 24332 25396 24388 25406
rect 24556 25396 24612 25788
rect 24668 25508 24724 25518
rect 24668 25414 24724 25452
rect 25676 25508 25732 27134
rect 26124 27188 26180 27692
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 26124 27186 26516 27188
rect 26124 27134 26126 27186
rect 26178 27134 26516 27186
rect 26124 27132 26516 27134
rect 26124 27122 26180 27132
rect 26348 26180 26404 26190
rect 25788 26178 26404 26180
rect 25788 26126 26350 26178
rect 26402 26126 26404 26178
rect 25788 26124 26404 26126
rect 25788 25618 25844 26124
rect 26348 26114 26404 26124
rect 25788 25566 25790 25618
rect 25842 25566 25844 25618
rect 25788 25554 25844 25566
rect 25900 25956 25956 25966
rect 25676 25442 25732 25452
rect 25900 25506 25956 25900
rect 25900 25454 25902 25506
rect 25954 25454 25956 25506
rect 25900 25442 25956 25454
rect 24332 25394 24612 25396
rect 24332 25342 24334 25394
rect 24386 25342 24612 25394
rect 24332 25340 24612 25342
rect 24892 25394 24948 25406
rect 24892 25342 24894 25394
rect 24946 25342 24948 25394
rect 24332 25060 24388 25340
rect 24108 25004 24388 25060
rect 24892 25284 24948 25342
rect 26124 25396 26180 25406
rect 26124 25302 26180 25340
rect 23716 24892 23940 24948
rect 23660 24882 23716 24892
rect 22764 23886 22766 23938
rect 22818 23886 22820 23938
rect 22764 23874 22820 23886
rect 23436 23996 23604 24052
rect 23436 23604 23492 23996
rect 23548 23826 23604 23838
rect 23548 23774 23550 23826
rect 23602 23774 23604 23826
rect 23548 23716 23604 23774
rect 23660 23716 23716 23726
rect 23548 23660 23660 23716
rect 23660 23650 23716 23660
rect 23436 23548 23604 23604
rect 23212 22260 23268 22270
rect 23212 22166 23268 22204
rect 22540 22148 22596 22158
rect 22540 20244 22596 22092
rect 22876 22148 22932 22158
rect 22876 22146 23044 22148
rect 22876 22094 22878 22146
rect 22930 22094 23044 22146
rect 22876 22092 23044 22094
rect 22876 22082 22932 22092
rect 22652 21474 22708 21486
rect 22652 21422 22654 21474
rect 22706 21422 22708 21474
rect 22652 20804 22708 21422
rect 22652 20710 22708 20748
rect 22876 20244 22932 20254
rect 22540 20242 22932 20244
rect 22540 20190 22878 20242
rect 22930 20190 22932 20242
rect 22540 20188 22932 20190
rect 22876 20178 22932 20188
rect 22428 20076 22596 20132
rect 22428 19908 22484 19918
rect 22428 19814 22484 19852
rect 22540 19460 22596 20076
rect 22764 20020 22820 20030
rect 22764 19926 22820 19964
rect 22876 19908 22932 19918
rect 22988 19908 23044 22092
rect 23436 20132 23492 20142
rect 23436 20038 23492 20076
rect 22932 19852 23044 19908
rect 23100 20018 23156 20030
rect 23100 19966 23102 20018
rect 23154 19966 23156 20018
rect 22876 19842 22932 19852
rect 23100 19460 23156 19966
rect 22540 19394 22596 19404
rect 22652 19404 23156 19460
rect 22428 19348 22484 19358
rect 22428 19254 22484 19292
rect 22316 19182 22318 19234
rect 22370 19182 22372 19234
rect 22316 19170 22372 19182
rect 22540 19234 22596 19246
rect 22540 19182 22542 19234
rect 22594 19182 22596 19234
rect 22092 18622 22094 18674
rect 22146 18622 22148 18674
rect 21868 18564 21924 18574
rect 21532 18398 21534 18450
rect 21586 18398 21588 18450
rect 21196 17714 21252 17724
rect 20860 17614 20862 17666
rect 20914 17614 20916 17666
rect 20860 17602 20916 17614
rect 21532 17666 21588 18398
rect 21532 17614 21534 17666
rect 21586 17614 21588 17666
rect 20524 17556 20580 17566
rect 20524 17462 20580 17500
rect 20636 17442 20692 17454
rect 20636 17390 20638 17442
rect 20690 17390 20692 17442
rect 20636 17108 20692 17390
rect 21532 17332 21588 17614
rect 21756 18562 21924 18564
rect 21756 18510 21870 18562
rect 21922 18510 21924 18562
rect 21756 18508 21924 18510
rect 21644 17556 21700 17566
rect 21644 17462 21700 17500
rect 21532 17276 21700 17332
rect 20524 17052 20692 17108
rect 20860 17108 20916 17118
rect 20524 16772 20580 17052
rect 20636 16884 20692 16894
rect 20636 16790 20692 16828
rect 20860 16882 20916 17052
rect 21196 17108 21252 17118
rect 21196 17014 21252 17052
rect 20860 16830 20862 16882
rect 20914 16830 20916 16882
rect 20860 16818 20916 16830
rect 21420 16884 21476 16894
rect 20524 15876 20580 16716
rect 20524 15810 20580 15820
rect 21420 15148 21476 16828
rect 21532 16882 21588 16894
rect 21532 16830 21534 16882
rect 21586 16830 21588 16882
rect 21532 16772 21588 16830
rect 21532 16706 21588 16716
rect 21644 16098 21700 17276
rect 21644 16046 21646 16098
rect 21698 16046 21700 16098
rect 21644 16034 21700 16046
rect 21756 17106 21812 18508
rect 21868 18498 21924 18508
rect 22092 18452 22148 18622
rect 21980 18396 22148 18452
rect 21868 17780 21924 17790
rect 21868 17686 21924 17724
rect 21756 17054 21758 17106
rect 21810 17054 21812 17106
rect 21756 15988 21812 17054
rect 21756 15894 21812 15932
rect 21868 17442 21924 17454
rect 21868 17390 21870 17442
rect 21922 17390 21924 17442
rect 21868 15148 21924 17390
rect 21980 17444 22036 18396
rect 22204 18228 22260 18238
rect 22204 18134 22260 18172
rect 22540 17780 22596 19182
rect 22428 17724 22596 17780
rect 22652 17778 22708 19404
rect 22764 19234 22820 19246
rect 22764 19182 22766 19234
rect 22818 19182 22820 19234
rect 22764 18004 22820 19182
rect 23100 18562 23156 19404
rect 23324 19234 23380 19246
rect 23324 19182 23326 19234
rect 23378 19182 23380 19234
rect 23324 19012 23380 19182
rect 23324 18946 23380 18956
rect 23548 18674 23604 23548
rect 23660 23492 23716 23502
rect 23660 23378 23716 23436
rect 23660 23326 23662 23378
rect 23714 23326 23716 23378
rect 23660 23314 23716 23326
rect 23884 23378 23940 24892
rect 23996 24836 24052 24846
rect 24108 24836 24164 25004
rect 24052 24780 24164 24836
rect 24220 24836 24276 24846
rect 23996 24742 24052 24780
rect 24108 24610 24164 24622
rect 24108 24558 24110 24610
rect 24162 24558 24164 24610
rect 23884 23326 23886 23378
rect 23938 23326 23940 23378
rect 23884 23314 23940 23326
rect 23996 23716 24052 23726
rect 23996 23378 24052 23660
rect 23996 23326 23998 23378
rect 24050 23326 24052 23378
rect 23996 23314 24052 23326
rect 24108 23378 24164 24558
rect 24220 23604 24276 24780
rect 24332 24724 24388 24734
rect 24332 24630 24388 24668
rect 24556 24722 24612 24734
rect 24556 24670 24558 24722
rect 24610 24670 24612 24722
rect 24220 23538 24276 23548
rect 24108 23326 24110 23378
rect 24162 23326 24164 23378
rect 24108 23314 24164 23326
rect 24220 23268 24276 23278
rect 23884 22370 23940 22382
rect 23884 22318 23886 22370
rect 23938 22318 23940 22370
rect 23884 22260 23940 22318
rect 24220 22372 24276 23212
rect 24556 23044 24612 24670
rect 24556 22978 24612 22988
rect 24220 22278 24276 22316
rect 24892 22482 24948 25228
rect 25564 25284 25620 25294
rect 25564 25190 25620 25228
rect 25676 25284 25732 25294
rect 25676 25282 25844 25284
rect 25676 25230 25678 25282
rect 25730 25230 25844 25282
rect 25676 25228 25844 25230
rect 25676 25218 25732 25228
rect 25676 24724 25732 24734
rect 25676 24052 25732 24668
rect 25676 23958 25732 23996
rect 25788 23828 25844 25228
rect 26460 24946 26516 27132
rect 40012 27186 40068 27198
rect 40012 27134 40014 27186
rect 40066 27134 40068 27186
rect 37660 27074 37716 27086
rect 37660 27022 37662 27074
rect 37714 27022 37716 27074
rect 27468 26180 27524 26190
rect 27244 25396 27300 25406
rect 27244 25302 27300 25340
rect 27468 25394 27524 26124
rect 28476 26180 28532 26190
rect 28476 26086 28532 26124
rect 28924 26178 28980 26190
rect 28924 26126 28926 26178
rect 28978 26126 28980 26178
rect 27468 25342 27470 25394
rect 27522 25342 27524 25394
rect 27468 25330 27524 25342
rect 27580 25394 27636 25406
rect 27580 25342 27582 25394
rect 27634 25342 27636 25394
rect 26460 24894 26462 24946
rect 26514 24894 26516 24946
rect 26460 24724 26516 24894
rect 26908 24836 26964 24846
rect 26908 24742 26964 24780
rect 26124 24668 26460 24724
rect 26124 24050 26180 24668
rect 26460 24658 26516 24668
rect 26796 24724 26852 24734
rect 26124 23998 26126 24050
rect 26178 23998 26180 24050
rect 26124 23986 26180 23998
rect 26684 24052 26740 24062
rect 26796 24052 26852 24668
rect 27020 24724 27076 24734
rect 27356 24724 27412 24734
rect 27020 24722 27300 24724
rect 27020 24670 27022 24722
rect 27074 24670 27300 24722
rect 27020 24668 27300 24670
rect 27020 24658 27076 24668
rect 26908 24500 26964 24510
rect 26908 24498 27188 24500
rect 26908 24446 26910 24498
rect 26962 24446 27188 24498
rect 26908 24444 27188 24446
rect 26908 24434 26964 24444
rect 26684 24050 27076 24052
rect 26684 23998 26686 24050
rect 26738 23998 27076 24050
rect 26684 23996 27076 23998
rect 26684 23986 26740 23996
rect 25788 23772 26292 23828
rect 26124 23154 26180 23166
rect 26124 23102 26126 23154
rect 26178 23102 26180 23154
rect 25340 23044 25396 23054
rect 24892 22430 24894 22482
rect 24946 22430 24948 22482
rect 23884 22194 23940 22204
rect 23996 19348 24052 19358
rect 23996 19254 24052 19292
rect 23548 18622 23550 18674
rect 23602 18622 23604 18674
rect 23548 18610 23604 18622
rect 23100 18510 23102 18562
rect 23154 18510 23156 18562
rect 23100 18498 23156 18510
rect 23324 18562 23380 18574
rect 23324 18510 23326 18562
rect 23378 18510 23380 18562
rect 22876 18450 22932 18462
rect 22876 18398 22878 18450
rect 22930 18398 22932 18450
rect 22876 18340 22932 18398
rect 23324 18340 23380 18510
rect 22876 18284 23156 18340
rect 22764 17938 22820 17948
rect 22876 17892 22932 17902
rect 22876 17798 22932 17836
rect 23100 17892 23156 18284
rect 23324 18274 23380 18284
rect 23996 18340 24052 18350
rect 24332 18340 24388 18350
rect 24052 18284 24164 18340
rect 23996 18274 24052 18284
rect 23884 18228 23940 18238
rect 22652 17726 22654 17778
rect 22706 17726 22708 17778
rect 22092 17668 22148 17678
rect 22092 17574 22148 17612
rect 21980 17106 22036 17388
rect 21980 17054 21982 17106
rect 22034 17054 22036 17106
rect 21980 17042 22036 17054
rect 22092 17108 22148 17118
rect 22428 17108 22484 17724
rect 22092 17106 22484 17108
rect 22092 17054 22094 17106
rect 22146 17054 22484 17106
rect 22092 17052 22484 17054
rect 22540 17556 22596 17566
rect 22652 17556 22708 17726
rect 22652 17500 23044 17556
rect 22092 17042 22148 17052
rect 22540 16884 22596 17500
rect 22988 17106 23044 17500
rect 22988 17054 22990 17106
rect 23042 17054 23044 17106
rect 22988 17042 23044 17054
rect 22764 16996 22820 17006
rect 22764 16902 22820 16940
rect 22204 16882 22596 16884
rect 22204 16830 22542 16882
rect 22594 16830 22596 16882
rect 22204 16828 22596 16830
rect 22204 16548 22260 16828
rect 22540 16818 22596 16828
rect 22876 16884 22932 16894
rect 22876 16770 22932 16828
rect 23100 16882 23156 17836
rect 23436 18004 23492 18014
rect 23212 17444 23268 17454
rect 23212 17350 23268 17388
rect 23436 17108 23492 17948
rect 23884 17892 23940 18172
rect 23884 17836 24052 17892
rect 23772 17666 23828 17678
rect 23772 17614 23774 17666
rect 23826 17614 23828 17666
rect 23772 17444 23828 17614
rect 23772 17378 23828 17388
rect 23884 17666 23940 17678
rect 23884 17614 23886 17666
rect 23938 17614 23940 17666
rect 23436 17042 23492 17052
rect 23772 17108 23828 17118
rect 23884 17108 23940 17614
rect 23996 17666 24052 17836
rect 23996 17614 23998 17666
rect 24050 17614 24052 17666
rect 23996 17602 24052 17614
rect 23828 17052 23940 17108
rect 23100 16830 23102 16882
rect 23154 16830 23156 16882
rect 23100 16818 23156 16830
rect 23548 16884 23604 16894
rect 23548 16790 23604 16828
rect 22876 16718 22878 16770
rect 22930 16718 22932 16770
rect 22876 16706 22932 16718
rect 23772 16658 23828 17052
rect 24108 16994 24164 18284
rect 24332 17666 24388 18284
rect 24332 17614 24334 17666
rect 24386 17614 24388 17666
rect 24332 17602 24388 17614
rect 24220 17556 24276 17566
rect 24220 17462 24276 17500
rect 24108 16942 24110 16994
rect 24162 16942 24164 16994
rect 24108 16930 24164 16942
rect 24332 17444 24388 17454
rect 24332 16994 24388 17388
rect 24332 16942 24334 16994
rect 24386 16942 24388 16994
rect 24332 16930 24388 16942
rect 23772 16606 23774 16658
rect 23826 16606 23828 16658
rect 23772 16594 23828 16606
rect 24220 16770 24276 16782
rect 24220 16718 24222 16770
rect 24274 16718 24276 16770
rect 21980 16492 22260 16548
rect 21980 16098 22036 16492
rect 24220 16212 24276 16718
rect 24780 16212 24836 16222
rect 24220 16210 24836 16212
rect 24220 16158 24782 16210
rect 24834 16158 24836 16210
rect 24220 16156 24836 16158
rect 24780 16146 24836 16156
rect 21980 16046 21982 16098
rect 22034 16046 22036 16098
rect 21980 16034 22036 16046
rect 23996 16098 24052 16110
rect 23996 16046 23998 16098
rect 24050 16046 24052 16098
rect 21420 15092 21812 15148
rect 21868 15092 23156 15148
rect 23996 15092 24052 16046
rect 24892 15148 24948 22430
rect 25228 22596 25284 22606
rect 25228 22370 25284 22540
rect 25228 22318 25230 22370
rect 25282 22318 25284 22370
rect 25228 22260 25284 22318
rect 25228 22194 25284 22204
rect 25340 21810 25396 22988
rect 25340 21758 25342 21810
rect 25394 21758 25396 21810
rect 25340 21746 25396 21758
rect 25452 22372 25508 22382
rect 25452 21810 25508 22316
rect 26124 22372 26180 23102
rect 26124 22306 26180 22316
rect 25452 21758 25454 21810
rect 25506 21758 25508 21810
rect 25452 21746 25508 21758
rect 25228 21362 25284 21374
rect 25228 21310 25230 21362
rect 25282 21310 25284 21362
rect 25228 19908 25284 21310
rect 25228 18674 25284 19852
rect 26124 20132 26180 20142
rect 26124 19348 26180 20076
rect 26236 19908 26292 23772
rect 26460 23380 26516 23390
rect 26460 23286 26516 23324
rect 27020 23156 27076 23996
rect 27132 23268 27188 24444
rect 27244 23492 27300 24668
rect 27356 24630 27412 24668
rect 27580 23716 27636 25342
rect 28924 24724 28980 26126
rect 37660 26180 37716 27022
rect 40012 26292 40068 27134
rect 40012 26226 40068 26236
rect 37660 26114 37716 26124
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 40012 25618 40068 25630
rect 40012 25566 40014 25618
rect 40066 25566 40068 25618
rect 37660 25508 37716 25518
rect 37436 25506 37716 25508
rect 37436 25454 37662 25506
rect 37714 25454 37716 25506
rect 37436 25452 37716 25454
rect 30940 24836 30996 24846
rect 30940 24742 30996 24780
rect 30716 24724 30772 24734
rect 28924 24658 28980 24668
rect 30268 24668 30716 24724
rect 28140 24610 28196 24622
rect 28140 24558 28142 24610
rect 28194 24558 28196 24610
rect 28028 24164 28084 24174
rect 28140 24164 28196 24558
rect 28028 24162 28196 24164
rect 28028 24110 28030 24162
rect 28082 24110 28196 24162
rect 28028 24108 28196 24110
rect 30268 24610 30324 24668
rect 30716 24630 30772 24668
rect 37436 24724 37492 25452
rect 37660 25442 37716 25452
rect 40012 24948 40068 25566
rect 40012 24882 40068 24892
rect 37436 24658 37492 24668
rect 37660 24724 37716 24734
rect 37660 24630 37716 24668
rect 30268 24558 30270 24610
rect 30322 24558 30324 24610
rect 28028 24098 28084 24108
rect 29260 24050 29316 24062
rect 29260 23998 29262 24050
rect 29314 23998 29316 24050
rect 28140 23940 28196 23950
rect 28140 23846 28196 23884
rect 29036 23938 29092 23950
rect 29036 23886 29038 23938
rect 29090 23886 29092 23938
rect 28028 23828 28084 23838
rect 28028 23734 28084 23772
rect 27580 23650 27636 23660
rect 27244 23436 28308 23492
rect 27132 23202 27188 23212
rect 27804 23268 27860 23278
rect 27804 23174 27860 23212
rect 26908 23154 27076 23156
rect 26908 23102 27022 23154
rect 27074 23102 27076 23154
rect 26908 23100 27076 23102
rect 26684 22260 26740 22270
rect 26684 22166 26740 22204
rect 26908 21812 26964 23100
rect 27020 23090 27076 23100
rect 28252 22594 28308 23436
rect 29036 23380 29092 23886
rect 29260 23940 29316 23998
rect 29260 23874 29316 23884
rect 29596 23828 29652 23838
rect 29596 23734 29652 23772
rect 30268 23828 30324 24558
rect 40012 24498 40068 24510
rect 40012 24446 40014 24498
rect 40066 24446 40068 24498
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 40012 24276 40068 24446
rect 40012 24210 40068 24220
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 37660 23940 37716 23950
rect 37660 23846 37716 23884
rect 30268 23762 30324 23772
rect 28252 22542 28254 22594
rect 28306 22542 28308 22594
rect 28252 22530 28308 22542
rect 28588 23044 28644 23054
rect 27020 22372 27076 22382
rect 27020 22258 27076 22316
rect 28364 22372 28420 22382
rect 28364 22278 28420 22316
rect 27020 22206 27022 22258
rect 27074 22206 27076 22258
rect 27020 22194 27076 22206
rect 28140 22260 28196 22270
rect 28140 22166 28196 22204
rect 28588 22258 28644 22988
rect 28588 22206 28590 22258
rect 28642 22206 28644 22258
rect 28588 22194 28644 22206
rect 29036 22260 29092 23324
rect 26908 21810 27300 21812
rect 26908 21758 26910 21810
rect 26962 21758 27300 21810
rect 26908 21756 27300 21758
rect 26796 20690 26852 20702
rect 26796 20638 26798 20690
rect 26850 20638 26852 20690
rect 26796 20188 26852 20638
rect 26908 20188 26964 21756
rect 27244 21586 27300 21756
rect 27244 21534 27246 21586
rect 27298 21534 27300 21586
rect 27244 21522 27300 21534
rect 28028 21476 28084 21486
rect 28028 21474 28196 21476
rect 28028 21422 28030 21474
rect 28082 21422 28196 21474
rect 28028 21420 28196 21422
rect 28028 21410 28084 21420
rect 28140 20802 28196 21420
rect 28140 20750 28142 20802
rect 28194 20750 28196 20802
rect 28140 20738 28196 20750
rect 28476 20916 28532 20926
rect 28476 20802 28532 20860
rect 28476 20750 28478 20802
rect 28530 20750 28532 20802
rect 28476 20738 28532 20750
rect 28588 20804 28644 20814
rect 28364 20580 28420 20590
rect 28364 20486 28420 20524
rect 28588 20188 28644 20748
rect 29036 20802 29092 22204
rect 29372 23714 29428 23726
rect 29372 23662 29374 23714
rect 29426 23662 29428 23714
rect 29372 22372 29428 23662
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 37660 23156 37716 23166
rect 37660 23062 37716 23100
rect 29932 23044 29988 23054
rect 29932 22950 29988 22988
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 29260 20916 29316 20926
rect 29260 20822 29316 20860
rect 29036 20750 29038 20802
rect 29090 20750 29092 20802
rect 29036 20738 29092 20750
rect 29372 20804 29428 22316
rect 37884 22370 37940 22382
rect 37884 22318 37886 22370
rect 37938 22318 37940 22370
rect 37660 21586 37716 21598
rect 37660 21534 37662 21586
rect 37714 21534 37716 21586
rect 29372 20710 29428 20748
rect 29596 21476 29652 21486
rect 29596 20690 29652 21420
rect 30156 21476 30212 21486
rect 30156 21382 30212 21420
rect 37436 21476 37492 21486
rect 37660 21476 37716 21534
rect 37436 21474 37716 21476
rect 37436 21422 37438 21474
rect 37490 21422 37716 21474
rect 37436 21420 37716 21422
rect 37884 21476 37940 22318
rect 40012 21588 40068 22430
rect 40012 21522 40068 21532
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 29596 20638 29598 20690
rect 29650 20638 29652 20690
rect 29596 20626 29652 20638
rect 26796 20132 26964 20188
rect 27132 20132 27188 20142
rect 26572 20020 26628 20030
rect 26572 19908 26628 19964
rect 26236 19852 26628 19908
rect 26124 19254 26180 19292
rect 25228 18622 25230 18674
rect 25282 18622 25284 18674
rect 25228 18610 25284 18622
rect 25452 18676 25508 18686
rect 25452 18582 25508 18620
rect 25900 18452 25956 18462
rect 25900 18358 25956 18396
rect 25340 18340 25396 18350
rect 25340 18246 25396 18284
rect 26460 18116 26516 19852
rect 26572 19012 26628 19022
rect 26572 18452 26628 18956
rect 26796 18452 26852 20132
rect 27132 20038 27188 20076
rect 28364 20130 28420 20142
rect 28364 20078 28366 20130
rect 28418 20078 28420 20130
rect 27356 20020 27412 20030
rect 27356 19926 27412 19964
rect 27804 20020 27860 20030
rect 28140 20020 28196 20030
rect 27804 20018 28196 20020
rect 27804 19966 27806 20018
rect 27858 19966 28142 20018
rect 28194 19966 28196 20018
rect 27804 19964 28196 19966
rect 27804 19954 27860 19964
rect 28140 19954 28196 19964
rect 28364 20020 28420 20078
rect 28476 20132 28644 20188
rect 29708 20132 29764 20142
rect 28476 20130 28532 20132
rect 28476 20078 28478 20130
rect 28530 20078 28532 20130
rect 28476 20066 28532 20078
rect 29708 20038 29764 20076
rect 28364 19954 28420 19964
rect 29372 20020 29428 20030
rect 27580 19908 27636 19918
rect 27580 19906 27748 19908
rect 27580 19854 27582 19906
rect 27634 19854 27748 19906
rect 27580 19852 27748 19854
rect 27580 19842 27636 19852
rect 27692 18564 27748 19852
rect 27916 19234 27972 19246
rect 27916 19182 27918 19234
rect 27970 19182 27972 19234
rect 27916 19012 27972 19182
rect 27916 18946 27972 18956
rect 28140 19010 28196 19022
rect 28140 18958 28142 19010
rect 28194 18958 28196 19010
rect 27804 18564 27860 18574
rect 27692 18562 27860 18564
rect 27692 18510 27806 18562
rect 27858 18510 27860 18562
rect 27692 18508 27860 18510
rect 27804 18498 27860 18508
rect 27020 18452 27076 18462
rect 26572 18450 27412 18452
rect 26572 18398 27022 18450
rect 27074 18398 27412 18450
rect 26572 18396 27412 18398
rect 26460 18050 26516 18060
rect 26684 18338 26740 18396
rect 27020 18386 27076 18396
rect 26684 18286 26686 18338
rect 26738 18286 26740 18338
rect 21532 14756 21588 14766
rect 21532 14662 21588 14700
rect 21756 14754 21812 15092
rect 21756 14702 21758 14754
rect 21810 14702 21812 14754
rect 21756 14690 21812 14702
rect 21420 14644 21476 14654
rect 21420 14550 21476 14588
rect 20412 14478 20414 14530
rect 20466 14478 20468 14530
rect 20412 14466 20468 14478
rect 21868 14418 21924 14430
rect 21868 14366 21870 14418
rect 21922 14366 21924 14418
rect 20748 14308 20804 14318
rect 20748 14306 21028 14308
rect 20748 14254 20750 14306
rect 20802 14254 21028 14306
rect 20748 14252 21028 14254
rect 20748 14242 20804 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19628 13806 19630 13858
rect 19682 13806 19684 13858
rect 19628 13794 19684 13806
rect 20412 13746 20468 13758
rect 20412 13694 20414 13746
rect 20466 13694 20468 13746
rect 20412 13636 20468 13694
rect 20860 13636 20916 13646
rect 18060 13570 18116 13580
rect 20300 13634 20916 13636
rect 20300 13582 20862 13634
rect 20914 13582 20916 13634
rect 20300 13580 20916 13582
rect 17500 13074 17892 13076
rect 17500 13022 17502 13074
rect 17554 13022 17892 13074
rect 17500 13020 17892 13022
rect 18060 13412 18116 13422
rect 18060 13074 18116 13356
rect 18060 13022 18062 13074
rect 18114 13022 18116 13074
rect 17500 11788 17556 13020
rect 18060 13010 18116 13022
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 20300 12178 20356 13580
rect 20860 13412 20916 13580
rect 20860 13346 20916 13356
rect 20972 12290 21028 14252
rect 21868 14084 21924 14366
rect 21868 14028 22372 14084
rect 22316 13860 22372 14028
rect 22428 13860 22484 13870
rect 22316 13858 22484 13860
rect 22316 13806 22430 13858
rect 22482 13806 22484 13858
rect 22316 13804 22484 13806
rect 22428 13794 22484 13804
rect 21756 13746 21812 13758
rect 21756 13694 21758 13746
rect 21810 13694 21812 13746
rect 21756 13412 21812 13694
rect 21756 13346 21812 13356
rect 20972 12238 20974 12290
rect 21026 12238 21028 12290
rect 20972 12226 21028 12238
rect 20300 12126 20302 12178
rect 20354 12126 20356 12178
rect 20300 12114 20356 12126
rect 23100 12066 23156 15092
rect 23548 15036 23996 15092
rect 23548 13412 23604 15036
rect 23996 15026 24052 15036
rect 24332 15092 24948 15148
rect 25340 17668 25396 17678
rect 25340 15092 25396 17612
rect 26684 17668 26740 18286
rect 26684 17602 26740 17612
rect 26124 17556 26180 17566
rect 26124 17462 26180 17500
rect 26908 17556 26964 17566
rect 26908 16996 26964 17500
rect 26908 16210 26964 16940
rect 26908 16158 26910 16210
rect 26962 16158 26964 16210
rect 26908 16146 26964 16158
rect 27356 17444 27412 18396
rect 28140 18340 28196 18958
rect 28140 18274 28196 18284
rect 28252 19012 28308 19022
rect 28252 18452 28308 18956
rect 29372 18676 29428 19964
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 37436 19348 37492 21420
rect 37884 21410 37940 21420
rect 39900 21474 39956 21486
rect 39900 21422 39902 21474
rect 39954 21422 39956 21474
rect 39900 20916 39956 21422
rect 39900 20850 39956 20860
rect 40012 20914 40068 20926
rect 40012 20862 40014 20914
rect 40066 20862 40068 20914
rect 37884 20802 37940 20814
rect 37884 20750 37886 20802
rect 37938 20750 37940 20802
rect 37660 20020 37716 20030
rect 37660 19926 37716 19964
rect 37436 19282 37492 19292
rect 37660 19236 37716 19246
rect 37660 19142 37716 19180
rect 29372 18610 29428 18620
rect 29932 18676 29988 18686
rect 28252 17778 28308 18396
rect 29932 18338 29988 18620
rect 37884 18676 37940 20750
rect 40012 20244 40068 20862
rect 40012 20178 40068 20188
rect 40012 19794 40068 19806
rect 40012 19742 40014 19794
rect 40066 19742 40068 19794
rect 40012 19572 40068 19742
rect 40012 19506 40068 19516
rect 40012 19346 40068 19358
rect 40012 19294 40014 19346
rect 40066 19294 40068 19346
rect 40012 18900 40068 19294
rect 40012 18834 40068 18844
rect 37884 18610 37940 18620
rect 37660 18452 37716 18462
rect 37660 18358 37716 18396
rect 29932 18286 29934 18338
rect 29986 18286 29988 18338
rect 29932 18274 29988 18286
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 28252 17726 28254 17778
rect 28306 17726 28308 17778
rect 28252 17714 28308 17726
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 37660 17668 37716 17678
rect 37660 17574 37716 17612
rect 27356 16210 27412 17388
rect 29260 17444 29316 17454
rect 29260 17350 29316 17388
rect 40012 16884 40068 17726
rect 40012 16818 40068 16828
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 27356 16158 27358 16210
rect 27410 16158 27412 16210
rect 27356 16146 27412 16158
rect 23996 14756 24052 14766
rect 23996 14662 24052 14700
rect 24332 14754 24388 15092
rect 24332 14702 24334 14754
rect 24386 14702 24388 14754
rect 24332 14690 24388 14702
rect 24108 14306 24164 14318
rect 24108 14254 24110 14306
rect 24162 14254 24164 14306
rect 24108 13636 24164 14254
rect 25340 13970 25396 15036
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 25340 13918 25342 13970
rect 25394 13918 25396 13970
rect 25340 13906 25396 13918
rect 24556 13636 24612 13646
rect 24108 13634 24612 13636
rect 24108 13582 24558 13634
rect 24610 13582 24612 13634
rect 24108 13580 24612 13582
rect 23548 12402 23604 13356
rect 23548 12350 23550 12402
rect 23602 12350 23604 12402
rect 23548 12338 23604 12350
rect 23100 12014 23102 12066
rect 23154 12014 23156 12066
rect 23100 11844 23156 12014
rect 23100 11788 23604 11844
rect 17500 11732 17668 11788
rect 17500 4340 17556 4350
rect 17388 4284 17500 4340
rect 17500 4274 17556 4284
rect 17500 3668 17556 3678
rect 17500 800 17556 3612
rect 17612 3554 17668 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19740 4340 19796 4350
rect 19740 4246 19796 4284
rect 19516 4116 19572 4126
rect 18620 3668 18676 3678
rect 18620 3574 18676 3612
rect 17612 3502 17614 3554
rect 17666 3502 17668 3554
rect 17612 3490 17668 3502
rect 19516 800 19572 4060
rect 20748 4116 20804 4126
rect 20748 4022 20804 4060
rect 23548 3554 23604 11788
rect 23548 3502 23550 3554
rect 23602 3502 23604 3554
rect 23548 3490 23604 3502
rect 24220 3668 24276 3678
rect 22204 3442 22260 3454
rect 22204 3390 22206 3442
rect 22258 3390 22260 3442
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 22204 800 22260 3390
rect 24220 800 24276 3612
rect 24556 3554 24612 13580
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 15456 0 15568 800
rect 17472 0 17584 800
rect 19488 0 19600 800
rect 22176 0 22288 800
rect 24192 0 24304 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 16828 38220 16884 38276
rect 18060 38274 18116 38276
rect 18060 38222 18062 38274
rect 18062 38222 18114 38274
rect 18114 38222 18116 38274
rect 18060 38220 18116 38222
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 18844 37436 18900 37492
rect 19852 37490 19908 37492
rect 19852 37438 19854 37490
rect 19854 37438 19906 37490
rect 19906 37438 19908 37490
rect 19852 37436 19908 37438
rect 25564 38556 25620 38612
rect 26796 38556 26852 38612
rect 24220 38220 24276 38276
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 21532 37436 21588 37492
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 14364 28588 14420 28644
rect 15148 28642 15204 28644
rect 15148 28590 15150 28642
rect 15150 28590 15202 28642
rect 15202 28590 15204 28642
rect 15148 28588 15204 28590
rect 4172 27580 4228 27636
rect 1932 25564 1988 25620
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 13692 26460 13748 26516
rect 14588 26460 14644 26516
rect 4284 26290 4340 26292
rect 4284 26238 4286 26290
rect 4286 26238 4338 26290
rect 4338 26238 4340 26290
rect 4284 26236 4340 26238
rect 11788 26236 11844 26292
rect 15148 26460 15204 26516
rect 14700 26236 14756 26292
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 13916 25676 13972 25732
rect 14812 25506 14868 25508
rect 14812 25454 14814 25506
rect 14814 25454 14866 25506
rect 14866 25454 14868 25506
rect 14812 25452 14868 25454
rect 12572 24444 12628 24500
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 14812 23884 14868 23940
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4172 21420 4228 21476
rect 12684 22988 12740 23044
rect 14700 22540 14756 22596
rect 14924 23548 14980 23604
rect 14700 21756 14756 21812
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 9996 21196 10052 21252
rect 9996 20914 10052 20916
rect 9996 20862 9998 20914
rect 9998 20862 10050 20914
rect 10050 20862 10052 20914
rect 9996 20860 10052 20862
rect 11900 20860 11956 20916
rect 12908 20860 12964 20916
rect 4284 20802 4340 20804
rect 4284 20750 4286 20802
rect 4286 20750 4338 20802
rect 4338 20750 4340 20802
rect 4284 20748 4340 20750
rect 13580 20914 13636 20916
rect 13580 20862 13582 20914
rect 13582 20862 13634 20914
rect 13634 20862 13636 20914
rect 13580 20860 13636 20862
rect 1932 20188 1988 20244
rect 12236 20018 12292 20020
rect 12236 19966 12238 20018
rect 12238 19966 12290 20018
rect 12290 19966 12292 20018
rect 12236 19964 12292 19966
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 11676 18562 11732 18564
rect 11676 18510 11678 18562
rect 11678 18510 11730 18562
rect 11730 18510 11732 18562
rect 11676 18508 11732 18510
rect 10108 18284 10164 18340
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 11004 18284 11060 18340
rect 10780 18172 10836 18228
rect 12908 17778 12964 17780
rect 12908 17726 12910 17778
rect 12910 17726 12962 17778
rect 12962 17726 12964 17778
rect 12908 17724 12964 17726
rect 15820 25730 15876 25732
rect 15820 25678 15822 25730
rect 15822 25678 15874 25730
rect 15874 25678 15876 25730
rect 15820 25676 15876 25678
rect 15260 25506 15316 25508
rect 15260 25454 15262 25506
rect 15262 25454 15314 25506
rect 15314 25454 15316 25506
rect 15260 25452 15316 25454
rect 15484 25116 15540 25172
rect 15708 24892 15764 24948
rect 15036 22146 15092 22148
rect 15036 22094 15038 22146
rect 15038 22094 15090 22146
rect 15090 22094 15092 22146
rect 15036 22092 15092 22094
rect 15484 23548 15540 23604
rect 15372 21868 15428 21924
rect 15148 20860 15204 20916
rect 14700 19458 14756 19460
rect 14700 19406 14702 19458
rect 14702 19406 14754 19458
rect 14754 19406 14756 19458
rect 14700 19404 14756 19406
rect 14924 19516 14980 19572
rect 15932 23266 15988 23268
rect 15932 23214 15934 23266
rect 15934 23214 15986 23266
rect 15986 23214 15988 23266
rect 15932 23212 15988 23214
rect 16380 26962 16436 26964
rect 16380 26910 16382 26962
rect 16382 26910 16434 26962
rect 16434 26910 16436 26962
rect 16380 26908 16436 26910
rect 17276 26460 17332 26516
rect 17052 26348 17108 26404
rect 17500 26908 17556 26964
rect 17500 26460 17556 26516
rect 17948 27020 18004 27076
rect 17836 26348 17892 26404
rect 18060 26962 18116 26964
rect 18060 26910 18062 26962
rect 18062 26910 18114 26962
rect 18114 26910 18116 26962
rect 18060 26908 18116 26910
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 18732 27692 18788 27748
rect 18844 27244 18900 27300
rect 18732 26908 18788 26964
rect 18172 26514 18228 26516
rect 18172 26462 18174 26514
rect 18174 26462 18226 26514
rect 18226 26462 18228 26514
rect 18172 26460 18228 26462
rect 18508 26460 18564 26516
rect 17388 25116 17444 25172
rect 16492 24946 16548 24948
rect 16492 24894 16494 24946
rect 16494 24894 16546 24946
rect 16546 24894 16548 24946
rect 16492 24892 16548 24894
rect 16716 24722 16772 24724
rect 16716 24670 16718 24722
rect 16718 24670 16770 24722
rect 16770 24670 16772 24722
rect 16716 24668 16772 24670
rect 17724 24668 17780 24724
rect 16156 23938 16212 23940
rect 16156 23886 16158 23938
rect 16158 23886 16210 23938
rect 16210 23886 16212 23938
rect 16156 23884 16212 23886
rect 17612 23884 17668 23940
rect 16604 23436 16660 23492
rect 15708 23042 15764 23044
rect 15708 22990 15710 23042
rect 15710 22990 15762 23042
rect 15762 22990 15764 23042
rect 15708 22988 15764 22990
rect 15596 22204 15652 22260
rect 15932 22540 15988 22596
rect 15708 21980 15764 22036
rect 16828 23154 16884 23156
rect 16828 23102 16830 23154
rect 16830 23102 16882 23154
rect 16882 23102 16884 23154
rect 16828 23100 16884 23102
rect 16380 22428 16436 22484
rect 16044 22258 16100 22260
rect 16044 22206 16046 22258
rect 16046 22206 16098 22258
rect 16098 22206 16100 22258
rect 16044 22204 16100 22206
rect 15932 21868 15988 21924
rect 17388 23266 17444 23268
rect 17388 23214 17390 23266
rect 17390 23214 17442 23266
rect 17442 23214 17444 23266
rect 17388 23212 17444 23214
rect 17612 23100 17668 23156
rect 17612 22540 17668 22596
rect 17948 24498 18004 24500
rect 17948 24446 17950 24498
rect 17950 24446 18002 24498
rect 18002 24446 18004 24498
rect 17948 24444 18004 24446
rect 19180 28476 19236 28532
rect 21644 28476 21700 28532
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 22764 37490 22820 37492
rect 22764 37438 22766 37490
rect 22766 37438 22818 37490
rect 22818 37438 22820 37490
rect 22764 37436 22820 37438
rect 20300 27746 20356 27748
rect 20300 27694 20302 27746
rect 20302 27694 20354 27746
rect 20354 27694 20356 27746
rect 20300 27692 20356 27694
rect 19964 27298 20020 27300
rect 19964 27246 19966 27298
rect 19966 27246 20018 27298
rect 20018 27246 20020 27298
rect 19964 27244 20020 27246
rect 18844 26348 18900 26404
rect 19068 26460 19124 26516
rect 19516 27074 19572 27076
rect 19516 27022 19518 27074
rect 19518 27022 19570 27074
rect 19570 27022 19572 27074
rect 19516 27020 19572 27022
rect 22540 28476 22596 28532
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 22764 27692 22820 27748
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19404 25452 19460 25508
rect 18620 24834 18676 24836
rect 18620 24782 18622 24834
rect 18622 24782 18674 24834
rect 18674 24782 18676 24834
rect 18620 24780 18676 24782
rect 18844 24780 18900 24836
rect 18396 24668 18452 24724
rect 18172 23436 18228 23492
rect 17052 22428 17108 22484
rect 17948 23212 18004 23268
rect 18284 23772 18340 23828
rect 16380 22092 16436 22148
rect 16604 21980 16660 22036
rect 16716 21868 16772 21924
rect 18060 22540 18116 22596
rect 17276 21980 17332 22036
rect 16268 21532 16324 21588
rect 14252 18338 14308 18340
rect 14252 18286 14254 18338
rect 14254 18286 14306 18338
rect 14306 18286 14308 18338
rect 14252 18284 14308 18286
rect 13580 16828 13636 16884
rect 13804 16940 13860 16996
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 1932 15484 1988 15540
rect 4284 15260 4340 15316
rect 11676 15820 11732 15876
rect 14476 17724 14532 17780
rect 14812 18060 14868 18116
rect 15820 19458 15876 19460
rect 15820 19406 15822 19458
rect 15822 19406 15874 19458
rect 15874 19406 15876 19458
rect 15820 19404 15876 19406
rect 16044 19516 16100 19572
rect 16156 19346 16212 19348
rect 16156 19294 16158 19346
rect 16158 19294 16210 19346
rect 16210 19294 16212 19346
rect 16156 19292 16212 19294
rect 16044 19180 16100 19236
rect 15820 18956 15876 19012
rect 15820 18674 15876 18676
rect 15820 18622 15822 18674
rect 15822 18622 15874 18674
rect 15874 18622 15876 18674
rect 15820 18620 15876 18622
rect 16044 18674 16100 18676
rect 16044 18622 16046 18674
rect 16046 18622 16098 18674
rect 16098 18622 16100 18674
rect 16044 18620 16100 18622
rect 16604 19346 16660 19348
rect 16604 19294 16606 19346
rect 16606 19294 16658 19346
rect 16658 19294 16660 19346
rect 16604 19292 16660 19294
rect 16492 19010 16548 19012
rect 16492 18958 16494 19010
rect 16494 18958 16546 19010
rect 16546 18958 16548 19010
rect 16492 18956 16548 18958
rect 16940 18620 16996 18676
rect 15708 18060 15764 18116
rect 15596 17836 15652 17892
rect 14252 16828 14308 16884
rect 14812 16828 14868 16884
rect 11676 15260 11732 15316
rect 15036 16156 15092 16212
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 13132 14252 13188 14308
rect 12460 13746 12516 13748
rect 12460 13694 12462 13746
rect 12462 13694 12514 13746
rect 12514 13694 12516 13746
rect 12460 13692 12516 13694
rect 15484 17164 15540 17220
rect 15484 16994 15540 16996
rect 15484 16942 15486 16994
rect 15486 16942 15538 16994
rect 15538 16942 15540 16994
rect 15484 16940 15540 16942
rect 15148 16156 15204 16212
rect 15260 15874 15316 15876
rect 15260 15822 15262 15874
rect 15262 15822 15314 15874
rect 15314 15822 15316 15874
rect 15260 15820 15316 15822
rect 15484 15820 15540 15876
rect 15148 15426 15204 15428
rect 15148 15374 15150 15426
rect 15150 15374 15202 15426
rect 15202 15374 15204 15426
rect 15148 15372 15204 15374
rect 14812 14306 14868 14308
rect 14812 14254 14814 14306
rect 14814 14254 14866 14306
rect 14866 14254 14868 14306
rect 14812 14252 14868 14254
rect 14588 13692 14644 13748
rect 16156 17724 16212 17780
rect 17500 21698 17556 21700
rect 17500 21646 17502 21698
rect 17502 21646 17554 21698
rect 17554 21646 17556 21698
rect 17500 21644 17556 21646
rect 17836 21586 17892 21588
rect 17836 21534 17838 21586
rect 17838 21534 17890 21586
rect 17890 21534 17892 21586
rect 17836 21532 17892 21534
rect 18284 22092 18340 22148
rect 18172 20524 18228 20580
rect 18620 22540 18676 22596
rect 18396 21644 18452 21700
rect 18284 19852 18340 19908
rect 18620 21586 18676 21588
rect 18620 21534 18622 21586
rect 18622 21534 18674 21586
rect 18674 21534 18676 21586
rect 18620 21532 18676 21534
rect 18620 19234 18676 19236
rect 18620 19182 18622 19234
rect 18622 19182 18674 19234
rect 18674 19182 18676 19234
rect 18620 19180 18676 19182
rect 17052 17778 17108 17780
rect 17052 17726 17054 17778
rect 17054 17726 17106 17778
rect 17106 17726 17108 17778
rect 17052 17724 17108 17726
rect 16268 17500 16324 17556
rect 16492 17612 16548 17668
rect 17164 17666 17220 17668
rect 17164 17614 17166 17666
rect 17166 17614 17218 17666
rect 17218 17614 17220 17666
rect 17164 17612 17220 17614
rect 15932 16994 15988 16996
rect 15932 16942 15934 16994
rect 15934 16942 15986 16994
rect 15986 16942 15988 16994
rect 15932 16940 15988 16942
rect 16380 16156 16436 16212
rect 17500 18396 17556 18452
rect 17388 17500 17444 17556
rect 18508 18450 18564 18452
rect 18508 18398 18510 18450
rect 18510 18398 18562 18450
rect 18562 18398 18564 18450
rect 18508 18396 18564 18398
rect 18060 17890 18116 17892
rect 18060 17838 18062 17890
rect 18062 17838 18114 17890
rect 18114 17838 18116 17890
rect 18060 17836 18116 17838
rect 18396 18226 18452 18228
rect 18396 18174 18398 18226
rect 18398 18174 18450 18226
rect 18450 18174 18452 18226
rect 18396 18172 18452 18174
rect 18620 17724 18676 17780
rect 18284 17666 18340 17668
rect 18284 17614 18286 17666
rect 18286 17614 18338 17666
rect 18338 17614 18340 17666
rect 18284 17612 18340 17614
rect 18508 17500 18564 17556
rect 17948 17052 18004 17108
rect 17500 16940 17556 16996
rect 16492 15874 16548 15876
rect 16492 15822 16494 15874
rect 16494 15822 16546 15874
rect 16546 15822 16548 15874
rect 16492 15820 16548 15822
rect 17724 15426 17780 15428
rect 17724 15374 17726 15426
rect 17726 15374 17778 15426
rect 17778 15374 17780 15426
rect 17724 15372 17780 15374
rect 17052 14642 17108 14644
rect 17052 14590 17054 14642
rect 17054 14590 17106 14642
rect 17106 14590 17108 14642
rect 17052 14588 17108 14590
rect 15596 14476 15652 14532
rect 16828 14530 16884 14532
rect 16828 14478 16830 14530
rect 16830 14478 16882 14530
rect 16882 14478 16884 14530
rect 16828 14476 16884 14478
rect 16492 14364 16548 14420
rect 16268 14252 16324 14308
rect 17164 14530 17220 14532
rect 17164 14478 17166 14530
rect 17166 14478 17218 14530
rect 17218 14478 17220 14530
rect 17164 14476 17220 14478
rect 18956 22930 19012 22932
rect 18956 22878 18958 22930
rect 18958 22878 19010 22930
rect 19010 22878 19012 22930
rect 18956 22876 19012 22878
rect 18956 21586 19012 21588
rect 18956 21534 18958 21586
rect 18958 21534 19010 21586
rect 19010 21534 19012 21586
rect 18956 21532 19012 21534
rect 21868 26850 21924 26852
rect 21868 26798 21870 26850
rect 21870 26798 21922 26850
rect 21922 26798 21924 26850
rect 21868 26796 21924 26798
rect 22204 26962 22260 26964
rect 22204 26910 22206 26962
rect 22206 26910 22258 26962
rect 22258 26910 22260 26962
rect 22204 26908 22260 26910
rect 22428 26236 22484 26292
rect 21308 25506 21364 25508
rect 21308 25454 21310 25506
rect 21310 25454 21362 25506
rect 21362 25454 21364 25506
rect 21308 25452 21364 25454
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 21420 24332 21476 24388
rect 21308 23826 21364 23828
rect 21308 23774 21310 23826
rect 21310 23774 21362 23826
rect 21362 23774 21364 23826
rect 21308 23772 21364 23774
rect 21644 23772 21700 23828
rect 21420 23714 21476 23716
rect 21420 23662 21422 23714
rect 21422 23662 21474 23714
rect 21474 23662 21476 23714
rect 21420 23660 21476 23662
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19516 23324 19572 23380
rect 21084 23378 21140 23380
rect 21084 23326 21086 23378
rect 21086 23326 21138 23378
rect 21138 23326 21140 23378
rect 21084 23324 21140 23326
rect 19068 19740 19124 19796
rect 20412 23266 20468 23268
rect 20412 23214 20414 23266
rect 20414 23214 20466 23266
rect 20466 23214 20468 23266
rect 20412 23212 20468 23214
rect 19740 23100 19796 23156
rect 19964 22652 20020 22708
rect 21980 24892 22036 24948
rect 22316 24332 22372 24388
rect 22204 23324 22260 23380
rect 20076 22540 20132 22596
rect 20412 22876 20468 22932
rect 19516 21420 19572 21476
rect 19292 20188 19348 20244
rect 19180 19180 19236 19236
rect 19292 19852 19348 19908
rect 19292 19628 19348 19684
rect 20860 22652 20916 22708
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20076 20802 20132 20804
rect 20076 20750 20078 20802
rect 20078 20750 20130 20802
rect 20130 20750 20132 20802
rect 20076 20748 20132 20750
rect 20188 20524 20244 20580
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20076 19852 20132 19908
rect 19628 19346 19684 19348
rect 19628 19294 19630 19346
rect 19630 19294 19682 19346
rect 19682 19294 19684 19346
rect 19628 19292 19684 19294
rect 19852 19516 19908 19572
rect 22092 23266 22148 23268
rect 22092 23214 22094 23266
rect 22094 23214 22146 23266
rect 22146 23214 22148 23266
rect 22092 23212 22148 23214
rect 21644 22540 21700 22596
rect 21756 23100 21812 23156
rect 20748 21868 20804 21924
rect 20524 20076 20580 20132
rect 20300 20018 20356 20020
rect 20300 19966 20302 20018
rect 20302 19966 20354 20018
rect 20354 19966 20356 20018
rect 20300 19964 20356 19966
rect 20412 19740 20468 19796
rect 20636 19852 20692 19908
rect 18956 18172 19012 18228
rect 19180 18396 19236 18452
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19628 18562 19684 18564
rect 19628 18510 19630 18562
rect 19630 18510 19682 18562
rect 19682 18510 19684 18562
rect 19628 18508 19684 18510
rect 20972 19516 21028 19572
rect 19516 17666 19572 17668
rect 19516 17614 19518 17666
rect 19518 17614 19570 17666
rect 19570 17614 19572 17666
rect 19516 17612 19572 17614
rect 19180 17500 19236 17556
rect 20076 17554 20132 17556
rect 20076 17502 20078 17554
rect 20078 17502 20130 17554
rect 20130 17502 20132 17554
rect 20076 17500 20132 17502
rect 19516 16940 19572 16996
rect 19628 17388 19684 17444
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19404 16828 19460 16884
rect 20300 17500 20356 17556
rect 19964 16994 20020 16996
rect 19964 16942 19966 16994
rect 19966 16942 20018 16994
rect 20018 16942 20020 16994
rect 19964 16940 20020 16942
rect 19180 15932 19236 15988
rect 18396 14754 18452 14756
rect 18396 14702 18398 14754
rect 18398 14702 18450 14754
rect 18450 14702 18452 14754
rect 18396 14700 18452 14702
rect 19628 15986 19684 15988
rect 19628 15934 19630 15986
rect 19630 15934 19682 15986
rect 19682 15934 19684 15986
rect 19628 15932 19684 15934
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 18956 14530 19012 14532
rect 18956 14478 18958 14530
rect 18958 14478 19010 14530
rect 19010 14478 19012 14530
rect 18956 14476 19012 14478
rect 17388 14306 17444 14308
rect 17388 14254 17390 14306
rect 17390 14254 17442 14306
rect 17442 14254 17444 14306
rect 17388 14252 17444 14254
rect 14700 13356 14756 13412
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 15708 13468 15764 13524
rect 17500 13634 17556 13636
rect 17500 13582 17502 13634
rect 17502 13582 17554 13634
rect 17554 13582 17556 13634
rect 17500 13580 17556 13582
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 15484 5180 15540 5236
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 16716 5234 16772 5236
rect 16716 5182 16718 5234
rect 16718 5182 16770 5234
rect 16770 5182 16772 5234
rect 16716 5180 16772 5182
rect 19740 14754 19796 14756
rect 19740 14702 19742 14754
rect 19742 14702 19794 14754
rect 19794 14702 19796 14754
rect 19740 14700 19796 14702
rect 20860 18060 20916 18116
rect 21532 22092 21588 22148
rect 21868 22204 21924 22260
rect 22092 21868 22148 21924
rect 21420 20188 21476 20244
rect 21532 20130 21588 20132
rect 21532 20078 21534 20130
rect 21534 20078 21586 20130
rect 21586 20078 21588 20130
rect 21532 20076 21588 20078
rect 21756 19794 21812 19796
rect 21756 19742 21758 19794
rect 21758 19742 21810 19794
rect 21810 19742 21812 19794
rect 21756 19740 21812 19742
rect 21532 19628 21588 19684
rect 21308 18172 21364 18228
rect 21532 18620 21588 18676
rect 22092 20076 22148 20132
rect 22092 19906 22148 19908
rect 22092 19854 22094 19906
rect 22094 19854 22146 19906
rect 22146 19854 22148 19906
rect 22092 19852 22148 19854
rect 22092 19628 22148 19684
rect 21980 18620 22036 18676
rect 22204 19404 22260 19460
rect 23436 26796 23492 26852
rect 25228 27692 25284 27748
rect 25452 26908 25508 26964
rect 24444 26236 24500 26292
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 25788 27692 25844 27748
rect 25452 25900 25508 25956
rect 24668 25506 24724 25508
rect 24668 25454 24670 25506
rect 24670 25454 24722 25506
rect 24722 25454 24724 25506
rect 24668 25452 24724 25454
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 25900 25900 25956 25956
rect 25676 25452 25732 25508
rect 26124 25394 26180 25396
rect 26124 25342 26126 25394
rect 26126 25342 26178 25394
rect 26178 25342 26180 25394
rect 26124 25340 26180 25342
rect 24892 25228 24948 25284
rect 23660 24892 23716 24948
rect 23660 23660 23716 23716
rect 23212 22258 23268 22260
rect 23212 22206 23214 22258
rect 23214 22206 23266 22258
rect 23266 22206 23268 22258
rect 23212 22204 23268 22206
rect 22540 22146 22596 22148
rect 22540 22094 22542 22146
rect 22542 22094 22594 22146
rect 22594 22094 22596 22146
rect 22540 22092 22596 22094
rect 22652 20802 22708 20804
rect 22652 20750 22654 20802
rect 22654 20750 22706 20802
rect 22706 20750 22708 20802
rect 22652 20748 22708 20750
rect 22428 19906 22484 19908
rect 22428 19854 22430 19906
rect 22430 19854 22482 19906
rect 22482 19854 22484 19906
rect 22428 19852 22484 19854
rect 22764 20018 22820 20020
rect 22764 19966 22766 20018
rect 22766 19966 22818 20018
rect 22818 19966 22820 20018
rect 22764 19964 22820 19966
rect 23436 20130 23492 20132
rect 23436 20078 23438 20130
rect 23438 20078 23490 20130
rect 23490 20078 23492 20130
rect 23436 20076 23492 20078
rect 22876 19852 22932 19908
rect 22540 19404 22596 19460
rect 22428 19346 22484 19348
rect 22428 19294 22430 19346
rect 22430 19294 22482 19346
rect 22482 19294 22484 19346
rect 22428 19292 22484 19294
rect 21196 17724 21252 17780
rect 20524 17554 20580 17556
rect 20524 17502 20526 17554
rect 20526 17502 20578 17554
rect 20578 17502 20580 17554
rect 20524 17500 20580 17502
rect 21644 17554 21700 17556
rect 21644 17502 21646 17554
rect 21646 17502 21698 17554
rect 21698 17502 21700 17554
rect 21644 17500 21700 17502
rect 20860 17052 20916 17108
rect 20636 16882 20692 16884
rect 20636 16830 20638 16882
rect 20638 16830 20690 16882
rect 20690 16830 20692 16882
rect 20636 16828 20692 16830
rect 21196 17106 21252 17108
rect 21196 17054 21198 17106
rect 21198 17054 21250 17106
rect 21250 17054 21252 17106
rect 21196 17052 21252 17054
rect 21420 16828 21476 16884
rect 20524 16716 20580 16772
rect 20524 15820 20580 15876
rect 21532 16716 21588 16772
rect 21868 17778 21924 17780
rect 21868 17726 21870 17778
rect 21870 17726 21922 17778
rect 21922 17726 21924 17778
rect 21868 17724 21924 17726
rect 21756 15986 21812 15988
rect 21756 15934 21758 15986
rect 21758 15934 21810 15986
rect 21810 15934 21812 15986
rect 21756 15932 21812 15934
rect 22204 18226 22260 18228
rect 22204 18174 22206 18226
rect 22206 18174 22258 18226
rect 22258 18174 22260 18226
rect 22204 18172 22260 18174
rect 23324 18956 23380 19012
rect 23660 23436 23716 23492
rect 23996 24834 24052 24836
rect 23996 24782 23998 24834
rect 23998 24782 24050 24834
rect 24050 24782 24052 24834
rect 23996 24780 24052 24782
rect 24220 24780 24276 24836
rect 23996 23660 24052 23716
rect 24332 24722 24388 24724
rect 24332 24670 24334 24722
rect 24334 24670 24386 24722
rect 24386 24670 24388 24722
rect 24332 24668 24388 24670
rect 24220 23548 24276 23604
rect 24220 23212 24276 23268
rect 24556 22988 24612 23044
rect 24220 22370 24276 22372
rect 24220 22318 24222 22370
rect 24222 22318 24274 22370
rect 24274 22318 24276 22370
rect 24220 22316 24276 22318
rect 25564 25282 25620 25284
rect 25564 25230 25566 25282
rect 25566 25230 25618 25282
rect 25618 25230 25620 25282
rect 25564 25228 25620 25230
rect 25676 24668 25732 24724
rect 25676 24050 25732 24052
rect 25676 23998 25678 24050
rect 25678 23998 25730 24050
rect 25730 23998 25732 24050
rect 25676 23996 25732 23998
rect 27468 26124 27524 26180
rect 27244 25394 27300 25396
rect 27244 25342 27246 25394
rect 27246 25342 27298 25394
rect 27298 25342 27300 25394
rect 27244 25340 27300 25342
rect 28476 26178 28532 26180
rect 28476 26126 28478 26178
rect 28478 26126 28530 26178
rect 28530 26126 28532 26178
rect 28476 26124 28532 26126
rect 26908 24834 26964 24836
rect 26908 24782 26910 24834
rect 26910 24782 26962 24834
rect 26962 24782 26964 24834
rect 26908 24780 26964 24782
rect 26460 24668 26516 24724
rect 26796 24668 26852 24724
rect 25340 22988 25396 23044
rect 23884 22204 23940 22260
rect 23996 19346 24052 19348
rect 23996 19294 23998 19346
rect 23998 19294 24050 19346
rect 24050 19294 24052 19346
rect 23996 19292 24052 19294
rect 22764 17948 22820 18004
rect 22876 17890 22932 17892
rect 22876 17838 22878 17890
rect 22878 17838 22930 17890
rect 22930 17838 22932 17890
rect 22876 17836 22932 17838
rect 23324 18284 23380 18340
rect 23996 18284 24052 18340
rect 23884 18172 23940 18228
rect 23100 17836 23156 17892
rect 22092 17666 22148 17668
rect 22092 17614 22094 17666
rect 22094 17614 22146 17666
rect 22146 17614 22148 17666
rect 22092 17612 22148 17614
rect 21980 17388 22036 17444
rect 22540 17500 22596 17556
rect 22764 16994 22820 16996
rect 22764 16942 22766 16994
rect 22766 16942 22818 16994
rect 22818 16942 22820 16994
rect 22764 16940 22820 16942
rect 22876 16828 22932 16884
rect 23436 17948 23492 18004
rect 23212 17442 23268 17444
rect 23212 17390 23214 17442
rect 23214 17390 23266 17442
rect 23266 17390 23268 17442
rect 23212 17388 23268 17390
rect 23772 17388 23828 17444
rect 23436 17052 23492 17108
rect 23772 17052 23828 17108
rect 23548 16882 23604 16884
rect 23548 16830 23550 16882
rect 23550 16830 23602 16882
rect 23602 16830 23604 16882
rect 23548 16828 23604 16830
rect 24332 18284 24388 18340
rect 24220 17554 24276 17556
rect 24220 17502 24222 17554
rect 24222 17502 24274 17554
rect 24274 17502 24276 17554
rect 24220 17500 24276 17502
rect 24332 17388 24388 17444
rect 25228 22540 25284 22596
rect 25228 22204 25284 22260
rect 25452 22316 25508 22372
rect 26124 22316 26180 22372
rect 25228 19852 25284 19908
rect 26124 20076 26180 20132
rect 26460 23378 26516 23380
rect 26460 23326 26462 23378
rect 26462 23326 26514 23378
rect 26514 23326 26516 23378
rect 26460 23324 26516 23326
rect 27356 24722 27412 24724
rect 27356 24670 27358 24722
rect 27358 24670 27410 24722
rect 27410 24670 27412 24722
rect 27356 24668 27412 24670
rect 40012 26236 40068 26292
rect 37660 26124 37716 26180
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 30940 24834 30996 24836
rect 30940 24782 30942 24834
rect 30942 24782 30994 24834
rect 30994 24782 30996 24834
rect 30940 24780 30996 24782
rect 28924 24668 28980 24724
rect 30716 24722 30772 24724
rect 30716 24670 30718 24722
rect 30718 24670 30770 24722
rect 30770 24670 30772 24722
rect 30716 24668 30772 24670
rect 40012 24892 40068 24948
rect 37436 24668 37492 24724
rect 37660 24722 37716 24724
rect 37660 24670 37662 24722
rect 37662 24670 37714 24722
rect 37714 24670 37716 24722
rect 37660 24668 37716 24670
rect 28140 23938 28196 23940
rect 28140 23886 28142 23938
rect 28142 23886 28194 23938
rect 28194 23886 28196 23938
rect 28140 23884 28196 23886
rect 28028 23826 28084 23828
rect 28028 23774 28030 23826
rect 28030 23774 28082 23826
rect 28082 23774 28084 23826
rect 28028 23772 28084 23774
rect 27580 23660 27636 23716
rect 27132 23212 27188 23268
rect 27804 23266 27860 23268
rect 27804 23214 27806 23266
rect 27806 23214 27858 23266
rect 27858 23214 27860 23266
rect 27804 23212 27860 23214
rect 26684 22258 26740 22260
rect 26684 22206 26686 22258
rect 26686 22206 26738 22258
rect 26738 22206 26740 22258
rect 26684 22204 26740 22206
rect 29260 23884 29316 23940
rect 29596 23826 29652 23828
rect 29596 23774 29598 23826
rect 29598 23774 29650 23826
rect 29650 23774 29652 23826
rect 29596 23772 29652 23774
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 40012 24220 40068 24276
rect 37660 23938 37716 23940
rect 37660 23886 37662 23938
rect 37662 23886 37714 23938
rect 37714 23886 37716 23938
rect 37660 23884 37716 23886
rect 30268 23772 30324 23828
rect 29036 23324 29092 23380
rect 28588 22988 28644 23044
rect 27020 22316 27076 22372
rect 28364 22370 28420 22372
rect 28364 22318 28366 22370
rect 28366 22318 28418 22370
rect 28418 22318 28420 22370
rect 28364 22316 28420 22318
rect 28140 22258 28196 22260
rect 28140 22206 28142 22258
rect 28142 22206 28194 22258
rect 28194 22206 28196 22258
rect 28140 22204 28196 22206
rect 29036 22204 29092 22260
rect 28476 20860 28532 20916
rect 28588 20748 28644 20804
rect 28364 20578 28420 20580
rect 28364 20526 28366 20578
rect 28366 20526 28418 20578
rect 28418 20526 28420 20578
rect 28364 20524 28420 20526
rect 40012 23548 40068 23604
rect 37660 23154 37716 23156
rect 37660 23102 37662 23154
rect 37662 23102 37714 23154
rect 37714 23102 37716 23154
rect 37660 23100 37716 23102
rect 29932 23042 29988 23044
rect 29932 22990 29934 23042
rect 29934 22990 29986 23042
rect 29986 22990 29988 23042
rect 29932 22988 29988 22990
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 29372 22316 29428 22372
rect 29260 20914 29316 20916
rect 29260 20862 29262 20914
rect 29262 20862 29314 20914
rect 29314 20862 29316 20914
rect 29260 20860 29316 20862
rect 29372 20802 29428 20804
rect 29372 20750 29374 20802
rect 29374 20750 29426 20802
rect 29426 20750 29428 20802
rect 29372 20748 29428 20750
rect 29596 21420 29652 21476
rect 30156 21474 30212 21476
rect 30156 21422 30158 21474
rect 30158 21422 30210 21474
rect 30210 21422 30212 21474
rect 30156 21420 30212 21422
rect 40012 21532 40068 21588
rect 37884 21420 37940 21476
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 26572 19964 26628 20020
rect 26124 19346 26180 19348
rect 26124 19294 26126 19346
rect 26126 19294 26178 19346
rect 26178 19294 26180 19346
rect 26124 19292 26180 19294
rect 25452 18674 25508 18676
rect 25452 18622 25454 18674
rect 25454 18622 25506 18674
rect 25506 18622 25508 18674
rect 25452 18620 25508 18622
rect 25900 18450 25956 18452
rect 25900 18398 25902 18450
rect 25902 18398 25954 18450
rect 25954 18398 25956 18450
rect 25900 18396 25956 18398
rect 25340 18338 25396 18340
rect 25340 18286 25342 18338
rect 25342 18286 25394 18338
rect 25394 18286 25396 18338
rect 25340 18284 25396 18286
rect 26572 19010 26628 19012
rect 26572 18958 26574 19010
rect 26574 18958 26626 19010
rect 26626 18958 26628 19010
rect 26572 18956 26628 18958
rect 27132 20130 27188 20132
rect 27132 20078 27134 20130
rect 27134 20078 27186 20130
rect 27186 20078 27188 20130
rect 27132 20076 27188 20078
rect 27356 20018 27412 20020
rect 27356 19966 27358 20018
rect 27358 19966 27410 20018
rect 27410 19966 27412 20018
rect 27356 19964 27412 19966
rect 29708 20130 29764 20132
rect 29708 20078 29710 20130
rect 29710 20078 29762 20130
rect 29762 20078 29764 20130
rect 29708 20076 29764 20078
rect 28364 19964 28420 20020
rect 29372 20018 29428 20020
rect 29372 19966 29374 20018
rect 29374 19966 29426 20018
rect 29426 19966 29428 20018
rect 29372 19964 29428 19966
rect 27916 18956 27972 19012
rect 26460 18060 26516 18116
rect 21532 14754 21588 14756
rect 21532 14702 21534 14754
rect 21534 14702 21586 14754
rect 21586 14702 21588 14754
rect 21532 14700 21588 14702
rect 21420 14642 21476 14644
rect 21420 14590 21422 14642
rect 21422 14590 21474 14642
rect 21474 14590 21476 14642
rect 21420 14588 21476 14590
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 18060 13580 18116 13636
rect 18060 13356 18116 13412
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 20860 13356 20916 13412
rect 21756 13356 21812 13412
rect 23996 15036 24052 15092
rect 25340 17666 25396 17668
rect 25340 17614 25342 17666
rect 25342 17614 25394 17666
rect 25394 17614 25396 17666
rect 25340 17612 25396 17614
rect 26684 17612 26740 17668
rect 26124 17554 26180 17556
rect 26124 17502 26126 17554
rect 26126 17502 26178 17554
rect 26178 17502 26180 17554
rect 26124 17500 26180 17502
rect 26908 17500 26964 17556
rect 26908 16940 26964 16996
rect 28140 18284 28196 18340
rect 28252 18956 28308 19012
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 39900 20860 39956 20916
rect 37660 20018 37716 20020
rect 37660 19966 37662 20018
rect 37662 19966 37714 20018
rect 37714 19966 37716 20018
rect 37660 19964 37716 19966
rect 37436 19292 37492 19348
rect 37660 19234 37716 19236
rect 37660 19182 37662 19234
rect 37662 19182 37714 19234
rect 37714 19182 37716 19234
rect 37660 19180 37716 19182
rect 29372 18620 29428 18676
rect 29932 18620 29988 18676
rect 28252 18396 28308 18452
rect 40012 20188 40068 20244
rect 40012 19516 40068 19572
rect 40012 18844 40068 18900
rect 37884 18620 37940 18676
rect 37660 18450 37716 18452
rect 37660 18398 37662 18450
rect 37662 18398 37714 18450
rect 37714 18398 37716 18450
rect 37660 18396 37716 18398
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 37660 17666 37716 17668
rect 37660 17614 37662 17666
rect 37662 17614 37714 17666
rect 37714 17614 37716 17666
rect 37660 17612 37716 17614
rect 27356 17388 27412 17444
rect 29260 17442 29316 17444
rect 29260 17390 29262 17442
rect 29262 17390 29314 17442
rect 29314 17390 29316 17442
rect 29260 17388 29316 17390
rect 40012 16828 40068 16884
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 23996 14754 24052 14756
rect 23996 14702 23998 14754
rect 23998 14702 24050 14754
rect 24050 14702 24052 14754
rect 23996 14700 24052 14702
rect 25340 15036 25396 15092
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 23548 13356 23604 13412
rect 17500 4284 17556 4340
rect 17500 3612 17556 3668
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 19740 4338 19796 4340
rect 19740 4286 19742 4338
rect 19742 4286 19794 4338
rect 19794 4286 19796 4338
rect 19740 4284 19796 4286
rect 19516 4060 19572 4116
rect 18620 3666 18676 3668
rect 18620 3614 18622 3666
rect 18622 3614 18674 3666
rect 18674 3614 18676 3666
rect 18620 3612 18676 3614
rect 20748 4114 20804 4116
rect 20748 4062 20750 4114
rect 20750 4062 20802 4114
rect 20802 4062 20804 4114
rect 20748 4060 20804 4062
rect 24220 3612 24276 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
<< metal3 >>
rect 25554 38556 25564 38612
rect 25620 38556 26796 38612
rect 26852 38556 26862 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 16818 38220 16828 38276
rect 16884 38220 18060 38276
rect 18116 38220 18126 38276
rect 24210 38220 24220 38276
rect 24276 38220 25564 38276
rect 25620 38220 25630 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 18834 37436 18844 37492
rect 18900 37436 19852 37492
rect 19908 37436 19918 37492
rect 21522 37436 21532 37492
rect 21588 37436 22764 37492
rect 22820 37436 22830 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 14354 28588 14364 28644
rect 14420 28588 15148 28644
rect 15204 28588 15214 28644
rect 19170 28476 19180 28532
rect 19236 28476 21644 28532
rect 21700 28476 22540 28532
rect 22596 28476 22606 28532
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 18722 27692 18732 27748
rect 18788 27692 20300 27748
rect 20356 27692 20366 27748
rect 22754 27692 22764 27748
rect 22820 27692 25228 27748
rect 25284 27692 25788 27748
rect 25844 27692 25854 27748
rect 0 27636 800 27664
rect 0 27580 4172 27636
rect 4228 27580 4238 27636
rect 0 27552 800 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 18834 27244 18844 27300
rect 18900 27244 19964 27300
rect 20020 27244 20030 27300
rect 17938 27020 17948 27076
rect 18004 27020 19516 27076
rect 19572 27020 19582 27076
rect 16370 26908 16380 26964
rect 16436 26908 17500 26964
rect 17556 26908 17566 26964
rect 18050 26908 18060 26964
rect 18116 26908 18732 26964
rect 18788 26908 22204 26964
rect 22260 26908 25452 26964
rect 25508 26908 25518 26964
rect 21858 26796 21868 26852
rect 21924 26796 23436 26852
rect 23492 26796 23502 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 13682 26460 13692 26516
rect 13748 26460 14588 26516
rect 14644 26460 15148 26516
rect 15204 26460 17276 26516
rect 17332 26460 17342 26516
rect 17490 26460 17500 26516
rect 17556 26460 18172 26516
rect 18228 26460 18508 26516
rect 18564 26460 19068 26516
rect 19124 26460 19134 26516
rect 17042 26348 17052 26404
rect 17108 26348 17836 26404
rect 17892 26348 18844 26404
rect 18900 26348 18910 26404
rect 41200 26292 42000 26320
rect 4274 26236 4284 26292
rect 4340 26236 11788 26292
rect 11844 26236 14700 26292
rect 14756 26236 14766 26292
rect 22418 26236 22428 26292
rect 22484 26236 24444 26292
rect 24500 26236 24510 26292
rect 40002 26236 40012 26292
rect 40068 26236 42000 26292
rect 41200 26208 42000 26236
rect 27458 26124 27468 26180
rect 27524 26124 28476 26180
rect 28532 26124 37660 26180
rect 37716 26124 37726 26180
rect 25442 25900 25452 25956
rect 25508 25900 25900 25956
rect 25956 25900 25966 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 13906 25676 13916 25732
rect 13972 25676 15820 25732
rect 15876 25676 15886 25732
rect 0 25620 800 25648
rect 0 25564 1932 25620
rect 1988 25564 1998 25620
rect 0 25536 800 25564
rect 14802 25452 14812 25508
rect 14868 25452 15260 25508
rect 15316 25452 15326 25508
rect 19394 25452 19404 25508
rect 19460 25452 21308 25508
rect 21364 25452 21374 25508
rect 24658 25452 24668 25508
rect 24724 25452 25676 25508
rect 25732 25452 25742 25508
rect 26114 25340 26124 25396
rect 26180 25340 27244 25396
rect 27300 25340 27310 25396
rect 24882 25228 24892 25284
rect 24948 25228 25564 25284
rect 25620 25228 25630 25284
rect 15474 25116 15484 25172
rect 15540 25116 17388 25172
rect 17444 25116 17454 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 41200 24948 42000 24976
rect 15698 24892 15708 24948
rect 15764 24892 16492 24948
rect 16548 24892 21980 24948
rect 22036 24892 23660 24948
rect 23716 24892 23726 24948
rect 40002 24892 40012 24948
rect 40068 24892 42000 24948
rect 41200 24864 42000 24892
rect 18610 24780 18620 24836
rect 18676 24780 18844 24836
rect 18900 24780 23996 24836
rect 24052 24780 24062 24836
rect 24210 24780 24220 24836
rect 24276 24780 26908 24836
rect 26964 24780 26974 24836
rect 30930 24780 30940 24836
rect 30996 24780 37716 24836
rect 37660 24724 37716 24780
rect 16706 24668 16716 24724
rect 16772 24668 17724 24724
rect 17780 24668 18396 24724
rect 18452 24668 18462 24724
rect 24322 24668 24332 24724
rect 24388 24668 25676 24724
rect 25732 24668 25742 24724
rect 26450 24668 26460 24724
rect 26516 24668 26796 24724
rect 26852 24668 27356 24724
rect 27412 24668 28924 24724
rect 28980 24668 28990 24724
rect 30706 24668 30716 24724
rect 30772 24668 37436 24724
rect 37492 24668 37502 24724
rect 37650 24668 37660 24724
rect 37716 24668 37726 24724
rect 12562 24444 12572 24500
rect 12628 24444 17948 24500
rect 18004 24444 18014 24500
rect 21410 24332 21420 24388
rect 21476 24332 22316 24388
rect 22372 24332 22382 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 41200 24276 42000 24304
rect 40002 24220 40012 24276
rect 40068 24220 42000 24276
rect 41200 24192 42000 24220
rect 25666 23996 25676 24052
rect 25732 23996 31948 24052
rect 31892 23940 31948 23996
rect 14802 23884 14812 23940
rect 14868 23884 16156 23940
rect 16212 23884 16222 23940
rect 17602 23884 17612 23940
rect 17668 23884 17678 23940
rect 28130 23884 28140 23940
rect 28196 23884 29260 23940
rect 29316 23884 29326 23940
rect 31892 23884 37660 23940
rect 37716 23884 37726 23940
rect 17612 23828 17668 23884
rect 17612 23772 18284 23828
rect 18340 23772 21308 23828
rect 21364 23772 21374 23828
rect 21634 23772 21644 23828
rect 21700 23772 28028 23828
rect 28084 23772 28094 23828
rect 29586 23772 29596 23828
rect 29652 23772 30268 23828
rect 30324 23772 30334 23828
rect 21410 23660 21420 23716
rect 21476 23660 21486 23716
rect 23650 23660 23660 23716
rect 23716 23660 23996 23716
rect 24052 23660 24062 23716
rect 27570 23660 27580 23716
rect 27636 23660 27646 23716
rect 21420 23604 21476 23660
rect 14914 23548 14924 23604
rect 14980 23548 15484 23604
rect 15540 23548 15550 23604
rect 21420 23548 24220 23604
rect 24276 23548 24286 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 23660 23492 23716 23548
rect 16594 23436 16604 23492
rect 16660 23436 18172 23492
rect 18228 23436 18238 23492
rect 23650 23436 23660 23492
rect 23716 23436 23726 23492
rect 27580 23380 27636 23660
rect 41200 23604 42000 23632
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 41200 23520 42000 23548
rect 19506 23324 19516 23380
rect 19572 23324 21084 23380
rect 21140 23324 22204 23380
rect 22260 23324 22270 23380
rect 26450 23324 26460 23380
rect 26516 23324 29036 23380
rect 29092 23324 29102 23380
rect 15922 23212 15932 23268
rect 15988 23212 17388 23268
rect 17444 23212 17948 23268
rect 18004 23212 18014 23268
rect 20402 23212 20412 23268
rect 20468 23212 22092 23268
rect 22148 23212 24220 23268
rect 24276 23212 24286 23268
rect 27122 23212 27132 23268
rect 27188 23212 27804 23268
rect 27860 23212 27870 23268
rect 16818 23100 16828 23156
rect 16884 23100 17612 23156
rect 17668 23100 17678 23156
rect 19730 23100 19740 23156
rect 19796 23100 21756 23156
rect 21812 23100 21822 23156
rect 31892 23100 37660 23156
rect 37716 23100 37726 23156
rect 31892 23044 31948 23100
rect 12674 22988 12684 23044
rect 12740 22988 15708 23044
rect 15764 22988 15774 23044
rect 24546 22988 24556 23044
rect 24612 22988 25340 23044
rect 25396 22988 25406 23044
rect 28578 22988 28588 23044
rect 28644 22988 29932 23044
rect 29988 22988 31948 23044
rect 41200 22932 42000 22960
rect 18946 22876 18956 22932
rect 19012 22876 20412 22932
rect 20468 22876 20478 22932
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 41200 22848 42000 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 19954 22652 19964 22708
rect 20020 22652 20860 22708
rect 20916 22652 20926 22708
rect 14690 22540 14700 22596
rect 14756 22540 15932 22596
rect 15988 22540 15998 22596
rect 17602 22540 17612 22596
rect 17668 22540 18060 22596
rect 18116 22540 18620 22596
rect 18676 22540 20076 22596
rect 20132 22540 20142 22596
rect 21634 22540 21644 22596
rect 21700 22540 25228 22596
rect 25284 22540 25294 22596
rect 21644 22484 21700 22540
rect 16370 22428 16380 22484
rect 16436 22428 17052 22484
rect 17108 22428 21700 22484
rect 24210 22316 24220 22372
rect 24276 22316 25452 22372
rect 25508 22316 26124 22372
rect 26180 22316 26190 22372
rect 27010 22316 27020 22372
rect 27076 22316 28364 22372
rect 28420 22316 29372 22372
rect 29428 22316 29438 22372
rect 15586 22204 15596 22260
rect 15652 22204 16044 22260
rect 16100 22204 16110 22260
rect 21858 22204 21868 22260
rect 21924 22204 23212 22260
rect 23268 22204 23884 22260
rect 23940 22204 23950 22260
rect 25218 22204 25228 22260
rect 25284 22204 26684 22260
rect 26740 22204 26750 22260
rect 28130 22204 28140 22260
rect 28196 22204 29036 22260
rect 29092 22204 29102 22260
rect 15596 22148 15652 22204
rect 15026 22092 15036 22148
rect 15092 22092 15652 22148
rect 16370 22092 16380 22148
rect 16436 22092 18284 22148
rect 18340 22092 18350 22148
rect 21522 22092 21532 22148
rect 21588 22092 22540 22148
rect 22596 22092 22606 22148
rect 15698 21980 15708 22036
rect 15764 21980 16604 22036
rect 16660 21980 17276 22036
rect 17332 21980 17342 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 15092 21868 15372 21924
rect 15428 21868 15438 21924
rect 15922 21868 15932 21924
rect 15988 21868 16716 21924
rect 16772 21868 16782 21924
rect 20738 21868 20748 21924
rect 20804 21868 22092 21924
rect 22148 21868 22158 21924
rect 15092 21812 15148 21868
rect 14690 21756 14700 21812
rect 14756 21756 15148 21812
rect 15092 21700 15148 21756
rect 15092 21644 17500 21700
rect 17556 21644 18396 21700
rect 18452 21644 18462 21700
rect 41200 21588 42000 21616
rect 16258 21532 16268 21588
rect 16324 21532 17836 21588
rect 17892 21532 17902 21588
rect 18610 21532 18620 21588
rect 18676 21532 18956 21588
rect 19012 21532 19022 21588
rect 40002 21532 40012 21588
rect 40068 21532 42000 21588
rect 18620 21476 18676 21532
rect 41200 21504 42000 21532
rect 4162 21420 4172 21476
rect 4228 21420 18676 21476
rect 19506 21420 19516 21476
rect 19572 21420 19582 21476
rect 29586 21420 29596 21476
rect 29652 21420 30156 21476
rect 30212 21420 37884 21476
rect 37940 21420 37950 21476
rect 19516 21252 19572 21420
rect 9986 21196 9996 21252
rect 10052 21196 19572 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 41200 20916 42000 20944
rect 8372 20860 9996 20916
rect 10052 20860 10062 20916
rect 11890 20860 11900 20916
rect 11956 20860 12908 20916
rect 12964 20860 13580 20916
rect 13636 20860 15148 20916
rect 15204 20860 15214 20916
rect 28466 20860 28476 20916
rect 28532 20860 29260 20916
rect 29316 20860 29326 20916
rect 39890 20860 39900 20916
rect 39956 20860 42000 20916
rect 8372 20804 8428 20860
rect 41200 20832 42000 20860
rect 4274 20748 4284 20804
rect 4340 20748 8428 20804
rect 20066 20748 20076 20804
rect 20132 20748 22652 20804
rect 22708 20748 22718 20804
rect 28578 20748 28588 20804
rect 28644 20748 29372 20804
rect 29428 20748 29438 20804
rect 18162 20524 18172 20580
rect 18228 20524 20188 20580
rect 20244 20524 28364 20580
rect 28420 20524 28430 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 0 20244 800 20272
rect 41200 20244 42000 20272
rect 0 20188 1932 20244
rect 1988 20188 1998 20244
rect 19282 20188 19292 20244
rect 19348 20188 21420 20244
rect 21476 20188 21486 20244
rect 40002 20188 40012 20244
rect 40068 20188 42000 20244
rect 0 20160 800 20188
rect 41200 20160 42000 20188
rect 20514 20076 20524 20132
rect 20580 20076 21532 20132
rect 21588 20076 21598 20132
rect 22082 20076 22092 20132
rect 22148 20076 23436 20132
rect 23492 20076 26124 20132
rect 26180 20076 26190 20132
rect 26348 20076 27132 20132
rect 27188 20076 27198 20132
rect 29698 20076 29708 20132
rect 29764 20076 31948 20132
rect 21532 20020 21588 20076
rect 12226 19964 12236 20020
rect 12292 19964 20300 20020
rect 20356 19964 20366 20020
rect 21532 19964 22764 20020
rect 22820 19964 22830 20020
rect 18274 19852 18284 19908
rect 18340 19852 19292 19908
rect 19348 19852 19358 19908
rect 20066 19852 20076 19908
rect 20132 19852 20636 19908
rect 20692 19852 22092 19908
rect 22148 19852 22158 19908
rect 22418 19852 22428 19908
rect 22484 19852 22876 19908
rect 22932 19852 25228 19908
rect 25284 19852 25294 19908
rect 22428 19796 22484 19852
rect 19058 19740 19068 19796
rect 19124 19740 20412 19796
rect 20468 19740 20478 19796
rect 21746 19740 21756 19796
rect 21812 19740 22484 19796
rect 19282 19628 19292 19684
rect 19348 19628 21532 19684
rect 21588 19628 22092 19684
rect 22148 19628 22158 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 26348 19572 26404 20076
rect 31892 20020 31948 20076
rect 26562 19964 26572 20020
rect 26628 19964 27356 20020
rect 27412 19964 27422 20020
rect 28354 19964 28364 20020
rect 28420 19964 29372 20020
rect 29428 19964 29438 20020
rect 31892 19964 37660 20020
rect 37716 19964 37726 20020
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 14914 19516 14924 19572
rect 14980 19516 16044 19572
rect 16100 19516 16110 19572
rect 19842 19516 19852 19572
rect 19908 19516 20972 19572
rect 21028 19516 26404 19572
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 41200 19488 42000 19516
rect 14690 19404 14700 19460
rect 14756 19404 15820 19460
rect 15876 19404 15886 19460
rect 22194 19404 22204 19460
rect 22260 19404 22540 19460
rect 22596 19404 22606 19460
rect 16146 19292 16156 19348
rect 16212 19292 16604 19348
rect 16660 19292 19628 19348
rect 19684 19292 19694 19348
rect 22418 19292 22428 19348
rect 22484 19292 23996 19348
rect 24052 19292 24062 19348
rect 26114 19292 26124 19348
rect 26180 19292 37436 19348
rect 37492 19292 37502 19348
rect 16034 19180 16044 19236
rect 16100 19180 18620 19236
rect 18676 19180 19180 19236
rect 19236 19180 19246 19236
rect 31892 19180 37660 19236
rect 37716 19180 37726 19236
rect 31892 19012 31948 19180
rect 15810 18956 15820 19012
rect 15876 18956 16492 19012
rect 16548 18956 16558 19012
rect 23314 18956 23324 19012
rect 23380 18956 26572 19012
rect 26628 18956 26638 19012
rect 27906 18956 27916 19012
rect 27972 18956 28252 19012
rect 28308 18956 31948 19012
rect 41200 18900 42000 18928
rect 40002 18844 40012 18900
rect 40068 18844 42000 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 41200 18816 42000 18844
rect 15092 18620 15820 18676
rect 15876 18620 15886 18676
rect 16034 18620 16044 18676
rect 16100 18620 16940 18676
rect 16996 18620 21532 18676
rect 21588 18620 21598 18676
rect 21970 18620 21980 18676
rect 22036 18620 25452 18676
rect 25508 18620 25518 18676
rect 29362 18620 29372 18676
rect 29428 18620 29932 18676
rect 29988 18620 37884 18676
rect 37940 18620 37950 18676
rect 15092 18564 15148 18620
rect 11666 18508 11676 18564
rect 11732 18508 15148 18564
rect 18284 18508 19628 18564
rect 19684 18508 19694 18564
rect 18284 18452 18340 18508
rect 17490 18396 17500 18452
rect 17556 18396 18340 18452
rect 18498 18396 18508 18452
rect 18564 18396 19180 18452
rect 19236 18396 19246 18452
rect 25890 18396 25900 18452
rect 25956 18396 28252 18452
rect 28308 18396 28318 18452
rect 31892 18396 37660 18452
rect 37716 18396 37726 18452
rect 31892 18340 31948 18396
rect 10098 18284 10108 18340
rect 10164 18284 11004 18340
rect 11060 18284 14252 18340
rect 14308 18284 14318 18340
rect 18396 18284 23324 18340
rect 23380 18284 23996 18340
rect 24052 18284 24062 18340
rect 24322 18284 24332 18340
rect 24388 18284 25340 18340
rect 25396 18284 25406 18340
rect 28130 18284 28140 18340
rect 28196 18284 31948 18340
rect 18396 18228 18452 18284
rect 41200 18228 42000 18256
rect 10770 18172 10780 18228
rect 10836 18172 18396 18228
rect 18452 18172 18462 18228
rect 18946 18172 18956 18228
rect 19012 18172 21308 18228
rect 21364 18172 21374 18228
rect 22194 18172 22204 18228
rect 22260 18172 23884 18228
rect 23940 18172 23950 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 18956 18116 19012 18172
rect 41200 18144 42000 18172
rect 14802 18060 14812 18116
rect 14868 18060 15708 18116
rect 15764 18060 19012 18116
rect 20850 18060 20860 18116
rect 20916 18060 26460 18116
rect 26516 18060 26526 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 22754 17948 22764 18004
rect 22820 17948 23436 18004
rect 23492 17948 23502 18004
rect 15484 17836 15596 17892
rect 15652 17836 15662 17892
rect 18050 17836 18060 17892
rect 18116 17836 22876 17892
rect 22932 17836 23100 17892
rect 23156 17836 23166 17892
rect 12898 17724 12908 17780
rect 12964 17724 14476 17780
rect 14532 17724 14542 17780
rect 15484 17220 15540 17836
rect 16146 17724 16156 17780
rect 16212 17724 17052 17780
rect 17108 17724 18620 17780
rect 18676 17724 18686 17780
rect 21186 17724 21196 17780
rect 21252 17724 21868 17780
rect 21924 17724 21934 17780
rect 16482 17612 16492 17668
rect 16548 17612 17164 17668
rect 17220 17612 17230 17668
rect 18274 17612 18284 17668
rect 18340 17612 19516 17668
rect 19572 17612 19582 17668
rect 22082 17612 22092 17668
rect 22148 17612 22596 17668
rect 25330 17612 25340 17668
rect 25396 17612 26684 17668
rect 26740 17612 26750 17668
rect 31892 17612 37660 17668
rect 37716 17612 37726 17668
rect 22540 17556 22596 17612
rect 31892 17556 31948 17612
rect 16258 17500 16268 17556
rect 16324 17500 17388 17556
rect 17444 17500 18508 17556
rect 18564 17500 18574 17556
rect 19170 17500 19180 17556
rect 19236 17500 20076 17556
rect 20132 17500 20142 17556
rect 20290 17500 20300 17556
rect 20356 17500 20524 17556
rect 20580 17500 21644 17556
rect 21700 17500 21710 17556
rect 22530 17500 22540 17556
rect 22596 17500 22606 17556
rect 24210 17500 24220 17556
rect 24276 17500 26124 17556
rect 26180 17500 26190 17556
rect 26898 17500 26908 17556
rect 26964 17500 31948 17556
rect 19618 17388 19628 17444
rect 19684 17388 21980 17444
rect 22036 17388 22046 17444
rect 23202 17388 23212 17444
rect 23268 17388 23772 17444
rect 23828 17388 24332 17444
rect 24388 17388 24398 17444
rect 27346 17388 27356 17444
rect 27412 17388 29260 17444
rect 29316 17388 29326 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 15474 17164 15484 17220
rect 15540 17164 15550 17220
rect 17938 17052 17948 17108
rect 18004 17052 20860 17108
rect 20916 17052 20926 17108
rect 21186 17052 21196 17108
rect 21252 17052 23436 17108
rect 23492 17052 23772 17108
rect 23828 17052 23838 17108
rect 13794 16940 13804 16996
rect 13860 16940 15484 16996
rect 15540 16940 15550 16996
rect 15922 16940 15932 16996
rect 15988 16940 17500 16996
rect 17556 16940 17566 16996
rect 19506 16940 19516 16996
rect 19572 16940 19964 16996
rect 20020 16940 20030 16996
rect 22754 16940 22764 16996
rect 22820 16940 26908 16996
rect 26964 16940 26974 16996
rect 41200 16884 42000 16912
rect 13570 16828 13580 16884
rect 13636 16828 14252 16884
rect 14308 16828 14812 16884
rect 14868 16828 14878 16884
rect 19394 16828 19404 16884
rect 19460 16828 20636 16884
rect 20692 16828 21420 16884
rect 21476 16828 21486 16884
rect 22866 16828 22876 16884
rect 22932 16828 23548 16884
rect 23604 16828 23614 16884
rect 40002 16828 40012 16884
rect 40068 16828 42000 16884
rect 41200 16800 42000 16828
rect 20514 16716 20524 16772
rect 20580 16716 21532 16772
rect 21588 16716 21598 16772
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 15026 16156 15036 16212
rect 15092 16156 15148 16212
rect 15204 16156 16380 16212
rect 16436 16156 16446 16212
rect 19170 15932 19180 15988
rect 19236 15932 19628 15988
rect 19684 15932 21756 15988
rect 21812 15932 21822 15988
rect 11666 15820 11676 15876
rect 11732 15820 15260 15876
rect 15316 15820 15326 15876
rect 15474 15820 15484 15876
rect 15540 15820 16492 15876
rect 16548 15820 20524 15876
rect 20580 15820 20590 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 0 15540 800 15568
rect 0 15484 1932 15540
rect 1988 15484 1998 15540
rect 0 15456 800 15484
rect 15138 15372 15148 15428
rect 15204 15372 17724 15428
rect 17780 15372 17790 15428
rect 4274 15260 4284 15316
rect 4340 15260 11676 15316
rect 11732 15260 11742 15316
rect 23986 15036 23996 15092
rect 24052 15036 25340 15092
rect 25396 15036 25406 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 18386 14700 18396 14756
rect 18452 14700 19740 14756
rect 19796 14700 19806 14756
rect 21522 14700 21532 14756
rect 21588 14700 23996 14756
rect 24052 14700 24062 14756
rect 17042 14588 17052 14644
rect 17108 14588 21420 14644
rect 21476 14588 21486 14644
rect 15586 14476 15596 14532
rect 15652 14476 16828 14532
rect 16884 14476 16894 14532
rect 17154 14476 17164 14532
rect 17220 14476 18956 14532
rect 19012 14476 19022 14532
rect 17164 14420 17220 14476
rect 16482 14364 16492 14420
rect 16548 14364 17220 14420
rect 13122 14252 13132 14308
rect 13188 14252 14812 14308
rect 14868 14252 14878 14308
rect 16258 14252 16268 14308
rect 16324 14252 17388 14308
rect 17444 14252 17454 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 12450 13692 12460 13748
rect 12516 13692 14588 13748
rect 14644 13692 14654 13748
rect 17490 13580 17500 13636
rect 17556 13580 18060 13636
rect 18116 13580 18126 13636
rect 15698 13468 15708 13524
rect 15764 13468 15774 13524
rect 15708 13412 15764 13468
rect 14690 13356 14700 13412
rect 14756 13356 18060 13412
rect 18116 13356 18126 13412
rect 20850 13356 20860 13412
rect 20916 13356 21756 13412
rect 21812 13356 23548 13412
rect 23604 13356 23614 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 15474 5180 15484 5236
rect 15540 5180 16716 5236
rect 16772 5180 16782 5236
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 17490 4284 17500 4340
rect 17556 4284 19740 4340
rect 19796 4284 19806 4340
rect 19506 4060 19516 4116
rect 19572 4060 20748 4116
rect 20804 4060 20814 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 17490 3612 17500 3668
rect 17556 3612 18620 3668
rect 18676 3612 18686 3668
rect 24210 3612 24220 3668
rect 24276 3612 25564 3668
rect 25620 3612 25630 3668
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _119_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14336 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18704 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform 1 0 19152 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _122_
timestamp 1698175906
transform 1 0 14448 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18816 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1698175906
transform -1 0 20160 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform 1 0 15232 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform 1 0 16016 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _127_
timestamp 1698175906
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698175906
transform -1 0 16016 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16240 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21392 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _131_
timestamp 1698175906
transform 1 0 19264 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform -1 0 22736 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _133_
timestamp 1698175906
transform -1 0 17696 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _134_
timestamp 1698175906
transform 1 0 17136 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _135_
timestamp 1698175906
transform -1 0 17024 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _136_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18256 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18256 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _138_
timestamp 1698175906
transform 1 0 20272 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _139_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21392 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _140_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18368 0 1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _141_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15456 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _142_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18928 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _143_
timestamp 1698175906
transform 1 0 20496 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _144_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22176 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _145_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17920 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _146_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _147_
timestamp 1698175906
transform 1 0 14560 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17696 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _149_
timestamp 1698175906
transform 1 0 16576 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _150_
timestamp 1698175906
transform 1 0 26544 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _151_
timestamp 1698175906
transform 1 0 19936 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _152_
timestamp 1698175906
transform 1 0 25984 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _153_
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _154_
timestamp 1698175906
transform -1 0 28672 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _155_
timestamp 1698175906
transform -1 0 17472 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _156_
timestamp 1698175906
transform 1 0 21504 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _157_
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _158_
timestamp 1698175906
transform -1 0 23408 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _159_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform 1 0 22624 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _161_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18368 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _162_
timestamp 1698175906
transform 1 0 22512 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _163_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24528 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _164_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18144 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _165_
timestamp 1698175906
transform -1 0 16240 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _166_
timestamp 1698175906
transform 1 0 15456 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _167_
timestamp 1698175906
transform -1 0 20496 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _168_
timestamp 1698175906
transform -1 0 22624 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _169_
timestamp 1698175906
transform 1 0 21504 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _170_
timestamp 1698175906
transform 1 0 19824 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _171_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21280 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _172_
timestamp 1698175906
transform -1 0 21392 0 -1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _173_
timestamp 1698175906
transform 1 0 20272 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _174_
timestamp 1698175906
transform 1 0 20384 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _175_
timestamp 1698175906
transform -1 0 28672 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _176_
timestamp 1698175906
transform -1 0 27888 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _177_
timestamp 1698175906
transform -1 0 18704 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _178_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16800 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _179_
timestamp 1698175906
transform 1 0 18032 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _180_
timestamp 1698175906
transform -1 0 18032 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _181_
timestamp 1698175906
transform 1 0 17808 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _182_
timestamp 1698175906
transform 1 0 16016 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _183_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _184_
timestamp 1698175906
transform 1 0 15904 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _185_
timestamp 1698175906
transform 1 0 15456 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _186_
timestamp 1698175906
transform -1 0 21952 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _187_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20160 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _188_
timestamp 1698175906
transform 1 0 19264 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _189_
timestamp 1698175906
transform -1 0 12432 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _190_
timestamp 1698175906
transform -1 0 22288 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _191_
timestamp 1698175906
transform -1 0 21840 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _192_
timestamp 1698175906
transform 1 0 19376 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _193_
timestamp 1698175906
transform -1 0 17024 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _194_
timestamp 1698175906
transform 1 0 18144 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _195_
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _196_
timestamp 1698175906
transform 1 0 23856 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _197_
timestamp 1698175906
transform 1 0 20720 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _198_
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _199_
timestamp 1698175906
transform -1 0 24304 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _200_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24080 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _201_
timestamp 1698175906
transform -1 0 25312 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _202_
timestamp 1698175906
transform 1 0 24192 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _203_
timestamp 1698175906
transform 1 0 23296 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _204_
timestamp 1698175906
transform -1 0 24528 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _205_
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _206_
timestamp 1698175906
transform -1 0 17360 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _207_
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _208_
timestamp 1698175906
transform 1 0 28000 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _209_
timestamp 1698175906
transform -1 0 27216 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _210_
timestamp 1698175906
transform 1 0 15456 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _211_
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _212_
timestamp 1698175906
transform -1 0 15568 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _213_
timestamp 1698175906
transform 1 0 15232 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _214_
timestamp 1698175906
transform -1 0 23408 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _215_
timestamp 1698175906
transform -1 0 24528 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _216_
timestamp 1698175906
transform -1 0 15904 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _217_
timestamp 1698175906
transform -1 0 15120 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _218_
timestamp 1698175906
transform -1 0 18704 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _219_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19936 0 1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _220_
timestamp 1698175906
transform -1 0 15120 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _221_
timestamp 1698175906
transform 1 0 15120 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _222_
timestamp 1698175906
transform 1 0 17136 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _223_
timestamp 1698175906
transform -1 0 27776 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _224_
timestamp 1698175906
transform -1 0 26320 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _225_
timestamp 1698175906
transform 1 0 24192 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _226_
timestamp 1698175906
transform -1 0 22624 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _227_
timestamp 1698175906
transform -1 0 19040 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _228_
timestamp 1698175906
transform 1 0 18704 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _229_
timestamp 1698175906
transform 1 0 18256 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _230_
timestamp 1698175906
transform 1 0 16240 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _231_
timestamp 1698175906
transform -1 0 16240 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _232_
timestamp 1698175906
transform -1 0 15456 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _233_
timestamp 1698175906
transform -1 0 17920 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _234_
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _235_
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _236_
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _237_
timestamp 1698175906
transform -1 0 28336 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23072 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform 1 0 27104 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _240_
timestamp 1698175906
transform 1 0 25200 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _241_
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _242_
timestamp 1698175906
transform 1 0 26880 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _243_
timestamp 1698175906
transform 1 0 9856 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _244_
timestamp 1698175906
transform 1 0 10752 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _245_
timestamp 1698175906
transform 1 0 11648 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _246_
timestamp 1698175906
transform 1 0 11648 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _247_
timestamp 1698175906
transform -1 0 13104 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _248_
timestamp 1698175906
transform 1 0 18928 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _249_
timestamp 1698175906
transform 1 0 22624 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _250_
timestamp 1698175906
transform 1 0 22624 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _251_
timestamp 1698175906
transform 1 0 21504 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _252_
timestamp 1698175906
transform 1 0 26880 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _253_
timestamp 1698175906
transform -1 0 14784 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _254_
timestamp 1698175906
transform 1 0 23856 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _255_
timestamp 1698175906
transform 1 0 12208 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _256_
timestamp 1698175906
transform -1 0 20608 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _257_
timestamp 1698175906
transform -1 0 14896 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _258_
timestamp 1698175906
transform 1 0 25424 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _259_
timestamp 1698175906
transform 1 0 21504 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _260_
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _261_
timestamp 1698175906
transform 1 0 13440 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _262_
timestamp 1698175906
transform 1 0 14448 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _263_
timestamp 1698175906
transform 1 0 27216 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _264_
timestamp 1698175906
transform -1 0 22288 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _265_
timestamp 1698175906
transform 1 0 27664 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _266_
timestamp 1698175906
transform 1 0 29232 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _267_
timestamp 1698175906
transform 1 0 30464 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__139__C dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform 1 0 26544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform 1 0 26880 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__CLK
timestamp 1698175906
transform 1 0 29232 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__CLK
timestamp 1698175906
transform 1 0 23520 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__CLK
timestamp 1698175906
transform 1 0 26656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__CLK
timestamp 1698175906
transform 1 0 13552 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__CLK
timestamp 1698175906
transform 1 0 14224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__CLK
timestamp 1698175906
transform 1 0 15120 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__CLK
timestamp 1698175906
transform 1 0 15120 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__CLK
timestamp 1698175906
transform 1 0 13552 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__CLK
timestamp 1698175906
transform -1 0 22624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__CLK
timestamp 1698175906
transform 1 0 26096 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__CLK
timestamp 1698175906
transform 1 0 26096 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__CLK
timestamp 1698175906
transform 1 0 26656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__CLK
timestamp 1698175906
transform 1 0 14784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__CLK
timestamp 1698175906
transform 1 0 27328 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__CLK
timestamp 1698175906
transform 1 0 15680 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__CLK
timestamp 1698175906
transform 1 0 20832 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__CLK
timestamp 1698175906
transform 1 0 15120 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__CLK
timestamp 1698175906
transform 1 0 28896 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__CLK
timestamp 1698175906
transform -1 0 17248 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__CLK
timestamp 1698175906
transform -1 0 17696 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__CLK
timestamp 1698175906
transform -1 0 18144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__CLK
timestamp 1698175906
transform 1 0 26432 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 18592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output22_I
timestamp 1698175906
transform -1 0 37520 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18816 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 20608 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 22512 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_158
timestamp 1698175906
transform 1 0 19040 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_162
timestamp 1698175906
transform 1 0 19488 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_189
timestamp 1698175906
transform 1 0 22512 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_205
timestamp 1698175906
transform 1 0 24304 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_123
timestamp 1698175906
transform 1 0 15120 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_153
timestamp 1698175906
transform 1 0 18480 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_169
timestamp 1698175906
transform 1 0 20272 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_173
timestamp 1698175906
transform 1 0 20720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_158 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19040 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_166
timestamp 1698175906
transform 1 0 19936 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_196
timestamp 1698175906
transform 1 0 23296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_200
timestamp 1698175906
transform 1 0 23744 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698175906
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_115
timestamp 1698175906
transform 1 0 14224 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_146
timestamp 1698175906
transform 1 0 17696 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_150
timestamp 1698175906
transform 1 0 18144 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_166
timestamp 1698175906
transform 1 0 19936 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_88
timestamp 1698175906
transform 1 0 11200 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_96
timestamp 1698175906
transform 1 0 12096 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_126
timestamp 1698175906
transform 1 0 15456 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_130
timestamp 1698175906
transform 1 0 15904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_172
timestamp 1698175906
transform 1 0 20608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_176
timestamp 1698175906
transform 1 0 21056 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_216
timestamp 1698175906
transform 1 0 25536 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_115
timestamp 1698175906
transform 1 0 14224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_131
timestamp 1698175906
transform 1 0 16016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_135
timestamp 1698175906
transform 1 0 16464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_166
timestamp 1698175906
transform 1 0 19936 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_168
timestamp 1698175906
transform 1 0 20160 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_185
timestamp 1698175906
transform 1 0 22064 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_207
timestamp 1698175906
transform 1 0 24528 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_239
timestamp 1698175906
transform 1 0 28112 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698175906
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_88
timestamp 1698175906
transform 1 0 11200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_90
timestamp 1698175906
transform 1 0 11424 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_120
timestamp 1698175906
transform 1 0 14784 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_130
timestamp 1698175906
transform 1 0 15904 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_134
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_148
timestamp 1698175906
transform 1 0 17920 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_180
timestamp 1698175906
transform 1 0 21504 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_196
timestamp 1698175906
transform 1 0 23296 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_204
timestamp 1698175906
transform 1 0 24192 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698175906
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_28
timestamp 1698175906
transform 1 0 4480 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698175906
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_115
timestamp 1698175906
transform 1 0 14224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_119
timestamp 1698175906
transform 1 0 14672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_127
timestamp 1698175906
transform 1 0 15568 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_131
timestamp 1698175906
transform 1 0 16016 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_143
timestamp 1698175906
transform 1 0 17360 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_159
timestamp 1698175906
transform 1 0 19152 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_161
timestamp 1698175906
transform 1 0 19376 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_168
timestamp 1698175906
transform 1 0 20160 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698175906
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_179
timestamp 1698175906
transform 1 0 21392 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_185
timestamp 1698175906
transform 1 0 22064 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_230
timestamp 1698175906
transform 1 0 27104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_234
timestamp 1698175906
transform 1 0 27552 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698175906
transform 1 0 28448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_104
timestamp 1698175906
transform 1 0 12992 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_120
timestamp 1698175906
transform 1 0 14784 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_132
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_158
timestamp 1698175906
transform 1 0 19040 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_186
timestamp 1698175906
transform 1 0 22176 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698175906
transform 1 0 24528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_69
timestamp 1698175906
transform 1 0 9072 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_73
timestamp 1698175906
transform 1 0 9520 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_75
timestamp 1698175906
transform 1 0 9744 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_111
timestamp 1698175906
transform 1 0 13776 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_115
timestamp 1698175906
transform 1 0 14224 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_122
timestamp 1698175906
transform 1 0 15008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_124
timestamp 1698175906
transform 1 0 15232 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_187
timestamp 1698175906
transform 1 0 22288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_207
timestamp 1698175906
transform 1 0 24528 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_211
timestamp 1698175906
transform 1 0 24976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_242
timestamp 1698175906
transform 1 0 28448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_251
timestamp 1698175906
transform 1 0 29456 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_80
timestamp 1698175906
transform 1 0 10304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_113
timestamp 1698175906
transform 1 0 14000 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_123
timestamp 1698175906
transform 1 0 15120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_125
timestamp 1698175906
transform 1 0 15344 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_135
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_150
timestamp 1698175906
transform 1 0 18144 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_179
timestamp 1698175906
transform 1 0 21392 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_187
timestamp 1698175906
transform 1 0 22288 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_189
timestamp 1698175906
transform 1 0 22512 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_203
timestamp 1698175906
transform 1 0 24080 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698175906
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_220
timestamp 1698175906
transform 1 0 25984 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_224
timestamp 1698175906
transform 1 0 26432 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_257
timestamp 1698175906
transform 1 0 30128 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_273
timestamp 1698175906
transform 1 0 31920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698175906
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_111
timestamp 1698175906
transform 1 0 13776 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_121
timestamp 1698175906
transform 1 0 14896 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_125
timestamp 1698175906
transform 1 0 15344 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_144
timestamp 1698175906
transform 1 0 17472 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698175906
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_185
timestamp 1698175906
transform 1 0 22064 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_223
timestamp 1698175906
transform 1 0 26320 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_227
timestamp 1698175906
transform 1 0 26768 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698175906
transform 1 0 28336 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_88
timestamp 1698175906
transform 1 0 11200 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_92
timestamp 1698175906
transform 1 0 11648 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_99
timestamp 1698175906
transform 1 0 12432 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_115
timestamp 1698175906
transform 1 0 14224 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_123
timestamp 1698175906
transform 1 0 15120 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_133
timestamp 1698175906
transform 1 0 16240 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_137
timestamp 1698175906
transform 1 0 16688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_148
timestamp 1698175906
transform 1 0 17920 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_156
timestamp 1698175906
transform 1 0 18816 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_195
timestamp 1698175906
transform 1 0 23184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_199
timestamp 1698175906
transform 1 0 23632 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_207
timestamp 1698175906
transform 1 0 24528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_228
timestamp 1698175906
transform 1 0 26880 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_237
timestamp 1698175906
transform 1 0 27888 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_244
timestamp 1698175906
transform 1 0 28672 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_248
timestamp 1698175906
transform 1 0 29120 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_255
timestamp 1698175906
transform 1 0 29904 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_271
timestamp 1698175906
transform 1 0 31696 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698175906
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698175906
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 9072 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 9520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 9744 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_111
timestamp 1698175906
transform 1 0 13776 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_119
timestamp 1698175906
transform 1 0 14672 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_121
timestamp 1698175906
transform 1 0 14896 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_172
timestamp 1698175906
transform 1 0 20608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698175906
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_254
timestamp 1698175906
transform 1 0 29792 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_286
timestamp 1698175906
transform 1 0 33376 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_302
timestamp 1698175906
transform 1 0 35168 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_310
timestamp 1698175906
transform 1 0 36064 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698175906
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_88
timestamp 1698175906
transform 1 0 11200 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_121
timestamp 1698175906
transform 1 0 14896 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_125
timestamp 1698175906
transform 1 0 15344 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_151
timestamp 1698175906
transform 1 0 18256 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_153
timestamp 1698175906
transform 1 0 18480 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698175906
transform 1 0 24416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_218
timestamp 1698175906
transform 1 0 25760 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_226
timestamp 1698175906
transform 1 0 26656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_259
timestamp 1698175906
transform 1 0 30352 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_275
timestamp 1698175906
transform 1 0 32144 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_318
timestamp 1698175906
transform 1 0 36960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_320
timestamp 1698175906
transform 1 0 37184 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_115
timestamp 1698175906
transform 1 0 14224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_117
timestamp 1698175906
transform 1 0 14448 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_157
timestamp 1698175906
transform 1 0 18928 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_168
timestamp 1698175906
transform 1 0 20160 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_197
timestamp 1698175906
transform 1 0 23408 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_214
timestamp 1698175906
transform 1 0 25312 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_222
timestamp 1698175906
transform 1 0 26208 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_224
timestamp 1698175906
transform 1 0 26432 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_231
timestamp 1698175906
transform 1 0 27216 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_235
timestamp 1698175906
transform 1 0 27664 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_237
timestamp 1698175906
transform 1 0 27888 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_88
timestamp 1698175906
transform 1 0 11200 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_121
timestamp 1698175906
transform 1 0 14896 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_125
timestamp 1698175906
transform 1 0 15344 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_159
timestamp 1698175906
transform 1 0 19152 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_172
timestamp 1698175906
transform 1 0 20608 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_187
timestamp 1698175906
transform 1 0 22288 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_195
timestamp 1698175906
transform 1 0 23184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_205
timestamp 1698175906
transform 1 0 24304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_226
timestamp 1698175906
transform 1 0 26656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_257
timestamp 1698175906
transform 1 0 30128 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698175906
transform 1 0 31920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_123
timestamp 1698175906
transform 1 0 15120 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_147
timestamp 1698175906
transform 1 0 17808 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_163
timestamp 1698175906
transform 1 0 19600 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698175906
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_185
timestamp 1698175906
transform 1 0 22064 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_189
timestamp 1698175906
transform 1 0 22512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_219
timestamp 1698175906
transform 1 0 25872 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_223
timestamp 1698175906
transform 1 0 26320 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_225
timestamp 1698175906
transform 1 0 26544 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_228
timestamp 1698175906
transform 1 0 26880 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698175906
transform 1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_254
timestamp 1698175906
transform 1 0 29792 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_286
timestamp 1698175906
transform 1 0 33376 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_302
timestamp 1698175906
transform 1 0 35168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_310
timestamp 1698175906
transform 1 0 36064 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698175906
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_104
timestamp 1698175906
transform 1 0 12992 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_120
timestamp 1698175906
transform 1 0 14784 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_128
timestamp 1698175906
transform 1 0 15680 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_132
timestamp 1698175906
transform 1 0 16128 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_156
timestamp 1698175906
transform 1 0 18816 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_188
timestamp 1698175906
transform 1 0 22400 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_196
timestamp 1698175906
transform 1 0 23296 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_200
timestamp 1698175906
transform 1 0 23744 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698175906
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_220
timestamp 1698175906
transform 1 0 25984 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_266
timestamp 1698175906
transform 1 0 31136 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_274
timestamp 1698175906
transform 1 0 32032 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698175906
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 36512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 37408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_115
timestamp 1698175906
transform 1 0 14224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_131
timestamp 1698175906
transform 1 0 16016 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_139
timestamp 1698175906
transform 1 0 16912 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_155
timestamp 1698175906
transform 1 0 18704 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698175906
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_182
timestamp 1698175906
transform 1 0 21728 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_198
timestamp 1698175906
transform 1 0 23520 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_202
timestamp 1698175906
transform 1 0 23968 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_212
timestamp 1698175906
transform 1 0 25088 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_223
timestamp 1698175906
transform 1 0 26320 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_236
timestamp 1698175906
transform 1 0 27776 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 4480 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_88
timestamp 1698175906
transform 1 0 11200 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_121
timestamp 1698175906
transform 1 0 14896 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_125
timestamp 1698175906
transform 1 0 15344 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_133
timestamp 1698175906
transform 1 0 16240 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_137
timestamp 1698175906
transform 1 0 16688 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_146
timestamp 1698175906
transform 1 0 17696 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_153
timestamp 1698175906
transform 1 0 18480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_163
timestamp 1698175906
transform 1 0 19600 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_171
timestamp 1698175906
transform 1 0 20496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_175
timestamp 1698175906
transform 1 0 20944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_183
timestamp 1698175906
transform 1 0 21840 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_191
timestamp 1698175906
transform 1 0 22736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_195
timestamp 1698175906
transform 1 0 23184 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_214
timestamp 1698175906
transform 1 0 25312 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_244
timestamp 1698175906
transform 1 0 28672 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_248
timestamp 1698175906
transform 1 0 29120 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_123
timestamp 1698175906
transform 1 0 15120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698175906
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_219
timestamp 1698175906
transform 1 0 25872 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_223
timestamp 1698175906
transform 1 0 26320 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_239
timestamp 1698175906
transform 1 0 28112 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698175906
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_104
timestamp 1698175906
transform 1 0 12992 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_137
timestamp 1698175906
transform 1 0 16688 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698175906
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_171
timestamp 1698175906
transform 1 0 20496 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_179
timestamp 1698175906
transform 1 0 21392 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_216
timestamp 1698175906
transform 1 0 25536 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_115
timestamp 1698175906
transform 1 0 14224 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_119
timestamp 1698175906
transform 1 0 14672 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_121
timestamp 1698175906
transform 1 0 14896 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_126
timestamp 1698175906
transform 1 0 15456 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_134
timestamp 1698175906
transform 1 0 16352 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_138
timestamp 1698175906
transform 1 0 16800 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_142
timestamp 1698175906
transform 1 0 17248 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_146
timestamp 1698175906
transform 1 0 17696 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_150
timestamp 1698175906
transform 1 0 18144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_152
timestamp 1698175906
transform 1 0 18368 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_158
timestamp 1698175906
transform 1 0 19040 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698175906
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_187
timestamp 1698175906
transform 1 0 22288 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_219
timestamp 1698175906
transform 1 0 25872 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_235
timestamp 1698175906
transform 1 0 27664 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_243
timestamp 1698175906
transform 1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_150
timestamp 1698175906
transform 1 0 18144 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_154
timestamp 1698175906
transform 1 0 18592 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_156
timestamp 1698175906
transform 1 0 18816 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_186
timestamp 1698175906
transform 1 0 22176 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_190
timestamp 1698175906
transform 1 0 22624 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_150
timestamp 1698175906
transform 1 0 18144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_154
timestamp 1698175906
transform 1 0 18592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 25536 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_243
timestamp 1698175906
transform 1 0 28560 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698175906
transform 1 0 32144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_165
timestamp 1698175906
transform 1 0 19824 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_169
timestamp 1698175906
transform 1 0 20272 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37520 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 25648 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 18704 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 4480 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 37520 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 37520 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 21280 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 21616 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform -1 0 4480 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 19600 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 4480 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 24192 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 15568 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 16912 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 17472 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698175906
transform 1 0 37520 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 41200 24864 42000 24976 0 FreeSans 448 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 25536 41200 25648 42000 0 FreeSans 448 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 24192 41200 24304 42000 0 FreeSans 448 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 18816 41200 18928 42000 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 0 15456 800 15568 0 FreeSans 448 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 41200 18816 42000 18928 0 FreeSans 448 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 41200 26208 42000 26320 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 41200 16800 42000 16912 0 FreeSans 448 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 41200 20160 42000 20272 0 FreeSans 448 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 21504 41200 21616 42000 0 FreeSans 448 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 41200 21504 42000 21616 0 FreeSans 448 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 16800 41200 16912 42000 0 FreeSans 448 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 41200 24192 42000 24304 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 27776 18536 27776 18536 0 _000_
rlabel metal2 10808 17976 10808 17976 0 _001_
rlabel metal3 13412 18536 13412 18536 0 _002_
rlabel metal2 12600 23856 12600 23856 0 _003_
rlabel metal2 12656 21672 12656 21672 0 _004_
rlabel metal2 11928 20440 11928 20440 0 _005_
rlabel metal2 19656 28224 19656 28224 0 _006_
rlabel metal2 24024 23520 24024 23520 0 _007_
rlabel metal2 23576 26712 23576 26712 0 _008_
rlabel metal2 21896 14224 21896 14224 0 _009_
rlabel metal3 27496 23240 27496 23240 0 _010_
rlabel metal2 13832 16184 13832 16184 0 _011_
rlabel metal2 24248 16464 24248 16464 0 _012_
rlabel metal2 13160 14056 13160 14056 0 _013_
rlabel metal2 19656 14280 19656 14280 0 _014_
rlabel metal2 13944 25928 13944 25928 0 _015_
rlabel metal2 25816 25872 25816 25872 0 _016_
rlabel metal2 22120 27440 22120 27440 0 _017_
rlabel metal2 18200 27300 18200 27300 0 _018_
rlabel metal2 14392 28280 14392 28280 0 _019_
rlabel metal2 15456 13048 15456 13048 0 _020_
rlabel metal2 28112 24136 28112 24136 0 _021_
rlabel metal3 23240 19320 23240 19320 0 _022_
rlabel metal2 28168 21112 28168 21112 0 _023_
rlabel metal3 25200 17528 25200 17528 0 _024_
rlabel metal2 21000 13272 21000 13272 0 _025_
rlabel metal2 19656 20832 19656 20832 0 _026_
rlabel metal3 19432 27272 19432 27272 0 _027_
rlabel metal2 20104 19936 20104 19936 0 _028_
rlabel metal2 22568 17192 22568 17192 0 _029_
rlabel metal3 21112 17528 21112 17528 0 _030_
rlabel metal3 21560 17752 21560 17752 0 _031_
rlabel metal2 20384 18312 20384 18312 0 _032_
rlabel metal2 26600 19936 26600 19936 0 _033_
rlabel metal2 28000 19992 28000 19992 0 _034_
rlabel metal2 17528 26992 17528 26992 0 _035_
rlabel metal2 18928 28504 18928 28504 0 _036_
rlabel metal3 18760 27048 18760 27048 0 _037_
rlabel metal2 16968 24360 16968 24360 0 _038_
rlabel metal2 16128 22456 16128 22456 0 _039_
rlabel metal2 21448 20048 21448 20048 0 _040_
rlabel metal2 19544 20608 19544 20608 0 _041_
rlabel metal3 16296 19992 16296 19992 0 _042_
rlabel metal2 21784 26040 21784 26040 0 _043_
rlabel metal2 20328 26964 20328 26964 0 _044_
rlabel metal3 16128 24920 16128 24920 0 _045_
rlabel metal3 18760 24808 18760 24808 0 _046_
rlabel metal2 25368 22400 25368 22400 0 _047_
rlabel metal2 24136 23968 24136 23968 0 _048_
rlabel metal2 21224 23240 21224 23240 0 _049_
rlabel metal2 23688 23408 23688 23408 0 _050_
rlabel metal2 23520 26264 23520 26264 0 _051_
rlabel metal2 24920 23912 24920 23912 0 _052_
rlabel metal2 24360 25592 24360 25592 0 _053_
rlabel metal3 22792 14728 22792 14728 0 _054_
rlabel metal2 16968 15204 16968 15204 0 _055_
rlabel metal3 19264 14616 19264 14616 0 _056_
rlabel metal2 28280 23016 28280 23016 0 _057_
rlabel metal2 15736 17304 15736 17304 0 _058_
rlabel metal3 16464 15400 16464 15400 0 _059_
rlabel metal2 15288 16576 15288 16576 0 _060_
rlabel metal2 22904 16800 22904 16800 0 _061_
rlabel metal2 15008 14728 15008 14728 0 _062_
rlabel metal3 19096 14728 19096 14728 0 _063_
rlabel metal3 15064 25480 15064 25480 0 _064_
rlabel metal3 23856 26936 23856 26936 0 _065_
rlabel metal3 26712 25368 26712 25368 0 _066_
rlabel metal2 24472 26152 24472 26152 0 _067_
rlabel metal2 18424 27832 18424 27832 0 _068_
rlabel metal2 19432 25760 19432 25760 0 _069_
rlabel metal2 16184 27160 16184 27160 0 _070_
rlabel metal2 15512 27888 15512 27888 0 _071_
rlabel metal2 16296 14056 16296 14056 0 _072_
rlabel metal2 21672 24528 21672 24528 0 _073_
rlabel metal3 28728 23912 28728 23912 0 _074_
rlabel metal2 14840 17808 14840 17808 0 _075_
rlabel metal2 19208 18480 19208 18480 0 _076_
rlabel metal2 22120 19040 22120 19040 0 _077_
rlabel metal2 14952 19096 14952 19096 0 _078_
rlabel metal2 18312 18032 18312 18032 0 _079_
rlabel metal2 21784 17808 21784 17808 0 _080_
rlabel metal2 16296 17584 16296 17584 0 _081_
rlabel metal2 16520 17584 16520 17584 0 _082_
rlabel metal2 17024 21672 17024 21672 0 _083_
rlabel metal2 14952 24472 14952 24472 0 _084_
rlabel metal2 15512 16128 15512 16128 0 _085_
rlabel metal2 22288 17080 22288 17080 0 _086_
rlabel metal2 22568 21168 22568 21168 0 _087_
rlabel metal2 19768 26908 19768 26908 0 _088_
rlabel metal3 17584 24696 17584 24696 0 _089_
rlabel via2 17640 23128 17640 23128 0 _090_
rlabel metal2 18312 24976 18312 24976 0 _091_
rlabel metal3 16688 23240 16688 23240 0 _092_
rlabel metal2 20440 22624 20440 22624 0 _093_
rlabel metal2 22008 19712 22008 19712 0 _094_
rlabel metal2 22344 20048 22344 20048 0 _095_
rlabel metal3 21056 16856 21056 16856 0 _096_
rlabel metal2 18312 23184 18312 23184 0 _097_
rlabel metal2 17976 17752 17976 17752 0 _098_
rlabel metal2 23800 16856 23800 16856 0 _099_
rlabel metal2 17640 21000 17640 21000 0 _100_
rlabel metal2 14840 23128 14840 23128 0 _101_
rlabel metal2 16184 22232 16184 22232 0 _102_
rlabel metal2 20216 19880 20216 19880 0 _103_
rlabel metal2 25256 22288 25256 22288 0 _104_
rlabel metal3 28896 22344 28896 22344 0 _105_
rlabel metal3 21280 23240 21280 23240 0 _106_
rlabel metal3 28616 22232 28616 22232 0 _107_
rlabel metal2 28504 20832 28504 20832 0 _108_
rlabel metal2 16968 18816 16968 18816 0 _109_
rlabel metal2 24024 17752 24024 17752 0 _110_
rlabel metal3 22568 22232 22568 22232 0 _111_
rlabel metal2 25256 19992 25256 19992 0 _112_
rlabel metal2 24360 17976 24360 17976 0 _113_
rlabel metal2 23128 19264 23128 19264 0 _114_
rlabel metal3 20496 17864 20496 17864 0 _115_
rlabel metal2 23800 17528 23800 17528 0 _116_
rlabel metal2 21000 19824 21000 19824 0 _117_
rlabel metal2 15680 19320 15680 19320 0 _118_
rlabel metal3 2478 27608 2478 27608 0 clk
rlabel metal2 22680 21112 22680 21112 0 clknet_0_clk
rlabel metal2 17416 28392 17416 28392 0 clknet_1_0__leaf_clk
rlabel metal2 21672 28168 21672 28168 0 clknet_1_1__leaf_clk
rlabel metal2 14504 18088 14504 18088 0 dut32.count\[0\]
rlabel metal2 14616 18928 14616 18928 0 dut32.count\[1\]
rlabel metal2 14728 22792 14728 22792 0 dut32.count\[2\]
rlabel metal2 14728 21616 14728 21616 0 dut32.count\[3\]
rlabel metal2 30296 24640 30296 24640 0 net1
rlabel metal2 29960 18480 29960 18480 0 net10
rlabel metal2 28616 22624 28616 22624 0 net11
rlabel metal3 31920 23968 31920 23968 0 net12
rlabel metal2 21784 33264 21784 33264 0 net13
rlabel metal2 22064 29288 22064 29288 0 net14
rlabel metal3 6356 20776 6356 20776 0 net15
rlabel metal2 17472 4312 17472 4312 0 net16
rlabel metal2 11816 26208 11816 26208 0 net17
rlabel metal2 28168 18648 28168 18648 0 net18
rlabel metal2 21896 16268 21896 16268 0 net19
rlabel metal2 25704 29540 25704 29540 0 net2
rlabel metal2 29624 21056 29624 21056 0 net20
rlabel metal2 15288 12432 15288 12432 0 net21
rlabel metal2 37688 21504 37688 21504 0 net22
rlabel metal3 30828 20104 30828 20104 0 net23
rlabel metal2 16520 28112 16520 28112 0 net24
rlabel metal2 17640 7644 17640 7644 0 net25
rlabel metal3 37688 24752 37688 24752 0 net26
rlabel metal2 24528 27720 24528 27720 0 net3
rlabel metal2 18760 28112 18760 28112 0 net4
rlabel metal2 24584 8568 24584 8568 0 net5
rlabel metal2 4312 15680 4312 15680 0 net6
rlabel metal2 27944 19096 27944 19096 0 net7
rlabel metal2 27496 25760 27496 25760 0 net8
rlabel metal2 26936 16856 26936 16856 0 net9
rlabel metal2 40040 25256 40040 25256 0 segm[0]
rlabel metal2 25592 39914 25592 39914 0 segm[10]
rlabel metal2 24248 39746 24248 39746 0 segm[11]
rlabel metal3 19376 37464 19376 37464 0 segm[12]
rlabel metal3 24920 3640 24920 3640 0 segm[13]
rlabel metal3 1358 15512 1358 15512 0 segm[1]
rlabel metal2 40040 19096 40040 19096 0 segm[2]
rlabel metal2 40040 26712 40040 26712 0 segm[3]
rlabel metal2 40040 17304 40040 17304 0 segm[4]
rlabel metal2 40040 20552 40040 20552 0 segm[5]
rlabel metal3 40642 22904 40642 22904 0 segm[6]
rlabel metal2 40040 23800 40040 23800 0 segm[7]
rlabel metal2 22232 39746 22232 39746 0 segm[8]
rlabel metal2 21560 39354 21560 39354 0 segm[9]
rlabel metal3 1358 20216 1358 20216 0 sel[0]
rlabel metal3 20160 4088 20160 4088 0 sel[10]
rlabel metal3 1358 25592 1358 25592 0 sel[11]
rlabel metal3 40642 18200 40642 18200 0 sel[1]
rlabel metal2 22232 2086 22232 2086 0 sel[2]
rlabel metal2 40040 22008 40040 22008 0 sel[3]
rlabel metal3 16128 5208 16128 5208 0 sel[4]
rlabel metal2 39928 21168 39928 21168 0 sel[5]
rlabel metal2 40040 19656 40040 19656 0 sel[6]
rlabel metal2 16856 39746 16856 39746 0 sel[7]
rlabel metal3 18088 3640 18088 3640 0 sel[8]
rlabel metal2 40040 24360 40040 24360 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
