magic
tech gf180mcuD
magscale 1 5
timestamp 1699641901
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9591 19137 9617 19143
rect 9591 19105 9617 19111
rect 11047 19137 11073 19143
rect 11047 19105 11073 19111
rect 13063 19137 13089 19143
rect 13063 19105 13089 19111
rect 9865 18999 9871 19025
rect 9897 18999 9903 19025
rect 10537 18999 10543 19025
rect 10569 18999 10575 19025
rect 12609 18999 12615 19025
rect 12641 18999 12647 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 9199 18745 9225 18751
rect 9199 18713 9225 18719
rect 10711 18745 10737 18751
rect 10711 18713 10737 18719
rect 13399 18745 13425 18751
rect 13399 18713 13425 18719
rect 855 18689 881 18695
rect 855 18657 881 18663
rect 8689 18607 8695 18633
rect 8721 18607 8727 18633
rect 10425 18607 10431 18633
rect 10457 18607 10463 18633
rect 12889 18607 12895 18633
rect 12921 18607 12927 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 10369 13567 10375 13593
rect 10401 13567 10407 13593
rect 8913 13511 8919 13537
rect 8945 13511 8951 13537
rect 10711 13481 10737 13487
rect 9305 13455 9311 13481
rect 9337 13455 9343 13481
rect 10711 13449 10737 13455
rect 8415 13425 8441 13431
rect 8415 13393 8441 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 10487 13257 10513 13263
rect 10487 13225 10513 13231
rect 10767 13201 10793 13207
rect 10767 13169 10793 13175
rect 10375 13145 10401 13151
rect 6897 13119 6903 13145
rect 6929 13119 6935 13145
rect 8857 13119 8863 13145
rect 8889 13119 8895 13145
rect 10375 13113 10401 13119
rect 10543 13145 10569 13151
rect 10543 13113 10569 13119
rect 10823 13145 10849 13151
rect 10823 13113 10849 13119
rect 11047 13089 11073 13095
rect 7233 13063 7239 13089
rect 7265 13063 7271 13089
rect 8297 13063 8303 13089
rect 8329 13063 8335 13089
rect 9193 13063 9199 13089
rect 9225 13063 9231 13089
rect 10257 13063 10263 13089
rect 10289 13063 10295 13089
rect 11047 13057 11073 13063
rect 10767 13033 10793 13039
rect 10767 13001 10793 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 8191 12865 8217 12871
rect 8191 12833 8217 12839
rect 10151 12865 10177 12871
rect 10151 12833 10177 12839
rect 967 12809 993 12815
rect 20007 12809 20033 12815
rect 12833 12783 12839 12809
rect 12865 12783 12871 12809
rect 967 12777 993 12783
rect 20007 12777 20033 12783
rect 7855 12753 7881 12759
rect 2137 12727 2143 12753
rect 2169 12727 2175 12753
rect 7855 12721 7881 12727
rect 9759 12753 9785 12759
rect 9759 12721 9785 12727
rect 9927 12753 9953 12759
rect 9927 12721 9953 12727
rect 10207 12753 10233 12759
rect 11321 12727 11327 12753
rect 11353 12727 11359 12753
rect 18825 12727 18831 12753
rect 18857 12727 18863 12753
rect 10207 12721 10233 12727
rect 7911 12697 7937 12703
rect 7911 12665 7937 12671
rect 8023 12697 8049 12703
rect 8023 12665 8049 12671
rect 8135 12697 8161 12703
rect 11713 12671 11719 12697
rect 11745 12671 11751 12697
rect 8135 12665 8161 12671
rect 8191 12641 8217 12647
rect 8191 12609 8217 12615
rect 9871 12641 9897 12647
rect 9871 12609 9897 12615
rect 10151 12641 10177 12647
rect 10151 12609 10177 12615
rect 11159 12641 11185 12647
rect 11159 12609 11185 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 7351 12473 7377 12479
rect 7351 12441 7377 12447
rect 12615 12473 12641 12479
rect 12615 12441 12641 12447
rect 12951 12473 12977 12479
rect 13113 12447 13119 12473
rect 13145 12447 13151 12473
rect 12951 12441 12977 12447
rect 12777 12391 12783 12417
rect 12809 12391 12815 12417
rect 7463 12361 7489 12367
rect 9871 12361 9897 12367
rect 7009 12335 7015 12361
rect 7041 12335 7047 12361
rect 7233 12335 7239 12361
rect 7265 12335 7271 12361
rect 7569 12335 7575 12361
rect 7601 12335 7607 12361
rect 7463 12329 7489 12335
rect 9871 12329 9897 12335
rect 9927 12361 9953 12367
rect 9927 12329 9953 12335
rect 9983 12361 10009 12367
rect 9983 12329 10009 12335
rect 10039 12361 10065 12367
rect 10039 12329 10065 12335
rect 10095 12361 10121 12367
rect 10929 12335 10935 12361
rect 10961 12335 10967 12361
rect 18825 12335 18831 12361
rect 18857 12335 18863 12361
rect 10095 12329 10121 12335
rect 7407 12305 7433 12311
rect 5609 12279 5615 12305
rect 5641 12279 5647 12305
rect 6673 12279 6679 12305
rect 6705 12279 6711 12305
rect 7407 12273 7433 12279
rect 10711 12305 10737 12311
rect 11265 12279 11271 12305
rect 11297 12279 11303 12305
rect 12329 12279 12335 12305
rect 12361 12279 12367 12305
rect 10711 12273 10737 12279
rect 20007 12249 20033 12255
rect 20007 12217 20033 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 6735 12081 6761 12087
rect 6735 12049 6761 12055
rect 6791 12025 6817 12031
rect 6791 11993 6817 11999
rect 7183 12025 7209 12031
rect 11439 12025 11465 12031
rect 9921 11999 9927 12025
rect 9953 11999 9959 12025
rect 7183 11993 7209 11999
rect 11439 11993 11465 11999
rect 11887 12025 11913 12031
rect 11887 11993 11913 11999
rect 11327 11969 11353 11975
rect 8521 11943 8527 11969
rect 8553 11943 8559 11969
rect 11327 11937 11353 11943
rect 11551 11969 11577 11975
rect 11551 11937 11577 11943
rect 11663 11969 11689 11975
rect 11663 11937 11689 11943
rect 11943 11969 11969 11975
rect 11943 11937 11969 11943
rect 12055 11969 12081 11975
rect 12055 11937 12081 11943
rect 12447 11969 12473 11975
rect 12447 11937 12473 11943
rect 10655 11913 10681 11919
rect 7625 11887 7631 11913
rect 7657 11887 7663 11913
rect 8857 11887 8863 11913
rect 8889 11887 8895 11913
rect 10655 11881 10681 11887
rect 10823 11913 10849 11919
rect 10823 11881 10849 11887
rect 11831 11913 11857 11919
rect 11831 11881 11857 11887
rect 12279 11913 12305 11919
rect 12279 11881 12305 11887
rect 12335 11913 12361 11919
rect 12335 11881 12361 11887
rect 7799 11857 7825 11863
rect 7799 11825 7825 11831
rect 10151 11857 10177 11863
rect 10151 11825 10177 11831
rect 10711 11857 10737 11863
rect 10711 11825 10737 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 7743 11689 7769 11695
rect 7743 11657 7769 11663
rect 11775 11689 11801 11695
rect 11775 11657 11801 11663
rect 11887 11689 11913 11695
rect 11887 11657 11913 11663
rect 11719 11577 11745 11583
rect 6113 11551 6119 11577
rect 6145 11551 6151 11577
rect 11377 11551 11383 11577
rect 11409 11551 11415 11577
rect 11719 11545 11745 11551
rect 6449 11495 6455 11521
rect 6481 11495 6487 11521
rect 7513 11495 7519 11521
rect 7545 11495 7551 11521
rect 10257 11495 10263 11521
rect 10289 11495 10295 11521
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 8807 11297 8833 11303
rect 8807 11265 8833 11271
rect 11159 11297 11185 11303
rect 11159 11265 11185 11271
rect 967 11241 993 11247
rect 6399 11241 6425 11247
rect 4713 11215 4719 11241
rect 4745 11215 4751 11241
rect 967 11209 993 11215
rect 6399 11209 6425 11215
rect 8415 11241 8441 11247
rect 8415 11209 8441 11215
rect 9535 11241 9561 11247
rect 20007 11241 20033 11247
rect 11041 11215 11047 11241
rect 11073 11215 11079 11241
rect 9535 11209 9561 11215
rect 20007 11209 20033 11215
rect 8471 11185 8497 11191
rect 2137 11159 2143 11185
rect 2169 11159 2175 11185
rect 6113 11159 6119 11185
rect 6145 11159 6151 11185
rect 7905 11159 7911 11185
rect 7937 11159 7943 11185
rect 8471 11153 8497 11159
rect 8639 11185 8665 11191
rect 9423 11185 9449 11191
rect 8969 11159 8975 11185
rect 9001 11159 9007 11185
rect 8639 11153 8665 11159
rect 9423 11153 9449 11159
rect 9647 11185 9673 11191
rect 9647 11153 9673 11159
rect 9759 11185 9785 11191
rect 9759 11153 9785 11159
rect 10039 11185 10065 11191
rect 10039 11153 10065 11159
rect 10207 11185 10233 11191
rect 10207 11153 10233 11159
rect 10319 11185 10345 11191
rect 11321 11159 11327 11185
rect 11353 11159 11359 11185
rect 11433 11159 11439 11185
rect 11465 11159 11471 11185
rect 11713 11159 11719 11185
rect 11745 11159 11751 11185
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 10319 11153 10345 11159
rect 8135 11129 8161 11135
rect 9927 11129 9953 11135
rect 5777 11103 5783 11129
rect 5809 11103 5815 11129
rect 9025 11103 9031 11129
rect 9057 11103 9063 11129
rect 8135 11097 8161 11103
rect 9927 11097 9953 11103
rect 10823 11129 10849 11135
rect 10873 11103 10879 11129
rect 10905 11103 10911 11129
rect 10823 11097 10849 11103
rect 8191 11073 8217 11079
rect 7793 11047 7799 11073
rect 7825 11047 7831 11073
rect 8191 11041 8217 11047
rect 8303 11073 8329 11079
rect 8303 11041 8329 11047
rect 8751 11073 8777 11079
rect 10375 11073 10401 11079
rect 9249 11047 9255 11073
rect 9281 11047 9287 11073
rect 8751 11041 8777 11047
rect 10375 11041 10401 11047
rect 10655 11073 10681 11079
rect 10655 11041 10681 11047
rect 10767 11073 10793 11079
rect 10767 11041 10793 11047
rect 11215 11073 11241 11079
rect 11601 11047 11607 11073
rect 11633 11047 11639 11073
rect 11215 11041 11241 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 6175 10905 6201 10911
rect 6175 10873 6201 10879
rect 6287 10905 6313 10911
rect 6287 10873 6313 10879
rect 6623 10905 6649 10911
rect 6623 10873 6649 10879
rect 6679 10905 6705 10911
rect 8415 10905 8441 10911
rect 7625 10879 7631 10905
rect 7657 10879 7663 10905
rect 8745 10879 8751 10905
rect 8777 10879 8783 10905
rect 9921 10879 9927 10905
rect 9953 10879 9959 10905
rect 6679 10873 6705 10879
rect 8415 10873 8441 10879
rect 5839 10849 5865 10855
rect 5839 10817 5865 10823
rect 7407 10849 7433 10855
rect 8241 10823 8247 10849
rect 8273 10823 8279 10849
rect 8969 10823 8975 10849
rect 9001 10823 9007 10849
rect 9081 10823 9087 10849
rect 9113 10823 9119 10849
rect 10369 10823 10375 10849
rect 10401 10823 10407 10849
rect 13337 10823 13343 10849
rect 13369 10823 13375 10849
rect 7407 10817 7433 10823
rect 6399 10793 6425 10799
rect 6399 10761 6425 10767
rect 6567 10793 6593 10799
rect 6567 10761 6593 10767
rect 6903 10793 6929 10799
rect 6903 10761 6929 10767
rect 7799 10793 7825 10799
rect 7799 10761 7825 10767
rect 8695 10793 8721 10799
rect 11047 10793 11073 10799
rect 11439 10793 11465 10799
rect 9809 10767 9815 10793
rect 9841 10767 9847 10793
rect 10537 10767 10543 10793
rect 10569 10767 10575 10793
rect 10817 10767 10823 10793
rect 10849 10767 10855 10793
rect 11209 10767 11215 10793
rect 11241 10767 11247 10793
rect 8695 10761 8721 10767
rect 11047 10761 11073 10767
rect 11439 10761 11465 10767
rect 11551 10793 11577 10799
rect 11551 10761 11577 10767
rect 13175 10793 13201 10799
rect 18825 10767 18831 10793
rect 18857 10767 18863 10793
rect 13175 10761 13201 10767
rect 5951 10737 5977 10743
rect 5777 10711 5783 10737
rect 5809 10711 5815 10737
rect 5951 10705 5977 10711
rect 6343 10737 6369 10743
rect 6343 10705 6369 10711
rect 7127 10737 7153 10743
rect 11495 10737 11521 10743
rect 10313 10711 10319 10737
rect 10345 10711 10351 10737
rect 7127 10705 7153 10711
rect 11495 10705 11521 10711
rect 7295 10681 7321 10687
rect 7295 10649 7321 10655
rect 11327 10681 11353 10687
rect 11327 10649 11353 10655
rect 20007 10681 20033 10687
rect 20007 10649 20033 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 9585 10487 9591 10513
rect 9617 10487 9623 10513
rect 10319 10457 10345 10463
rect 10319 10425 10345 10431
rect 10935 10457 10961 10463
rect 11265 10431 11271 10457
rect 11297 10431 11303 10457
rect 12273 10431 12279 10457
rect 12305 10431 12311 10457
rect 13337 10431 13343 10457
rect 13369 10431 13375 10457
rect 10935 10425 10961 10431
rect 6119 10401 6145 10407
rect 6119 10369 6145 10375
rect 6231 10401 6257 10407
rect 6231 10369 6257 10375
rect 6679 10401 6705 10407
rect 6679 10369 6705 10375
rect 6847 10401 6873 10407
rect 6847 10369 6873 10375
rect 9759 10401 9785 10407
rect 9759 10369 9785 10375
rect 9871 10401 9897 10407
rect 10263 10401 10289 10407
rect 10089 10375 10095 10401
rect 10121 10375 10127 10401
rect 9871 10369 9897 10375
rect 10263 10369 10289 10375
rect 10991 10401 11017 10407
rect 10991 10369 11017 10375
rect 11159 10401 11185 10407
rect 11159 10369 11185 10375
rect 11719 10401 11745 10407
rect 11881 10375 11887 10401
rect 11913 10375 11919 10401
rect 11719 10369 11745 10375
rect 6791 10345 6817 10351
rect 8079 10345 8105 10351
rect 8863 10345 8889 10351
rect 7905 10319 7911 10345
rect 7937 10319 7943 10345
rect 8689 10319 8695 10345
rect 8721 10319 8727 10345
rect 6791 10313 6817 10319
rect 8079 10313 8105 10319
rect 8863 10313 8889 10319
rect 10767 10345 10793 10351
rect 10767 10313 10793 10319
rect 6175 10289 6201 10295
rect 6175 10257 6201 10263
rect 6343 10289 6369 10295
rect 6343 10257 6369 10263
rect 8527 10289 8553 10295
rect 9255 10289 9281 10295
rect 9025 10263 9031 10289
rect 9057 10263 9063 10289
rect 8527 10257 8553 10263
rect 9255 10257 9281 10263
rect 10375 10289 10401 10295
rect 10375 10257 10401 10263
rect 10879 10289 10905 10295
rect 10879 10257 10905 10263
rect 11271 10289 11297 10295
rect 11271 10257 11297 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 6343 10121 6369 10127
rect 6343 10089 6369 10095
rect 7351 10121 7377 10127
rect 7351 10089 7377 10095
rect 7463 10121 7489 10127
rect 7463 10089 7489 10095
rect 6455 10065 6481 10071
rect 5833 10039 5839 10065
rect 5865 10039 5871 10065
rect 6455 10033 6481 10039
rect 6735 10065 6761 10071
rect 6735 10033 6761 10039
rect 8695 10065 8721 10071
rect 8695 10033 8721 10039
rect 8751 10065 8777 10071
rect 8751 10033 8777 10039
rect 9143 10065 9169 10071
rect 9143 10033 9169 10039
rect 12671 10065 12697 10071
rect 12671 10033 12697 10039
rect 12727 10065 12753 10071
rect 12727 10033 12753 10039
rect 6511 10009 6537 10015
rect 2137 9983 2143 10009
rect 2169 9983 2175 10009
rect 6225 9983 6231 10009
rect 6257 9983 6263 10009
rect 6511 9977 6537 9983
rect 7687 10009 7713 10015
rect 7687 9977 7713 9983
rect 8863 10009 8889 10015
rect 8969 9983 8975 10009
rect 9001 9983 9007 10009
rect 9305 9983 9311 10009
rect 9337 9983 9343 10009
rect 8863 9977 8889 9983
rect 7407 9953 7433 9959
rect 4769 9927 4775 9953
rect 4801 9927 4807 9953
rect 7407 9921 7433 9927
rect 9087 9953 9113 9959
rect 11713 9927 11719 9953
rect 11745 9927 11751 9953
rect 9087 9921 9113 9927
rect 967 9897 993 9903
rect 967 9865 993 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 8023 9729 8049 9735
rect 8241 9703 8247 9729
rect 8273 9703 8279 9729
rect 8023 9697 8049 9703
rect 20007 9673 20033 9679
rect 8409 9647 8415 9673
rect 8441 9647 8447 9673
rect 11601 9647 11607 9673
rect 11633 9647 11639 9673
rect 12217 9647 12223 9673
rect 12249 9647 12255 9673
rect 13281 9647 13287 9673
rect 13313 9647 13319 9673
rect 20007 9641 20033 9647
rect 7351 9617 7377 9623
rect 9815 9617 9841 9623
rect 8465 9591 8471 9617
rect 8497 9591 8503 9617
rect 8801 9591 8807 9617
rect 8833 9591 8839 9617
rect 9305 9591 9311 9617
rect 9337 9591 9343 9617
rect 7351 9585 7377 9591
rect 9815 9585 9841 9591
rect 10599 9617 10625 9623
rect 10599 9585 10625 9591
rect 10879 9617 10905 9623
rect 10879 9585 10905 9591
rect 10991 9617 11017 9623
rect 10991 9585 11017 9591
rect 11103 9617 11129 9623
rect 11657 9591 11663 9617
rect 11689 9591 11695 9617
rect 11825 9591 11831 9617
rect 11857 9591 11863 9617
rect 18825 9591 18831 9617
rect 18857 9591 18863 9617
rect 11103 9585 11129 9591
rect 7967 9561 7993 9567
rect 11495 9561 11521 9567
rect 7177 9535 7183 9561
rect 7209 9535 7215 9561
rect 10033 9535 10039 9561
rect 10065 9535 10071 9561
rect 10313 9535 10319 9561
rect 10345 9535 10351 9561
rect 10761 9535 10767 9561
rect 10793 9535 10799 9561
rect 7967 9529 7993 9535
rect 11495 9529 11521 9535
rect 8913 9479 8919 9505
rect 8945 9479 8951 9505
rect 9417 9479 9423 9505
rect 9449 9479 9455 9505
rect 9977 9479 9983 9505
rect 10009 9479 10015 9505
rect 10817 9479 10823 9505
rect 10849 9479 10855 9505
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 9031 9337 9057 9343
rect 9031 9305 9057 9311
rect 10375 9337 10401 9343
rect 10375 9305 10401 9311
rect 8695 9281 8721 9287
rect 7233 9255 7239 9281
rect 7265 9255 7271 9281
rect 8695 9249 8721 9255
rect 8807 9281 8833 9287
rect 9983 9281 10009 9287
rect 9193 9255 9199 9281
rect 9225 9255 9231 9281
rect 8807 9249 8833 9255
rect 9983 9249 10009 9255
rect 10655 9281 10681 9287
rect 10655 9249 10681 9255
rect 10711 9281 10737 9287
rect 10711 9249 10737 9255
rect 8751 9225 8777 9231
rect 2137 9199 2143 9225
rect 2169 9199 2175 9225
rect 6337 9199 6343 9225
rect 6369 9199 6375 9225
rect 6841 9199 6847 9225
rect 6873 9199 6879 9225
rect 8751 9193 8777 9199
rect 10151 9225 10177 9231
rect 10151 9193 10177 9199
rect 10207 9225 10233 9231
rect 10823 9225 10849 9231
rect 10313 9199 10319 9225
rect 10345 9199 10351 9225
rect 10207 9193 10233 9199
rect 10823 9193 10849 9199
rect 10935 9225 10961 9231
rect 10935 9193 10961 9199
rect 10991 9225 11017 9231
rect 10991 9193 11017 9199
rect 11215 9225 11241 9231
rect 11215 9193 11241 9199
rect 11327 9225 11353 9231
rect 18825 9199 18831 9225
rect 18857 9199 18863 9225
rect 11327 9193 11353 9199
rect 4881 9143 4887 9169
rect 4913 9143 4919 9169
rect 5945 9143 5951 9169
rect 5977 9143 5983 9169
rect 8297 9143 8303 9169
rect 8329 9143 8335 9169
rect 11097 9143 11103 9169
rect 11129 9143 11135 9169
rect 967 9113 993 9119
rect 967 9081 993 9087
rect 20007 9113 20033 9119
rect 20007 9081 20033 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 5783 8945 5809 8951
rect 5783 8913 5809 8919
rect 5727 8889 5753 8895
rect 6841 8863 6847 8889
rect 6873 8863 6879 8889
rect 9697 8863 9703 8889
rect 9729 8863 9735 8889
rect 11881 8863 11887 8889
rect 11913 8863 11919 8889
rect 12945 8863 12951 8889
rect 12977 8863 12983 8889
rect 5727 8857 5753 8863
rect 6791 8833 6817 8839
rect 6791 8801 6817 8807
rect 6959 8833 6985 8839
rect 7065 8807 7071 8833
rect 7097 8807 7103 8833
rect 9641 8807 9647 8833
rect 9673 8807 9679 8833
rect 11545 8807 11551 8833
rect 11577 8807 11583 8833
rect 6959 8801 6985 8807
rect 6847 8777 6873 8783
rect 6847 8745 6873 8751
rect 9815 8777 9841 8783
rect 10817 8751 10823 8777
rect 10849 8751 10855 8777
rect 10985 8751 10991 8777
rect 11017 8751 11023 8777
rect 9815 8745 9841 8751
rect 10655 8721 10681 8727
rect 10655 8689 10681 8695
rect 11159 8721 11185 8727
rect 11159 8689 11185 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 6679 8553 6705 8559
rect 6679 8521 6705 8527
rect 6959 8497 6985 8503
rect 10593 8471 10599 8497
rect 10625 8471 10631 8497
rect 6959 8465 6985 8471
rect 6735 8441 6761 8447
rect 6735 8409 6761 8415
rect 6847 8441 6873 8447
rect 11489 8415 11495 8441
rect 11521 8415 11527 8441
rect 6847 8409 6873 8415
rect 6791 8385 6817 8391
rect 6791 8353 6817 8359
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 10655 8161 10681 8167
rect 10655 8129 10681 8135
rect 11439 8161 11465 8167
rect 11439 8129 11465 8135
rect 967 8105 993 8111
rect 967 8073 993 8079
rect 6287 8105 6313 8111
rect 6287 8073 6313 8079
rect 9927 8105 9953 8111
rect 9927 8073 9953 8079
rect 9311 8049 9337 8055
rect 11271 8049 11297 8055
rect 2137 8023 2143 8049
rect 2169 8023 2175 8049
rect 6785 8023 6791 8049
rect 6817 8023 6823 8049
rect 7121 8023 7127 8049
rect 7153 8023 7159 8049
rect 9081 8023 9087 8049
rect 9113 8023 9119 8049
rect 9417 8023 9423 8049
rect 9449 8023 9455 8049
rect 11153 8023 11159 8049
rect 11185 8023 11191 8049
rect 9311 8017 9337 8023
rect 11271 8017 11297 8023
rect 9871 7993 9897 7999
rect 9871 7961 9897 7967
rect 9983 7993 10009 7999
rect 10375 7993 10401 7999
rect 10201 7967 10207 7993
rect 10233 7967 10239 7993
rect 9983 7961 10009 7967
rect 10375 7961 10401 7967
rect 10711 7993 10737 7999
rect 10711 7961 10737 7967
rect 11495 7993 11521 7999
rect 11495 7961 11521 7967
rect 6343 7937 6369 7943
rect 6343 7905 6369 7911
rect 6903 7937 6929 7943
rect 6903 7905 6929 7911
rect 6959 7937 6985 7943
rect 6959 7905 6985 7911
rect 7015 7937 7041 7943
rect 7015 7905 7041 7911
rect 9199 7937 9225 7943
rect 9199 7905 9225 7911
rect 9255 7937 9281 7943
rect 9255 7905 9281 7911
rect 11215 7937 11241 7943
rect 11215 7905 11241 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 8751 7769 8777 7775
rect 8751 7737 8777 7743
rect 8919 7769 8945 7775
rect 8919 7737 8945 7743
rect 10095 7769 10121 7775
rect 10095 7737 10121 7743
rect 8303 7713 8329 7719
rect 8303 7681 8329 7687
rect 9031 7713 9057 7719
rect 9031 7681 9057 7687
rect 9479 7713 9505 7719
rect 9479 7681 9505 7687
rect 10207 7713 10233 7719
rect 11265 7687 11271 7713
rect 11297 7687 11303 7713
rect 10207 7681 10233 7687
rect 8415 7657 8441 7663
rect 2137 7631 2143 7657
rect 2169 7631 2175 7657
rect 7065 7631 7071 7657
rect 7097 7631 7103 7657
rect 8415 7625 8441 7631
rect 8807 7657 8833 7663
rect 8807 7625 8833 7631
rect 8863 7657 8889 7663
rect 8863 7625 8889 7631
rect 9591 7657 9617 7663
rect 10929 7631 10935 7657
rect 10961 7631 10967 7657
rect 9591 7625 9617 7631
rect 5609 7575 5615 7601
rect 5641 7575 5647 7601
rect 6673 7575 6679 7601
rect 6705 7575 6711 7601
rect 10089 7575 10095 7601
rect 10121 7575 10127 7601
rect 12329 7575 12335 7601
rect 12361 7575 12367 7601
rect 967 7545 993 7551
rect 967 7513 993 7519
rect 8247 7545 8273 7551
rect 8247 7513 8273 7519
rect 9759 7545 9785 7551
rect 9759 7513 9785 7519
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 6455 7377 6481 7383
rect 6455 7345 6481 7351
rect 6399 7321 6425 7327
rect 7793 7295 7799 7321
rect 7825 7295 7831 7321
rect 8857 7295 8863 7321
rect 8889 7295 8895 7321
rect 6399 7289 6425 7295
rect 9031 7265 9057 7271
rect 7457 7239 7463 7265
rect 7489 7239 7495 7265
rect 9031 7233 9057 7239
rect 9199 7265 9225 7271
rect 9199 7233 9225 7239
rect 9367 7265 9393 7271
rect 9983 7265 10009 7271
rect 9697 7239 9703 7265
rect 9729 7239 9735 7265
rect 9367 7233 9393 7239
rect 9983 7233 10009 7239
rect 9585 7183 9591 7209
rect 9617 7183 9623 7209
rect 9199 7153 9225 7159
rect 9199 7121 9225 7127
rect 10151 7153 10177 7159
rect 10151 7121 10177 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 9423 6985 9449 6991
rect 9423 6953 9449 6959
rect 9535 6929 9561 6935
rect 6561 6903 6567 6929
rect 6593 6903 6599 6929
rect 9535 6897 9561 6903
rect 9591 6929 9617 6935
rect 10257 6903 10263 6929
rect 10289 6903 10295 6929
rect 9591 6897 9617 6903
rect 6953 6847 6959 6873
rect 6985 6847 6991 6873
rect 9865 6847 9871 6873
rect 9897 6847 9903 6873
rect 5497 6791 5503 6817
rect 5529 6791 5535 6817
rect 11321 6791 11327 6817
rect 11353 6791 11359 6817
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 8409 6511 8415 6537
rect 8441 6511 8447 6537
rect 9473 6511 9479 6537
rect 9505 6511 9511 6537
rect 8073 6455 8079 6481
rect 8105 6455 8111 6481
rect 9647 6369 9673 6375
rect 9809 6343 9815 6369
rect 9841 6343 9847 6369
rect 9647 6337 9673 6343
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 9473 6119 9479 6145
rect 9505 6119 9511 6145
rect 9361 6063 9367 6089
rect 9393 6063 9399 6089
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 20119 5361 20145 5367
rect 20119 5329 20145 5335
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 9367 2617 9393 2623
rect 9367 2585 9393 2591
rect 8857 2535 8863 2561
rect 8889 2535 8895 2561
rect 20119 2449 20145 2455
rect 20119 2417 20145 2423
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 9367 2225 9393 2231
rect 9367 2193 9393 2199
rect 9529 2143 9535 2169
rect 9561 2143 9567 2169
rect 10039 2057 10065 2063
rect 10039 2025 10065 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 9081 1807 9087 1833
rect 9113 1807 9119 1833
rect 9865 1751 9871 1777
rect 9897 1751 9903 1777
rect 10369 1751 10375 1777
rect 10401 1751 10407 1777
rect 10879 1665 10905 1671
rect 10879 1633 10905 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9591 19111 9617 19137
rect 11047 19111 11073 19137
rect 13063 19111 13089 19137
rect 9871 18999 9897 19025
rect 10543 18999 10569 19025
rect 12615 18999 12641 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 9199 18719 9225 18745
rect 10711 18719 10737 18745
rect 13399 18719 13425 18745
rect 855 18663 881 18689
rect 8695 18607 8721 18633
rect 10431 18607 10457 18633
rect 12895 18607 12921 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 10375 13567 10401 13593
rect 8919 13511 8945 13537
rect 9311 13455 9337 13481
rect 10711 13455 10737 13481
rect 8415 13399 8441 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 10487 13231 10513 13257
rect 10767 13175 10793 13201
rect 6903 13119 6929 13145
rect 8863 13119 8889 13145
rect 10375 13119 10401 13145
rect 10543 13119 10569 13145
rect 10823 13119 10849 13145
rect 7239 13063 7265 13089
rect 8303 13063 8329 13089
rect 9199 13063 9225 13089
rect 10263 13063 10289 13089
rect 11047 13063 11073 13089
rect 10767 13007 10793 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 8191 12839 8217 12865
rect 10151 12839 10177 12865
rect 967 12783 993 12809
rect 12839 12783 12865 12809
rect 20007 12783 20033 12809
rect 2143 12727 2169 12753
rect 7855 12727 7881 12753
rect 9759 12727 9785 12753
rect 9927 12727 9953 12753
rect 10207 12727 10233 12753
rect 11327 12727 11353 12753
rect 18831 12727 18857 12753
rect 7911 12671 7937 12697
rect 8023 12671 8049 12697
rect 8135 12671 8161 12697
rect 11719 12671 11745 12697
rect 8191 12615 8217 12641
rect 9871 12615 9897 12641
rect 10151 12615 10177 12641
rect 11159 12615 11185 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 7351 12447 7377 12473
rect 12615 12447 12641 12473
rect 12951 12447 12977 12473
rect 13119 12447 13145 12473
rect 12783 12391 12809 12417
rect 7015 12335 7041 12361
rect 7239 12335 7265 12361
rect 7463 12335 7489 12361
rect 7575 12335 7601 12361
rect 9871 12335 9897 12361
rect 9927 12335 9953 12361
rect 9983 12335 10009 12361
rect 10039 12335 10065 12361
rect 10095 12335 10121 12361
rect 10935 12335 10961 12361
rect 18831 12335 18857 12361
rect 5615 12279 5641 12305
rect 6679 12279 6705 12305
rect 7407 12279 7433 12305
rect 10711 12279 10737 12305
rect 11271 12279 11297 12305
rect 12335 12279 12361 12305
rect 20007 12223 20033 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 6735 12055 6761 12081
rect 6791 11999 6817 12025
rect 7183 11999 7209 12025
rect 9927 11999 9953 12025
rect 11439 11999 11465 12025
rect 11887 11999 11913 12025
rect 8527 11943 8553 11969
rect 11327 11943 11353 11969
rect 11551 11943 11577 11969
rect 11663 11943 11689 11969
rect 11943 11943 11969 11969
rect 12055 11943 12081 11969
rect 12447 11943 12473 11969
rect 7631 11887 7657 11913
rect 8863 11887 8889 11913
rect 10655 11887 10681 11913
rect 10823 11887 10849 11913
rect 11831 11887 11857 11913
rect 12279 11887 12305 11913
rect 12335 11887 12361 11913
rect 7799 11831 7825 11857
rect 10151 11831 10177 11857
rect 10711 11831 10737 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 7743 11663 7769 11689
rect 11775 11663 11801 11689
rect 11887 11663 11913 11689
rect 6119 11551 6145 11577
rect 11383 11551 11409 11577
rect 11719 11551 11745 11577
rect 6455 11495 6481 11521
rect 7519 11495 7545 11521
rect 10263 11495 10289 11521
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 8807 11271 8833 11297
rect 11159 11271 11185 11297
rect 967 11215 993 11241
rect 4719 11215 4745 11241
rect 6399 11215 6425 11241
rect 8415 11215 8441 11241
rect 9535 11215 9561 11241
rect 11047 11215 11073 11241
rect 20007 11215 20033 11241
rect 2143 11159 2169 11185
rect 6119 11159 6145 11185
rect 7911 11159 7937 11185
rect 8471 11159 8497 11185
rect 8639 11159 8665 11185
rect 8975 11159 9001 11185
rect 9423 11159 9449 11185
rect 9647 11159 9673 11185
rect 9759 11159 9785 11185
rect 10039 11159 10065 11185
rect 10207 11159 10233 11185
rect 10319 11159 10345 11185
rect 11327 11159 11353 11185
rect 11439 11159 11465 11185
rect 11719 11159 11745 11185
rect 18831 11159 18857 11185
rect 5783 11103 5809 11129
rect 8135 11103 8161 11129
rect 9031 11103 9057 11129
rect 9927 11103 9953 11129
rect 10823 11103 10849 11129
rect 10879 11103 10905 11129
rect 7799 11047 7825 11073
rect 8191 11047 8217 11073
rect 8303 11047 8329 11073
rect 8751 11047 8777 11073
rect 9255 11047 9281 11073
rect 10375 11047 10401 11073
rect 10655 11047 10681 11073
rect 10767 11047 10793 11073
rect 11215 11047 11241 11073
rect 11607 11047 11633 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 6175 10879 6201 10905
rect 6287 10879 6313 10905
rect 6623 10879 6649 10905
rect 6679 10879 6705 10905
rect 7631 10879 7657 10905
rect 8415 10879 8441 10905
rect 8751 10879 8777 10905
rect 9927 10879 9953 10905
rect 5839 10823 5865 10849
rect 7407 10823 7433 10849
rect 8247 10823 8273 10849
rect 8975 10823 9001 10849
rect 9087 10823 9113 10849
rect 10375 10823 10401 10849
rect 13343 10823 13369 10849
rect 6399 10767 6425 10793
rect 6567 10767 6593 10793
rect 6903 10767 6929 10793
rect 7799 10767 7825 10793
rect 8695 10767 8721 10793
rect 9815 10767 9841 10793
rect 10543 10767 10569 10793
rect 10823 10767 10849 10793
rect 11047 10767 11073 10793
rect 11215 10767 11241 10793
rect 11439 10767 11465 10793
rect 11551 10767 11577 10793
rect 13175 10767 13201 10793
rect 18831 10767 18857 10793
rect 5783 10711 5809 10737
rect 5951 10711 5977 10737
rect 6343 10711 6369 10737
rect 7127 10711 7153 10737
rect 10319 10711 10345 10737
rect 11495 10711 11521 10737
rect 7295 10655 7321 10681
rect 11327 10655 11353 10681
rect 20007 10655 20033 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 9591 10487 9617 10513
rect 10319 10431 10345 10457
rect 10935 10431 10961 10457
rect 11271 10431 11297 10457
rect 12279 10431 12305 10457
rect 13343 10431 13369 10457
rect 6119 10375 6145 10401
rect 6231 10375 6257 10401
rect 6679 10375 6705 10401
rect 6847 10375 6873 10401
rect 9759 10375 9785 10401
rect 9871 10375 9897 10401
rect 10095 10375 10121 10401
rect 10263 10375 10289 10401
rect 10991 10375 11017 10401
rect 11159 10375 11185 10401
rect 11719 10375 11745 10401
rect 11887 10375 11913 10401
rect 6791 10319 6817 10345
rect 7911 10319 7937 10345
rect 8079 10319 8105 10345
rect 8695 10319 8721 10345
rect 8863 10319 8889 10345
rect 10767 10319 10793 10345
rect 6175 10263 6201 10289
rect 6343 10263 6369 10289
rect 8527 10263 8553 10289
rect 9031 10263 9057 10289
rect 9255 10263 9281 10289
rect 10375 10263 10401 10289
rect 10879 10263 10905 10289
rect 11271 10263 11297 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 6343 10095 6369 10121
rect 7351 10095 7377 10121
rect 7463 10095 7489 10121
rect 5839 10039 5865 10065
rect 6455 10039 6481 10065
rect 6735 10039 6761 10065
rect 8695 10039 8721 10065
rect 8751 10039 8777 10065
rect 9143 10039 9169 10065
rect 12671 10039 12697 10065
rect 12727 10039 12753 10065
rect 2143 9983 2169 10009
rect 6231 9983 6257 10009
rect 6511 9983 6537 10009
rect 7687 9983 7713 10009
rect 8863 9983 8889 10009
rect 8975 9983 9001 10009
rect 9311 9983 9337 10009
rect 4775 9927 4801 9953
rect 7407 9927 7433 9953
rect 9087 9927 9113 9953
rect 11719 9927 11745 9953
rect 967 9871 993 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 8023 9703 8049 9729
rect 8247 9703 8273 9729
rect 8415 9647 8441 9673
rect 11607 9647 11633 9673
rect 12223 9647 12249 9673
rect 13287 9647 13313 9673
rect 20007 9647 20033 9673
rect 7351 9591 7377 9617
rect 8471 9591 8497 9617
rect 8807 9591 8833 9617
rect 9311 9591 9337 9617
rect 9815 9591 9841 9617
rect 10599 9591 10625 9617
rect 10879 9591 10905 9617
rect 10991 9591 11017 9617
rect 11103 9591 11129 9617
rect 11663 9591 11689 9617
rect 11831 9591 11857 9617
rect 18831 9591 18857 9617
rect 7183 9535 7209 9561
rect 7967 9535 7993 9561
rect 10039 9535 10065 9561
rect 10319 9535 10345 9561
rect 10767 9535 10793 9561
rect 11495 9535 11521 9561
rect 8919 9479 8945 9505
rect 9423 9479 9449 9505
rect 9983 9479 10009 9505
rect 10823 9479 10849 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 9031 9311 9057 9337
rect 10375 9311 10401 9337
rect 7239 9255 7265 9281
rect 8695 9255 8721 9281
rect 8807 9255 8833 9281
rect 9199 9255 9225 9281
rect 9983 9255 10009 9281
rect 10655 9255 10681 9281
rect 10711 9255 10737 9281
rect 2143 9199 2169 9225
rect 6343 9199 6369 9225
rect 6847 9199 6873 9225
rect 8751 9199 8777 9225
rect 10151 9199 10177 9225
rect 10207 9199 10233 9225
rect 10319 9199 10345 9225
rect 10823 9199 10849 9225
rect 10935 9199 10961 9225
rect 10991 9199 11017 9225
rect 11215 9199 11241 9225
rect 11327 9199 11353 9225
rect 18831 9199 18857 9225
rect 4887 9143 4913 9169
rect 5951 9143 5977 9169
rect 8303 9143 8329 9169
rect 11103 9143 11129 9169
rect 967 9087 993 9113
rect 20007 9087 20033 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 5783 8919 5809 8945
rect 5727 8863 5753 8889
rect 6847 8863 6873 8889
rect 9703 8863 9729 8889
rect 11887 8863 11913 8889
rect 12951 8863 12977 8889
rect 6791 8807 6817 8833
rect 6959 8807 6985 8833
rect 7071 8807 7097 8833
rect 9647 8807 9673 8833
rect 11551 8807 11577 8833
rect 6847 8751 6873 8777
rect 9815 8751 9841 8777
rect 10823 8751 10849 8777
rect 10991 8751 11017 8777
rect 10655 8695 10681 8721
rect 11159 8695 11185 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 6679 8527 6705 8553
rect 6959 8471 6985 8497
rect 10599 8471 10625 8497
rect 6735 8415 6761 8441
rect 6847 8415 6873 8441
rect 11495 8415 11521 8441
rect 6791 8359 6817 8385
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 10655 8135 10681 8161
rect 11439 8135 11465 8161
rect 967 8079 993 8105
rect 6287 8079 6313 8105
rect 9927 8079 9953 8105
rect 2143 8023 2169 8049
rect 6791 8023 6817 8049
rect 7127 8023 7153 8049
rect 9087 8023 9113 8049
rect 9311 8023 9337 8049
rect 9423 8023 9449 8049
rect 11159 8023 11185 8049
rect 11271 8023 11297 8049
rect 9871 7967 9897 7993
rect 9983 7967 10009 7993
rect 10207 7967 10233 7993
rect 10375 7967 10401 7993
rect 10711 7967 10737 7993
rect 11495 7967 11521 7993
rect 6343 7911 6369 7937
rect 6903 7911 6929 7937
rect 6959 7911 6985 7937
rect 7015 7911 7041 7937
rect 9199 7911 9225 7937
rect 9255 7911 9281 7937
rect 11215 7911 11241 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 8751 7743 8777 7769
rect 8919 7743 8945 7769
rect 10095 7743 10121 7769
rect 8303 7687 8329 7713
rect 9031 7687 9057 7713
rect 9479 7687 9505 7713
rect 10207 7687 10233 7713
rect 11271 7687 11297 7713
rect 2143 7631 2169 7657
rect 7071 7631 7097 7657
rect 8415 7631 8441 7657
rect 8807 7631 8833 7657
rect 8863 7631 8889 7657
rect 9591 7631 9617 7657
rect 10935 7631 10961 7657
rect 5615 7575 5641 7601
rect 6679 7575 6705 7601
rect 10095 7575 10121 7601
rect 12335 7575 12361 7601
rect 967 7519 993 7545
rect 8247 7519 8273 7545
rect 9759 7519 9785 7545
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 6455 7351 6481 7377
rect 6399 7295 6425 7321
rect 7799 7295 7825 7321
rect 8863 7295 8889 7321
rect 7463 7239 7489 7265
rect 9031 7239 9057 7265
rect 9199 7239 9225 7265
rect 9367 7239 9393 7265
rect 9703 7239 9729 7265
rect 9983 7239 10009 7265
rect 9591 7183 9617 7209
rect 9199 7127 9225 7153
rect 10151 7127 10177 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 9423 6959 9449 6985
rect 6567 6903 6593 6929
rect 9535 6903 9561 6929
rect 9591 6903 9617 6929
rect 10263 6903 10289 6929
rect 6959 6847 6985 6873
rect 9871 6847 9897 6873
rect 5503 6791 5529 6817
rect 11327 6791 11353 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 8415 6511 8441 6537
rect 9479 6511 9505 6537
rect 8079 6455 8105 6481
rect 9647 6343 9673 6369
rect 9815 6343 9841 6369
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 9479 6119 9505 6145
rect 9367 6063 9393 6089
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 20119 5335 20145 5361
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9367 2591 9393 2617
rect 8863 2535 8889 2561
rect 20119 2423 20145 2449
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 9367 2199 9393 2225
rect 9535 2143 9561 2169
rect 10039 2031 10065 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 9087 1807 9113 1833
rect 9871 1751 9897 1777
rect 10375 1751 10401 1777
rect 10879 1639 10905 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8064 20600 8120 21000
rect 9744 20600 9800 21000
rect 10080 20600 10136 21000
rect 10416 20600 10472 21000
rect 12432 20600 12488 21000
rect 12768 20600 12824 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 8078 18746 8106 20600
rect 9590 19138 9618 19143
rect 9758 19138 9786 20600
rect 9590 19137 9786 19138
rect 9590 19111 9591 19137
rect 9617 19111 9786 19137
rect 9590 19110 9786 19111
rect 9590 19105 9618 19110
rect 9870 19026 9898 19031
rect 9646 19025 9898 19026
rect 9646 18999 9871 19025
rect 9897 18999 9898 19025
rect 9646 18998 9898 18999
rect 8078 18713 8106 18718
rect 9198 18746 9226 18751
rect 9198 18699 9226 18718
rect 854 18689 882 18695
rect 854 18663 855 18689
rect 881 18663 882 18689
rect 854 18522 882 18663
rect 854 18489 882 18494
rect 8694 18633 8722 18639
rect 8694 18607 8695 18633
rect 8721 18607 8722 18633
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 8414 13425 8442 13431
rect 8414 13399 8415 13425
rect 8441 13399 8442 13425
rect 2478 13146 2506 13151
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 966 12809 994 12815
rect 966 12783 967 12809
rect 993 12783 994 12809
rect 966 12474 994 12783
rect 966 12441 994 12446
rect 2142 12753 2170 12759
rect 2142 12727 2143 12753
rect 2169 12727 2170 12753
rect 2142 12306 2170 12727
rect 2142 12273 2170 12278
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 966 11242 994 11247
rect 966 11195 994 11214
rect 2142 11186 2170 11191
rect 2142 11139 2170 11158
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 2478 10290 2506 13118
rect 6902 13146 6930 13151
rect 7854 13146 7882 13151
rect 6902 13145 7042 13146
rect 6902 13119 6903 13145
rect 6929 13119 7042 13145
rect 6902 13118 7042 13119
rect 6902 13113 6930 13118
rect 7014 12362 7042 13118
rect 7238 13090 7266 13095
rect 7238 13043 7266 13062
rect 7854 12753 7882 13118
rect 8190 13090 8218 13095
rect 7854 12727 7855 12753
rect 7881 12727 7882 12753
rect 7350 12474 7378 12479
rect 7350 12427 7378 12446
rect 7630 12474 7658 12479
rect 7014 12361 7210 12362
rect 7014 12335 7015 12361
rect 7041 12335 7210 12361
rect 7014 12334 7210 12335
rect 7014 12329 7042 12334
rect 5614 12306 5642 12311
rect 5614 12259 5642 12278
rect 6678 12306 6706 12311
rect 6678 12305 6762 12306
rect 6678 12279 6679 12305
rect 6705 12279 6762 12305
rect 6678 12278 6762 12279
rect 6678 12273 6706 12278
rect 6734 12081 6762 12278
rect 6734 12055 6735 12081
rect 6761 12055 6762 12081
rect 6734 12049 6762 12055
rect 6790 12026 6818 12031
rect 6790 11979 6818 11998
rect 7182 12025 7210 12334
rect 7238 12361 7266 12367
rect 7238 12335 7239 12361
rect 7265 12335 7266 12361
rect 7238 12306 7266 12335
rect 7462 12361 7490 12367
rect 7462 12335 7463 12361
rect 7489 12335 7490 12361
rect 7238 12273 7266 12278
rect 7406 12305 7434 12311
rect 7406 12279 7407 12305
rect 7433 12279 7434 12305
rect 7182 11999 7183 12025
rect 7209 11999 7210 12025
rect 7182 11802 7210 11999
rect 7406 12026 7434 12279
rect 7406 11993 7434 11998
rect 7182 11769 7210 11774
rect 6118 11690 6146 11695
rect 6118 11577 6146 11662
rect 6118 11551 6119 11577
rect 6145 11551 6146 11577
rect 4718 11241 4746 11247
rect 4718 11215 4719 11241
rect 4745 11215 4746 11241
rect 4718 11186 4746 11215
rect 4718 11153 4746 11158
rect 6118 11185 6146 11551
rect 6398 11690 6426 11695
rect 6398 11242 6426 11662
rect 6454 11522 6482 11527
rect 6454 11521 6650 11522
rect 6454 11495 6455 11521
rect 6481 11495 6650 11521
rect 6454 11494 6650 11495
rect 6454 11489 6482 11494
rect 6398 11241 6538 11242
rect 6398 11215 6399 11241
rect 6425 11215 6538 11241
rect 6398 11214 6538 11215
rect 6398 11209 6426 11214
rect 6118 11159 6119 11185
rect 6145 11159 6146 11185
rect 6118 11153 6146 11159
rect 6286 11186 6314 11191
rect 5782 11129 5810 11135
rect 5782 11103 5783 11129
rect 5809 11103 5810 11129
rect 5782 10737 5810 11103
rect 6174 10906 6202 10911
rect 5782 10711 5783 10737
rect 5809 10711 5810 10737
rect 5782 10705 5810 10711
rect 5838 10849 5866 10855
rect 5838 10823 5839 10849
rect 5865 10823 5866 10849
rect 5838 10626 5866 10823
rect 5950 10738 5978 10743
rect 5950 10691 5978 10710
rect 5838 10593 5866 10598
rect 6118 10402 6146 10407
rect 6174 10402 6202 10878
rect 6286 10905 6314 11158
rect 6286 10879 6287 10905
rect 6313 10879 6314 10905
rect 6286 10873 6314 10879
rect 6398 10794 6426 10799
rect 6398 10747 6426 10766
rect 6342 10738 6370 10743
rect 6342 10691 6370 10710
rect 6510 10570 6538 11214
rect 6622 10905 6650 11494
rect 7462 10962 7490 12335
rect 7574 12362 7602 12367
rect 7574 12315 7602 12334
rect 7630 11913 7658 12446
rect 7854 12474 7882 12727
rect 7910 13034 7938 13039
rect 7910 12697 7938 13006
rect 8190 12865 8218 13062
rect 8302 13090 8330 13095
rect 8302 13043 8330 13062
rect 8190 12839 8191 12865
rect 8217 12839 8218 12865
rect 8190 12833 8218 12839
rect 7910 12671 7911 12697
rect 7937 12671 7938 12697
rect 7910 12665 7938 12671
rect 8022 12698 8050 12703
rect 8134 12698 8162 12703
rect 8022 12697 8162 12698
rect 8022 12671 8023 12697
rect 8049 12671 8135 12697
rect 8161 12671 8162 12697
rect 8022 12670 8162 12671
rect 8022 12665 8050 12670
rect 8134 12665 8162 12670
rect 7854 12441 7882 12446
rect 8190 12641 8218 12647
rect 8190 12615 8191 12641
rect 8217 12615 8218 12641
rect 7630 11887 7631 11913
rect 7657 11887 7658 11913
rect 7630 11881 7658 11887
rect 7798 11857 7826 11863
rect 7798 11831 7799 11857
rect 7825 11831 7826 11857
rect 7742 11690 7770 11695
rect 7742 11643 7770 11662
rect 7518 11522 7546 11527
rect 7518 11475 7546 11494
rect 7798 11298 7826 11831
rect 8190 11802 8218 12615
rect 8414 11970 8442 13399
rect 8694 13090 8722 18607
rect 8918 13537 8946 13543
rect 8918 13511 8919 13537
rect 8945 13511 8946 13537
rect 8862 13146 8890 13151
rect 8918 13146 8946 13511
rect 8862 13145 8946 13146
rect 8862 13119 8863 13145
rect 8889 13119 8946 13145
rect 8862 13118 8946 13119
rect 8862 13113 8890 13118
rect 8694 13057 8722 13062
rect 8526 11970 8554 11975
rect 8414 11942 8526 11970
rect 8526 11923 8554 11942
rect 8918 11970 8946 13118
rect 9310 13481 9338 13487
rect 9310 13455 9311 13481
rect 9337 13455 9338 13481
rect 9198 13090 9226 13095
rect 9198 13043 9226 13062
rect 9310 12922 9338 13455
rect 9310 12889 9338 12894
rect 9646 12418 9674 18998
rect 9870 18993 9898 18998
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 10094 18746 10122 20600
rect 10430 19138 10458 20600
rect 10430 19105 10458 19110
rect 11046 19138 11074 19143
rect 11046 19091 11074 19110
rect 12446 19138 12474 20600
rect 12446 19105 12474 19110
rect 10542 19026 10570 19031
rect 10094 18713 10122 18718
rect 10374 19025 10570 19026
rect 10374 18999 10543 19025
rect 10569 18999 10570 19025
rect 10374 18998 10570 18999
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 10374 13594 10402 18998
rect 10542 18993 10570 18998
rect 12614 19025 12642 19031
rect 12614 18999 12615 19025
rect 12641 18999 12642 19025
rect 10710 18746 10738 18751
rect 10710 18699 10738 18718
rect 10430 18633 10458 18639
rect 10430 18607 10431 18633
rect 10457 18607 10458 18633
rect 10430 17290 10458 18607
rect 10430 17262 10626 17290
rect 10598 15974 10626 17262
rect 10598 15946 10794 15974
rect 10374 13593 10514 13594
rect 10374 13567 10375 13593
rect 10401 13567 10514 13593
rect 10374 13566 10514 13567
rect 10374 13561 10402 13566
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 10486 13257 10514 13566
rect 10486 13231 10487 13257
rect 10513 13231 10514 13257
rect 10486 13225 10514 13231
rect 10710 13481 10738 13487
rect 10710 13455 10711 13481
rect 10737 13455 10738 13481
rect 10262 13202 10290 13207
rect 9758 13090 9786 13095
rect 9758 12753 9786 13062
rect 10262 13089 10290 13174
rect 10374 13146 10402 13151
rect 10262 13063 10263 13089
rect 10289 13063 10290 13089
rect 10262 13057 10290 13063
rect 10318 13145 10402 13146
rect 10318 13119 10375 13145
rect 10401 13119 10402 13145
rect 10318 13118 10402 13119
rect 9758 12727 9759 12753
rect 9785 12727 9786 12753
rect 9758 12721 9786 12727
rect 9926 13034 9954 13039
rect 9926 12753 9954 13006
rect 10094 12922 10122 12927
rect 10122 12894 10178 12922
rect 10094 12889 10122 12894
rect 10150 12865 10178 12894
rect 10150 12839 10151 12865
rect 10177 12839 10178 12865
rect 10150 12833 10178 12839
rect 9926 12727 9927 12753
rect 9953 12727 9954 12753
rect 9926 12721 9954 12727
rect 10206 12754 10234 12759
rect 10318 12754 10346 13118
rect 10374 13113 10402 13118
rect 10542 13146 10570 13151
rect 10542 13099 10570 13118
rect 10206 12753 10346 12754
rect 10206 12727 10207 12753
rect 10233 12727 10346 12753
rect 10206 12726 10346 12727
rect 10206 12721 10234 12726
rect 9870 12642 9898 12647
rect 9814 12641 9898 12642
rect 9814 12615 9871 12641
rect 9897 12615 9898 12641
rect 9814 12614 9898 12615
rect 9814 12586 9842 12614
rect 9870 12609 9898 12614
rect 10150 12642 10178 12647
rect 10150 12641 10234 12642
rect 10150 12615 10151 12641
rect 10177 12615 10234 12641
rect 10150 12614 10234 12615
rect 10150 12609 10178 12614
rect 9814 12553 9842 12558
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9646 12385 9674 12390
rect 10094 12418 10122 12423
rect 8862 11913 8890 11919
rect 8862 11887 8863 11913
rect 8889 11887 8890 11913
rect 8190 11769 8218 11774
rect 8638 11802 8666 11807
rect 8666 11774 8722 11802
rect 8638 11769 8666 11774
rect 7798 11265 7826 11270
rect 7910 11522 7938 11527
rect 7910 11242 7938 11494
rect 7910 11185 7938 11214
rect 8414 11242 8442 11247
rect 8414 11195 8442 11214
rect 7910 11159 7911 11185
rect 7937 11159 7938 11185
rect 7910 11153 7938 11159
rect 8470 11186 8498 11191
rect 8638 11186 8666 11191
rect 8470 11185 8638 11186
rect 8470 11159 8471 11185
rect 8497 11159 8638 11185
rect 8470 11158 8638 11159
rect 8134 11129 8162 11135
rect 8134 11103 8135 11129
rect 8161 11103 8162 11129
rect 7798 11073 7826 11079
rect 7798 11047 7799 11073
rect 7825 11047 7826 11073
rect 7462 10934 7546 10962
rect 6622 10879 6623 10905
rect 6649 10879 6650 10905
rect 6622 10873 6650 10879
rect 6678 10906 6706 10911
rect 6678 10859 6706 10878
rect 7406 10850 7434 10855
rect 7406 10803 7434 10822
rect 6566 10793 6594 10799
rect 6566 10767 6567 10793
rect 6593 10767 6594 10793
rect 6566 10626 6594 10767
rect 6790 10794 6818 10799
rect 6566 10598 6706 10626
rect 6510 10542 6650 10570
rect 6230 10402 6258 10407
rect 6174 10401 6258 10402
rect 6174 10375 6231 10401
rect 6257 10375 6258 10401
rect 6174 10374 6258 10375
rect 6118 10355 6146 10374
rect 6230 10369 6258 10374
rect 2478 10257 2506 10262
rect 6174 10289 6202 10295
rect 6174 10263 6175 10289
rect 6201 10263 6202 10289
rect 6174 10122 6202 10263
rect 5838 10094 6202 10122
rect 6342 10289 6370 10295
rect 6342 10263 6343 10289
rect 6369 10263 6370 10289
rect 6342 10121 6370 10263
rect 6622 10178 6650 10542
rect 6678 10402 6706 10598
rect 6678 10355 6706 10374
rect 6790 10346 6818 10766
rect 6902 10794 6930 10799
rect 6902 10793 7154 10794
rect 6902 10767 6903 10793
rect 6929 10767 7154 10793
rect 6902 10766 7154 10767
rect 6902 10761 6930 10766
rect 7126 10737 7154 10766
rect 7126 10711 7127 10737
rect 7153 10711 7154 10737
rect 7126 10705 7154 10711
rect 7294 10681 7322 10687
rect 7294 10655 7295 10681
rect 7321 10655 7322 10681
rect 6846 10514 6874 10519
rect 6846 10401 6874 10486
rect 7294 10514 7322 10655
rect 7322 10486 7378 10514
rect 7294 10481 7322 10486
rect 6846 10375 6847 10401
rect 6873 10375 6874 10401
rect 6846 10369 6874 10375
rect 6790 10299 6818 10318
rect 6622 10150 6706 10178
rect 6342 10095 6343 10121
rect 6369 10095 6370 10121
rect 5838 10065 5866 10094
rect 6342 10089 6370 10095
rect 5838 10039 5839 10065
rect 5865 10039 5866 10065
rect 5838 10033 5866 10039
rect 6230 10066 6258 10071
rect 2142 10010 2170 10015
rect 2142 9963 2170 9982
rect 4774 10010 4802 10015
rect 4774 9953 4802 9982
rect 6230 10009 6258 10038
rect 6230 9983 6231 10009
rect 6257 9983 6258 10009
rect 6230 9977 6258 9983
rect 6454 10065 6482 10071
rect 6454 10039 6455 10065
rect 6481 10039 6482 10065
rect 6454 10010 6482 10039
rect 6678 10066 6706 10150
rect 7350 10121 7378 10486
rect 7350 10095 7351 10121
rect 7377 10095 7378 10121
rect 7350 10089 7378 10095
rect 7462 10346 7490 10351
rect 7462 10121 7490 10318
rect 7462 10095 7463 10121
rect 7489 10095 7490 10121
rect 7462 10089 7490 10095
rect 6734 10066 6762 10071
rect 6706 10065 6762 10066
rect 6706 10039 6735 10065
rect 6761 10039 6762 10065
rect 6706 10038 6762 10039
rect 6678 10019 6706 10038
rect 6734 10033 6762 10038
rect 6454 9977 6482 9982
rect 6510 10009 6538 10015
rect 6510 9983 6511 10009
rect 6537 9983 6538 10009
rect 4774 9927 4775 9953
rect 4801 9927 4802 9953
rect 4774 9921 4802 9927
rect 966 9898 994 9903
rect 966 9851 994 9870
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 6510 9562 6538 9983
rect 7406 9953 7434 9959
rect 7406 9927 7407 9953
rect 7433 9927 7434 9953
rect 7350 9842 7378 9847
rect 6958 9674 6986 9679
rect 6510 9529 6538 9534
rect 6790 9562 6818 9567
rect 2142 9226 2170 9231
rect 2142 9179 2170 9198
rect 4886 9226 4914 9231
rect 4886 9169 4914 9198
rect 6342 9226 6370 9231
rect 6342 9179 6370 9198
rect 5950 9170 5978 9175
rect 4886 9143 4887 9169
rect 4913 9143 4914 9169
rect 966 9114 994 9119
rect 966 9067 994 9086
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 4886 8778 4914 9143
rect 5782 9169 5978 9170
rect 5782 9143 5951 9169
rect 5977 9143 5978 9169
rect 5782 9142 5978 9143
rect 5782 8945 5810 9142
rect 5950 9137 5978 9142
rect 5782 8919 5783 8945
rect 5809 8919 5810 8945
rect 5782 8913 5810 8919
rect 5726 8890 5754 8895
rect 5726 8843 5754 8862
rect 6790 8834 6818 9534
rect 6846 9226 6874 9231
rect 6846 9179 6874 9198
rect 6846 8890 6874 8895
rect 6846 8843 6874 8862
rect 4886 8745 4914 8750
rect 6678 8833 6818 8834
rect 6678 8807 6791 8833
rect 6817 8807 6818 8833
rect 6678 8806 6818 8807
rect 6678 8554 6706 8806
rect 6790 8801 6818 8806
rect 6958 8833 6986 9646
rect 7350 9617 7378 9814
rect 7350 9591 7351 9617
rect 7377 9591 7378 9617
rect 7350 9585 7378 9591
rect 7182 9562 7210 9567
rect 7182 9515 7210 9534
rect 7406 9506 7434 9927
rect 7238 9478 7434 9506
rect 7238 9281 7266 9478
rect 7238 9255 7239 9281
rect 7265 9255 7266 9281
rect 7238 9249 7266 9255
rect 6958 8807 6959 8833
rect 6985 8807 6986 8833
rect 6846 8778 6874 8783
rect 6846 8731 6874 8750
rect 6622 8553 6706 8554
rect 6622 8527 6679 8553
rect 6705 8527 6706 8553
rect 6622 8526 6706 8527
rect 6286 8386 6314 8391
rect 5502 8330 5530 8335
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 966 8105 994 8111
rect 966 8079 967 8105
rect 993 8079 994 8105
rect 966 7770 994 8079
rect 2142 8050 2170 8055
rect 2142 8003 2170 8022
rect 966 7737 994 7742
rect 2142 7658 2170 7663
rect 2142 7611 2170 7630
rect 5502 7658 5530 8302
rect 6286 8105 6314 8358
rect 6622 8162 6650 8526
rect 6678 8521 6706 8526
rect 6958 8497 6986 8807
rect 6958 8471 6959 8497
rect 6985 8471 6986 8497
rect 6958 8465 6986 8471
rect 7014 9226 7042 9231
rect 6734 8441 6762 8447
rect 6734 8415 6735 8441
rect 6761 8415 6762 8441
rect 6734 8330 6762 8415
rect 6846 8441 6874 8447
rect 6846 8415 6847 8441
rect 6873 8415 6874 8441
rect 6790 8386 6818 8391
rect 6790 8339 6818 8358
rect 6734 8297 6762 8302
rect 6622 8134 6818 8162
rect 6286 8079 6287 8105
rect 6313 8079 6314 8105
rect 6286 8073 6314 8079
rect 966 7546 994 7551
rect 966 7499 994 7518
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 5502 6817 5530 7630
rect 5614 8050 5642 8055
rect 5614 7882 5642 8022
rect 6790 8049 6818 8134
rect 6790 8023 6791 8049
rect 6817 8023 6818 8049
rect 6790 8017 6818 8023
rect 6846 8050 6874 8415
rect 7014 8442 7042 9198
rect 7126 9170 7154 9175
rect 7070 9002 7098 9007
rect 7070 8833 7098 8974
rect 7070 8807 7071 8833
rect 7097 8807 7098 8833
rect 7070 8801 7098 8807
rect 7014 8414 7098 8442
rect 6846 8022 7042 8050
rect 5614 7601 5642 7854
rect 5614 7575 5615 7601
rect 5641 7575 5642 7601
rect 5614 7569 5642 7575
rect 6342 7937 6370 7943
rect 6342 7911 6343 7937
rect 6369 7911 6370 7937
rect 6342 7098 6370 7911
rect 6398 7938 6426 7943
rect 6398 7321 6426 7910
rect 6902 7937 6930 7943
rect 6902 7911 6903 7937
rect 6929 7911 6930 7937
rect 6902 7882 6930 7911
rect 6958 7938 6986 7943
rect 6958 7891 6986 7910
rect 7014 7937 7042 8022
rect 7014 7911 7015 7937
rect 7041 7911 7042 7937
rect 6902 7849 6930 7854
rect 7014 7770 7042 7911
rect 7014 7737 7042 7742
rect 7070 7657 7098 8414
rect 7126 8049 7154 9142
rect 7518 9002 7546 10934
rect 7630 10906 7658 10911
rect 7630 10859 7658 10878
rect 7798 10794 7826 11047
rect 8134 10906 8162 11103
rect 8134 10873 8162 10878
rect 8190 11073 8218 11079
rect 8190 11047 8191 11073
rect 8217 11047 8218 11073
rect 7798 10747 7826 10766
rect 8190 10570 8218 11047
rect 8302 11074 8330 11079
rect 8302 11027 8330 11046
rect 8470 11018 8498 11158
rect 8638 11139 8666 11158
rect 8414 10990 8498 11018
rect 8414 10905 8442 10990
rect 8414 10879 8415 10905
rect 8441 10879 8442 10905
rect 8414 10873 8442 10879
rect 8638 10962 8666 10967
rect 8246 10850 8274 10855
rect 8246 10803 8274 10822
rect 7910 10542 8218 10570
rect 8414 10794 8442 10799
rect 7910 10346 7938 10542
rect 8078 10346 8106 10351
rect 7910 10299 7938 10318
rect 8022 10318 8078 10346
rect 7686 10066 7714 10071
rect 7686 10009 7714 10038
rect 7686 9983 7687 10009
rect 7713 9983 7714 10009
rect 7686 9977 7714 9983
rect 8022 9730 8050 10318
rect 8078 10299 8106 10318
rect 8414 10290 8442 10766
rect 8526 10290 8554 10295
rect 8414 10289 8554 10290
rect 8414 10263 8527 10289
rect 8553 10263 8554 10289
rect 8414 10262 8554 10263
rect 7910 9729 8050 9730
rect 7910 9703 8023 9729
rect 8049 9703 8050 9729
rect 7910 9702 8050 9703
rect 7910 9226 7938 9702
rect 8022 9697 8050 9702
rect 8246 9729 8274 9735
rect 8246 9703 8247 9729
rect 8273 9703 8274 9729
rect 8246 9674 8274 9703
rect 8246 9641 8274 9646
rect 8414 9673 8442 10262
rect 8526 10257 8554 10262
rect 8638 9842 8666 10934
rect 8694 10906 8722 11774
rect 8862 11466 8890 11887
rect 8918 11690 8946 11942
rect 8918 11657 8946 11662
rect 9422 12362 9450 12367
rect 8862 11433 8890 11438
rect 8806 11298 8834 11303
rect 8806 11251 8834 11270
rect 8918 11298 8946 11303
rect 8750 11073 8778 11079
rect 8750 11047 8751 11073
rect 8777 11047 8778 11073
rect 8750 11018 8778 11047
rect 8750 10990 8834 11018
rect 8750 10906 8778 10911
rect 8694 10905 8778 10906
rect 8694 10879 8751 10905
rect 8777 10879 8778 10905
rect 8694 10878 8778 10879
rect 8694 10793 8722 10799
rect 8694 10767 8695 10793
rect 8721 10767 8722 10793
rect 8694 10514 8722 10767
rect 8694 10481 8722 10486
rect 8694 10402 8722 10407
rect 8694 10345 8722 10374
rect 8694 10319 8695 10345
rect 8721 10319 8722 10345
rect 8694 10313 8722 10319
rect 8750 10234 8778 10878
rect 8806 10850 8834 10990
rect 8918 10962 8946 11270
rect 8974 11186 9002 11191
rect 8974 11139 9002 11158
rect 9422 11185 9450 12334
rect 9870 12362 9898 12381
rect 9870 12329 9898 12334
rect 9926 12361 9954 12367
rect 9926 12335 9927 12361
rect 9953 12335 9954 12361
rect 9870 12250 9898 12255
rect 9814 12222 9870 12250
rect 9702 12026 9730 12031
rect 9534 11466 9562 11471
rect 9534 11241 9562 11438
rect 9534 11215 9535 11241
rect 9561 11215 9562 11241
rect 9534 11209 9562 11215
rect 9422 11159 9423 11185
rect 9449 11159 9450 11185
rect 8918 10929 8946 10934
rect 9030 11130 9058 11135
rect 8974 10850 9002 10855
rect 8806 10849 9002 10850
rect 8806 10823 8975 10849
rect 9001 10823 9002 10849
rect 8806 10822 9002 10823
rect 8974 10794 9002 10822
rect 8974 10761 9002 10766
rect 8694 10206 8778 10234
rect 8806 10458 8834 10463
rect 8694 10066 8722 10206
rect 8694 10033 8722 10038
rect 8750 10066 8778 10071
rect 8806 10066 8834 10430
rect 9030 10402 9058 11102
rect 9254 11073 9282 11079
rect 9254 11047 9255 11073
rect 9281 11047 9282 11073
rect 9142 10906 9170 10911
rect 8974 10374 9058 10402
rect 9086 10878 9142 10906
rect 9086 10849 9114 10878
rect 9142 10873 9170 10878
rect 9086 10823 9087 10849
rect 9113 10823 9114 10849
rect 9086 10402 9114 10823
rect 9198 10850 9226 10855
rect 8862 10346 8890 10351
rect 8862 10299 8890 10318
rect 8750 10065 8834 10066
rect 8750 10039 8751 10065
rect 8777 10039 8834 10065
rect 8750 10038 8834 10039
rect 8750 10033 8778 10038
rect 8862 10009 8890 10015
rect 8974 10010 9002 10374
rect 9086 10369 9114 10374
rect 9142 10794 9170 10799
rect 9030 10290 9058 10295
rect 9142 10290 9170 10766
rect 9030 10289 9170 10290
rect 9030 10263 9031 10289
rect 9057 10263 9170 10289
rect 9030 10262 9170 10263
rect 9198 10402 9226 10822
rect 9254 10458 9282 11047
rect 9254 10425 9282 10430
rect 9030 10257 9058 10262
rect 9142 10066 9170 10071
rect 9198 10066 9226 10374
rect 9254 10290 9282 10295
rect 9282 10262 9338 10290
rect 9254 10243 9282 10262
rect 9142 10065 9226 10066
rect 9142 10039 9143 10065
rect 9169 10039 9226 10065
rect 9142 10038 9226 10039
rect 9142 10033 9170 10038
rect 8862 9983 8863 10009
rect 8889 9983 8890 10009
rect 8694 9842 8722 9847
rect 8638 9814 8694 9842
rect 8694 9809 8722 9814
rect 8862 9730 8890 9983
rect 8862 9697 8890 9702
rect 8918 10009 9002 10010
rect 8918 9983 8975 10009
rect 9001 9983 9002 10009
rect 8918 9982 9002 9983
rect 8414 9647 8415 9673
rect 8441 9647 8442 9673
rect 8358 9618 8386 9623
rect 8302 9590 8358 9618
rect 7966 9562 7994 9567
rect 8302 9562 8330 9590
rect 8358 9585 8386 9590
rect 7966 9561 8330 9562
rect 7966 9535 7967 9561
rect 7993 9535 8330 9561
rect 7966 9534 8330 9535
rect 7966 9529 7994 9534
rect 7910 9193 7938 9198
rect 8302 9169 8330 9534
rect 8414 9506 8442 9647
rect 8470 9618 8498 9623
rect 8470 9571 8498 9590
rect 8806 9618 8834 9637
rect 8806 9585 8834 9590
rect 8806 9506 8834 9511
rect 8414 9478 8722 9506
rect 8694 9281 8722 9478
rect 8694 9255 8695 9281
rect 8721 9255 8722 9281
rect 8694 9249 8722 9255
rect 8750 9478 8806 9506
rect 8750 9225 8778 9478
rect 8806 9473 8834 9478
rect 8918 9505 8946 9982
rect 8974 9977 9002 9982
rect 9310 10009 9338 10262
rect 9310 9983 9311 10009
rect 9337 9983 9338 10009
rect 9310 9977 9338 9983
rect 9086 9953 9114 9959
rect 9086 9927 9087 9953
rect 9113 9927 9114 9953
rect 8918 9479 8919 9505
rect 8945 9479 8946 9505
rect 8750 9199 8751 9225
rect 8777 9199 8778 9225
rect 8750 9193 8778 9199
rect 8806 9281 8834 9287
rect 8806 9255 8807 9281
rect 8833 9255 8834 9281
rect 8806 9226 8834 9255
rect 8806 9193 8834 9198
rect 8918 9226 8946 9479
rect 9030 9618 9058 9623
rect 9030 9337 9058 9590
rect 9030 9311 9031 9337
rect 9057 9311 9058 9337
rect 9030 9305 9058 9311
rect 8918 9193 8946 9198
rect 8302 9143 8303 9169
rect 8329 9143 8330 9169
rect 8302 9137 8330 9143
rect 7518 8969 7546 8974
rect 8750 9114 8778 9119
rect 7126 8023 7127 8049
rect 7153 8023 7154 8049
rect 7126 8017 7154 8023
rect 8750 7769 8778 9086
rect 9086 8050 9114 9927
rect 9030 8049 9114 8050
rect 9030 8023 9087 8049
rect 9113 8023 9114 8049
rect 9030 8022 9114 8023
rect 8750 7743 8751 7769
rect 8777 7743 8778 7769
rect 7070 7631 7071 7657
rect 7097 7631 7098 7657
rect 6678 7601 6706 7607
rect 6678 7575 6679 7601
rect 6705 7575 6706 7601
rect 6678 7574 6706 7575
rect 6454 7546 6706 7574
rect 6454 7377 6482 7546
rect 6454 7351 6455 7377
rect 6481 7351 6482 7377
rect 6454 7345 6482 7351
rect 6398 7295 6399 7321
rect 6425 7295 6426 7321
rect 6398 7289 6426 7295
rect 7070 7266 7098 7631
rect 8302 7713 8330 7719
rect 8302 7687 8303 7713
rect 8329 7687 8330 7713
rect 8302 7602 8330 7687
rect 8414 7658 8442 7663
rect 8414 7611 8442 7630
rect 8302 7569 8330 7574
rect 8246 7546 8274 7551
rect 7798 7545 8274 7546
rect 7798 7519 8247 7545
rect 8273 7519 8274 7545
rect 7798 7518 8274 7519
rect 7798 7321 7826 7518
rect 8246 7513 8274 7518
rect 7798 7295 7799 7321
rect 7825 7295 7826 7321
rect 7798 7289 7826 7295
rect 7462 7266 7490 7271
rect 6958 7265 7490 7266
rect 6958 7239 7463 7265
rect 7489 7239 7490 7265
rect 6958 7238 7490 7239
rect 6342 7070 6594 7098
rect 6566 6929 6594 7070
rect 6566 6903 6567 6929
rect 6593 6903 6594 6929
rect 6566 6897 6594 6903
rect 6958 6873 6986 7238
rect 6958 6847 6959 6873
rect 6985 6847 6986 6873
rect 6958 6841 6986 6847
rect 5502 6791 5503 6817
rect 5529 6791 5530 6817
rect 5502 6785 5530 6791
rect 7462 6706 7490 7238
rect 8414 7154 8442 7159
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 7462 6673 7490 6678
rect 8078 6706 8106 6711
rect 2238 6645 2370 6650
rect 8078 6481 8106 6678
rect 8414 6537 8442 7126
rect 8750 7098 8778 7743
rect 8918 7770 8946 7775
rect 8918 7723 8946 7742
rect 9030 7713 9058 8022
rect 9086 8017 9114 8022
rect 9142 9730 9170 9735
rect 9030 7687 9031 7713
rect 9057 7687 9058 7713
rect 9030 7681 9058 7687
rect 8806 7657 8834 7663
rect 8806 7631 8807 7657
rect 8833 7631 8834 7657
rect 8806 7322 8834 7631
rect 8862 7658 8890 7663
rect 8862 7611 8890 7630
rect 9030 7602 9058 7607
rect 9142 7574 9170 9702
rect 9254 9674 9282 9679
rect 9198 9281 9226 9287
rect 9198 9255 9199 9281
rect 9225 9255 9226 9281
rect 9198 9114 9226 9255
rect 9198 9081 9226 9086
rect 9254 8050 9282 9646
rect 9310 9618 9338 9623
rect 9310 9571 9338 9590
rect 9422 9505 9450 11159
rect 9646 11186 9674 11191
rect 9590 10626 9618 10631
rect 9422 9479 9423 9505
rect 9449 9479 9450 9505
rect 9422 9170 9450 9479
rect 9534 10598 9590 10626
rect 9534 9226 9562 10598
rect 9590 10593 9618 10598
rect 9590 10514 9618 10519
rect 9590 10467 9618 10486
rect 9646 10402 9674 11158
rect 9702 10850 9730 11998
rect 9758 11186 9786 11191
rect 9814 11186 9842 12222
rect 9870 12217 9898 12222
rect 9926 12194 9954 12335
rect 9982 12362 10010 12367
rect 9982 12315 10010 12334
rect 10038 12361 10066 12367
rect 10038 12335 10039 12361
rect 10065 12335 10066 12361
rect 10038 12250 10066 12335
rect 9926 12161 9954 12166
rect 9982 12222 10066 12250
rect 10094 12361 10122 12390
rect 10094 12335 10095 12361
rect 10121 12335 10122 12361
rect 9926 12082 9954 12087
rect 9926 12025 9954 12054
rect 9926 11999 9927 12025
rect 9953 11999 9954 12025
rect 9926 11993 9954 11999
rect 9982 12026 10010 12222
rect 9982 11993 10010 11998
rect 10038 12138 10066 12143
rect 10038 11970 10066 12110
rect 10094 12082 10122 12335
rect 10094 12049 10122 12054
rect 10150 12306 10178 12311
rect 10038 11942 10122 11970
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9758 11185 9842 11186
rect 9758 11159 9759 11185
rect 9785 11159 9842 11185
rect 9758 11158 9842 11159
rect 10038 11186 10066 11191
rect 10094 11186 10122 11942
rect 10150 11857 10178 12278
rect 10150 11831 10151 11857
rect 10177 11831 10178 11857
rect 10150 11690 10178 11831
rect 10206 11746 10234 12614
rect 10710 12306 10738 13455
rect 10766 13202 10794 15946
rect 10766 13155 10794 13174
rect 10822 13146 10850 13151
rect 10822 13099 10850 13118
rect 11046 13089 11074 13095
rect 11046 13063 11047 13089
rect 11073 13063 11074 13089
rect 10766 13034 10794 13039
rect 10766 12987 10794 13006
rect 10710 12259 10738 12278
rect 10766 12474 10794 12479
rect 10654 11914 10682 11919
rect 10206 11713 10234 11718
rect 10598 11913 10682 11914
rect 10598 11887 10655 11913
rect 10681 11887 10682 11913
rect 10598 11886 10682 11887
rect 10150 11522 10178 11662
rect 10262 11522 10290 11527
rect 10150 11521 10290 11522
rect 10150 11495 10263 11521
rect 10289 11495 10290 11521
rect 10150 11494 10290 11495
rect 10038 11185 10122 11186
rect 10038 11159 10039 11185
rect 10065 11159 10122 11185
rect 10038 11158 10122 11159
rect 9758 11153 9786 11158
rect 10038 11153 10066 11158
rect 9926 11130 9954 11135
rect 9926 11083 9954 11102
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 9926 10906 9954 10911
rect 10094 10906 10122 11158
rect 10206 11186 10234 11191
rect 10206 11139 10234 11158
rect 10262 10962 10290 11494
rect 10318 11186 10346 11191
rect 10318 11018 10346 11158
rect 10374 11130 10402 11135
rect 10374 11073 10402 11102
rect 10598 11130 10626 11886
rect 10654 11881 10682 11886
rect 10710 11857 10738 11863
rect 10710 11831 10711 11857
rect 10737 11831 10738 11857
rect 10710 11746 10738 11831
rect 10710 11713 10738 11718
rect 10766 11242 10794 12446
rect 10934 12362 10962 12367
rect 11046 12362 11074 13063
rect 11326 12753 11354 12759
rect 11326 12727 11327 12753
rect 11353 12727 11354 12753
rect 11158 12642 11186 12647
rect 11326 12642 11354 12727
rect 11718 12698 11746 12703
rect 11158 12641 11354 12642
rect 11158 12615 11159 12641
rect 11185 12615 11354 12641
rect 11158 12614 11354 12615
rect 11438 12697 11746 12698
rect 11438 12671 11719 12697
rect 11745 12671 11746 12697
rect 11438 12670 11746 12671
rect 11158 12362 11186 12614
rect 10934 12361 11186 12362
rect 10934 12335 10935 12361
rect 10961 12335 11186 12361
rect 10934 12334 11186 12335
rect 10934 12306 10962 12334
rect 10934 12273 10962 12278
rect 11270 12306 11298 12311
rect 11270 12259 11298 12278
rect 11270 12026 11298 12031
rect 11046 11970 11074 11975
rect 10822 11914 10850 11919
rect 10822 11867 10850 11886
rect 10766 11214 10850 11242
rect 10598 11097 10626 11102
rect 10822 11129 10850 11214
rect 11046 11241 11074 11942
rect 11158 11746 11186 11751
rect 11158 11297 11186 11718
rect 11158 11271 11159 11297
rect 11185 11271 11186 11297
rect 11158 11265 11186 11271
rect 11046 11215 11047 11241
rect 11073 11215 11074 11241
rect 11046 11209 11074 11215
rect 10822 11103 10823 11129
rect 10849 11103 10850 11129
rect 10374 11047 10375 11073
rect 10401 11047 10402 11073
rect 10374 11041 10402 11047
rect 10654 11074 10682 11079
rect 10654 11027 10682 11046
rect 10766 11073 10794 11079
rect 10766 11047 10767 11073
rect 10793 11047 10794 11073
rect 10318 10985 10346 10990
rect 10262 10929 10290 10934
rect 10206 10906 10234 10911
rect 9926 10905 10206 10906
rect 9926 10879 9927 10905
rect 9953 10879 10206 10905
rect 9926 10878 10206 10879
rect 9926 10873 9954 10878
rect 9702 10817 9730 10822
rect 9814 10793 9842 10799
rect 9814 10767 9815 10793
rect 9841 10767 9842 10793
rect 9758 10402 9786 10407
rect 9646 10401 9786 10402
rect 9646 10375 9759 10401
rect 9785 10375 9786 10401
rect 9646 10374 9786 10375
rect 9814 10402 9842 10767
rect 9870 10402 9898 10407
rect 9814 10401 9898 10402
rect 9814 10375 9871 10401
rect 9897 10375 9898 10401
rect 9814 10374 9898 10375
rect 9534 9198 9730 9226
rect 9422 9137 9450 9142
rect 9646 9114 9674 9119
rect 9646 8833 9674 9086
rect 9702 8889 9730 9198
rect 9702 8863 9703 8889
rect 9729 8863 9730 8889
rect 9702 8857 9730 8863
rect 9646 8807 9647 8833
rect 9673 8807 9674 8833
rect 9646 8801 9674 8807
rect 9646 8498 9674 8503
rect 9590 8106 9618 8111
rect 9422 8078 9590 8106
rect 9310 8050 9338 8055
rect 9254 8049 9338 8050
rect 9254 8023 9311 8049
rect 9337 8023 9338 8049
rect 9254 8022 9338 8023
rect 9310 8017 9338 8022
rect 9422 8049 9450 8078
rect 9422 8023 9423 8049
rect 9449 8023 9450 8049
rect 9422 8017 9450 8023
rect 9198 7938 9226 7943
rect 9198 7891 9226 7910
rect 9254 7937 9282 7943
rect 9254 7911 9255 7937
rect 9281 7911 9282 7937
rect 9254 7826 9282 7911
rect 9030 7546 9170 7574
rect 9198 7798 9282 7826
rect 8862 7322 8890 7327
rect 8806 7321 8890 7322
rect 8806 7295 8863 7321
rect 8889 7295 8890 7321
rect 8806 7294 8890 7295
rect 8750 7065 8778 7070
rect 8414 6511 8415 6537
rect 8441 6511 8442 6537
rect 8414 6505 8442 6511
rect 8078 6455 8079 6481
rect 8105 6455 8106 6481
rect 8078 6449 8106 6455
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 8750 2618 8778 2623
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8750 400 8778 2590
rect 8862 2561 8890 7294
rect 9030 7265 9058 7546
rect 9030 7239 9031 7265
rect 9057 7239 9058 7265
rect 9030 7233 9058 7239
rect 9198 7265 9226 7798
rect 9478 7770 9506 7775
rect 9478 7713 9506 7742
rect 9478 7687 9479 7713
rect 9505 7687 9506 7713
rect 9478 7574 9506 7687
rect 9590 7657 9618 8078
rect 9590 7631 9591 7657
rect 9617 7631 9618 7657
rect 9590 7625 9618 7631
rect 9478 7546 9562 7574
rect 9198 7239 9199 7265
rect 9225 7239 9226 7265
rect 9198 7233 9226 7239
rect 9366 7266 9394 7271
rect 9366 7265 9450 7266
rect 9366 7239 9367 7265
rect 9393 7239 9450 7265
rect 9366 7238 9450 7239
rect 9366 7233 9394 7238
rect 9198 7154 9226 7159
rect 9198 7107 9226 7126
rect 9422 6985 9450 7238
rect 9534 7210 9562 7546
rect 9590 7210 9618 7215
rect 9534 7209 9618 7210
rect 9534 7183 9591 7209
rect 9617 7183 9618 7209
rect 9534 7182 9618 7183
rect 9590 7177 9618 7182
rect 9422 6959 9423 6985
rect 9449 6959 9450 6985
rect 9422 6953 9450 6959
rect 9590 7098 9618 7103
rect 9534 6929 9562 6935
rect 9534 6903 9535 6929
rect 9561 6903 9562 6929
rect 9478 6537 9506 6543
rect 9478 6511 9479 6537
rect 9505 6511 9506 6537
rect 9478 6370 9506 6511
rect 9534 6370 9562 6903
rect 9590 6929 9618 7070
rect 9590 6903 9591 6929
rect 9617 6903 9618 6929
rect 9590 6897 9618 6903
rect 9646 6986 9674 8470
rect 9758 7994 9786 10374
rect 9814 10290 9842 10295
rect 9870 10290 9898 10374
rect 10094 10402 10122 10407
rect 10206 10402 10234 10878
rect 10766 10906 10794 11047
rect 10822 10906 10850 11103
rect 10878 11130 10906 11135
rect 10878 11083 10906 11102
rect 11214 11074 11242 11079
rect 11158 11073 11242 11074
rect 11158 11047 11215 11073
rect 11241 11047 11242 11073
rect 11158 11046 11242 11047
rect 10822 10878 10906 10906
rect 10766 10873 10794 10878
rect 10318 10850 10346 10855
rect 10318 10737 10346 10822
rect 10318 10711 10319 10737
rect 10345 10711 10346 10737
rect 10318 10705 10346 10711
rect 10374 10849 10402 10855
rect 10374 10823 10375 10849
rect 10401 10823 10402 10849
rect 10318 10458 10346 10463
rect 10318 10411 10346 10430
rect 10262 10402 10290 10407
rect 10206 10401 10290 10402
rect 10206 10375 10263 10401
rect 10289 10375 10290 10401
rect 10206 10374 10290 10375
rect 10094 10355 10122 10374
rect 10262 10369 10290 10374
rect 10374 10402 10402 10823
rect 10374 10369 10402 10374
rect 10542 10793 10570 10799
rect 10542 10767 10543 10793
rect 10569 10767 10570 10793
rect 9870 10262 10122 10290
rect 9814 9786 9842 10262
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9982 10122 10010 10127
rect 10094 10122 10122 10262
rect 9814 9758 9898 9786
rect 9814 9674 9842 9679
rect 9814 9617 9842 9646
rect 9814 9591 9815 9617
rect 9841 9591 9842 9617
rect 9814 9585 9842 9591
rect 9870 9506 9898 9758
rect 9814 9478 9898 9506
rect 9982 9505 10010 10094
rect 9982 9479 9983 9505
rect 10009 9479 10010 9505
rect 9814 9338 9842 9478
rect 9982 9473 10010 9479
rect 10038 10094 10122 10122
rect 10374 10289 10402 10295
rect 10374 10263 10375 10289
rect 10401 10263 10402 10289
rect 10038 9561 10066 10094
rect 10038 9535 10039 9561
rect 10065 9535 10066 9561
rect 10038 9506 10066 9535
rect 10262 9562 10290 9567
rect 10038 9478 10122 9506
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 10094 9338 10122 9478
rect 9814 9310 10010 9338
rect 9982 9281 10010 9310
rect 9982 9255 9983 9281
rect 10009 9255 10010 9281
rect 9982 9249 10010 9255
rect 10038 9310 10122 9338
rect 10038 8834 10066 9310
rect 10038 8801 10066 8806
rect 10150 9225 10178 9231
rect 10150 9199 10151 9225
rect 10177 9199 10178 9225
rect 10150 9170 10178 9199
rect 10206 9226 10234 9231
rect 10206 9179 10234 9198
rect 9814 8777 9842 8783
rect 9814 8751 9815 8777
rect 9841 8751 9842 8777
rect 9814 8106 9842 8751
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9982 8386 10010 8391
rect 9926 8106 9954 8111
rect 9842 8105 9954 8106
rect 9842 8079 9927 8105
rect 9953 8079 9954 8105
rect 9842 8078 9954 8079
rect 9814 8059 9842 8078
rect 9926 8073 9954 8078
rect 9870 7994 9898 7999
rect 9758 7966 9870 7994
rect 9870 7947 9898 7966
rect 9982 7993 10010 8358
rect 10150 8386 10178 9142
rect 10262 9002 10290 9534
rect 10318 9562 10346 9567
rect 10374 9562 10402 10263
rect 10542 10290 10570 10767
rect 10822 10794 10850 10799
rect 10822 10747 10850 10766
rect 10878 10682 10906 10878
rect 11046 10793 11074 10799
rect 11046 10767 11047 10793
rect 11073 10767 11074 10793
rect 10542 10257 10570 10262
rect 10766 10654 10906 10682
rect 10934 10682 10962 10687
rect 10766 10345 10794 10654
rect 10934 10457 10962 10654
rect 11046 10626 11074 10767
rect 11158 10794 11186 11046
rect 11214 11041 11242 11046
rect 11158 10761 11186 10766
rect 11214 10793 11242 10799
rect 11214 10767 11215 10793
rect 11241 10767 11242 10793
rect 11046 10593 11074 10598
rect 10934 10431 10935 10457
rect 10961 10431 10962 10457
rect 10934 10425 10962 10431
rect 10990 10514 11018 10519
rect 10990 10402 11018 10486
rect 11214 10458 11242 10767
rect 11214 10425 11242 10430
rect 11270 10458 11298 11998
rect 11438 12025 11466 12670
rect 11718 12665 11746 12670
rect 12614 12586 12642 18999
rect 12782 18746 12810 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 13062 19138 13090 19143
rect 13062 19091 13090 19110
rect 12782 18713 12810 18718
rect 13398 18746 13426 18751
rect 13398 18699 13426 18718
rect 12894 18633 12922 18639
rect 12894 18607 12895 18633
rect 12921 18607 12922 18633
rect 12894 13454 12922 18607
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 12838 13426 12922 13454
rect 12838 12810 12866 13426
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 12838 12809 12978 12810
rect 12838 12783 12839 12809
rect 12865 12783 12978 12809
rect 12838 12782 12978 12783
rect 12838 12777 12866 12782
rect 12334 12558 12642 12586
rect 11886 12306 11914 12311
rect 11774 12250 11802 12255
rect 11438 11999 11439 12025
rect 11465 11999 11466 12025
rect 11438 11993 11466 11999
rect 11662 12026 11690 12031
rect 11326 11970 11354 11975
rect 11326 11923 11354 11942
rect 11550 11970 11578 11975
rect 11550 11923 11578 11942
rect 11662 11969 11690 11998
rect 11662 11943 11663 11969
rect 11689 11943 11690 11969
rect 11662 11937 11690 11943
rect 11718 11802 11746 11807
rect 11382 11577 11410 11583
rect 11382 11551 11383 11577
rect 11409 11551 11410 11577
rect 11326 11186 11354 11191
rect 11326 11139 11354 11158
rect 11326 10682 11354 10687
rect 11326 10635 11354 10654
rect 11270 10457 11354 10458
rect 11270 10431 11271 10457
rect 11297 10431 11354 10457
rect 11270 10430 11354 10431
rect 11270 10425 11298 10430
rect 11158 10402 11186 10407
rect 10990 10401 11186 10402
rect 10990 10375 10991 10401
rect 11017 10375 11159 10401
rect 11185 10375 11186 10401
rect 10990 10374 11186 10375
rect 10990 10369 11018 10374
rect 10766 10319 10767 10345
rect 10793 10319 10794 10345
rect 10766 10178 10794 10319
rect 10878 10290 10906 10295
rect 10878 10234 10906 10262
rect 10878 10206 11074 10234
rect 10766 10145 10794 10150
rect 10766 10066 10794 10071
rect 10654 9842 10682 9847
rect 10598 9618 10626 9623
rect 10598 9571 10626 9590
rect 10318 9561 10402 9562
rect 10318 9535 10319 9561
rect 10345 9535 10402 9561
rect 10318 9534 10402 9535
rect 10318 9226 10346 9534
rect 10374 9338 10402 9343
rect 10374 9291 10402 9310
rect 10654 9281 10682 9814
rect 10766 9562 10794 10038
rect 10766 9515 10794 9534
rect 10878 9617 10906 9623
rect 10878 9591 10879 9617
rect 10905 9591 10906 9617
rect 10822 9506 10850 9511
rect 10822 9459 10850 9478
rect 10766 9338 10794 9343
rect 10878 9338 10906 9591
rect 10794 9310 10906 9338
rect 10990 9617 11018 9623
rect 10990 9591 10991 9617
rect 11017 9591 11018 9617
rect 10990 9338 11018 9591
rect 11046 9450 11074 10206
rect 11158 9786 11186 10374
rect 11270 10289 11298 10295
rect 11270 10263 11271 10289
rect 11297 10263 11298 10289
rect 11270 10066 11298 10263
rect 11270 10033 11298 10038
rect 11326 9842 11354 10430
rect 11382 9898 11410 11551
rect 11718 11577 11746 11774
rect 11774 11689 11802 12222
rect 11886 12025 11914 12278
rect 12334 12305 12362 12558
rect 12334 12279 12335 12305
rect 12361 12279 12362 12305
rect 12334 12250 12362 12279
rect 12334 12217 12362 12222
rect 12390 12474 12418 12479
rect 11886 11999 11887 12025
rect 11913 11999 11914 12025
rect 11886 11993 11914 11999
rect 12054 12026 12082 12031
rect 11942 11969 11970 11975
rect 11942 11943 11943 11969
rect 11969 11943 11970 11969
rect 11774 11663 11775 11689
rect 11801 11663 11802 11689
rect 11774 11657 11802 11663
rect 11830 11913 11858 11919
rect 11830 11887 11831 11913
rect 11857 11887 11858 11913
rect 11830 11690 11858 11887
rect 11942 11914 11970 11943
rect 12054 11969 12082 11998
rect 12054 11943 12055 11969
rect 12081 11943 12082 11969
rect 12054 11937 12082 11943
rect 11942 11881 11970 11886
rect 12278 11913 12306 11919
rect 12278 11887 12279 11913
rect 12305 11887 12306 11913
rect 12278 11802 12306 11887
rect 12334 11914 12362 11919
rect 12390 11914 12418 12446
rect 12614 12474 12642 12479
rect 12614 12427 12642 12446
rect 12950 12474 12978 12782
rect 20006 12809 20034 12815
rect 20006 12783 20007 12809
rect 20033 12783 20034 12809
rect 18830 12753 18858 12759
rect 18830 12727 18831 12753
rect 18857 12727 18858 12753
rect 12950 12427 12978 12446
rect 13118 12530 13146 12535
rect 13118 12473 13146 12502
rect 18830 12530 18858 12727
rect 18830 12497 18858 12502
rect 13118 12447 13119 12473
rect 13145 12447 13146 12473
rect 13118 12441 13146 12447
rect 20006 12474 20034 12783
rect 20006 12441 20034 12446
rect 12782 12418 12810 12423
rect 12782 12371 12810 12390
rect 18830 12362 18858 12367
rect 18830 12315 18858 12334
rect 20006 12249 20034 12255
rect 20006 12223 20007 12249
rect 20033 12223 20034 12249
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 20006 12138 20034 12223
rect 20006 12105 20034 12110
rect 12446 11970 12474 11975
rect 12446 11923 12474 11942
rect 12334 11913 12418 11914
rect 12334 11887 12335 11913
rect 12361 11887 12418 11913
rect 12334 11886 12418 11887
rect 12334 11881 12362 11886
rect 12278 11769 12306 11774
rect 11886 11690 11914 11695
rect 11830 11689 11914 11690
rect 11830 11663 11887 11689
rect 11913 11663 11914 11689
rect 11830 11662 11914 11663
rect 11886 11657 11914 11662
rect 11718 11551 11719 11577
rect 11745 11551 11746 11577
rect 11718 11298 11746 11551
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 11718 11270 11802 11298
rect 11438 11186 11466 11191
rect 11718 11186 11746 11191
rect 11438 11185 11746 11186
rect 11438 11159 11439 11185
rect 11465 11159 11719 11185
rect 11745 11159 11746 11185
rect 11438 11158 11746 11159
rect 11438 11153 11466 11158
rect 11606 11073 11634 11079
rect 11606 11047 11607 11073
rect 11633 11047 11634 11073
rect 11438 10850 11466 10855
rect 11438 10793 11466 10822
rect 11438 10767 11439 10793
rect 11465 10767 11466 10793
rect 11438 10761 11466 10767
rect 11550 10793 11578 10799
rect 11550 10767 11551 10793
rect 11577 10767 11578 10793
rect 11494 10738 11522 10743
rect 11494 10691 11522 10710
rect 11550 10066 11578 10767
rect 11550 10033 11578 10038
rect 11606 10010 11634 11047
rect 11662 10290 11690 11158
rect 11718 11153 11746 11158
rect 11718 10906 11746 10911
rect 11718 10402 11746 10878
rect 11774 10850 11802 11270
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 18830 11185 18858 11191
rect 18830 11159 18831 11185
rect 18857 11159 18858 11185
rect 18830 10906 18858 11159
rect 18830 10873 18858 10878
rect 11774 10817 11802 10822
rect 13342 10850 13370 10855
rect 13342 10803 13370 10822
rect 13174 10794 13202 10799
rect 12278 10738 12306 10743
rect 12278 10457 12306 10710
rect 12278 10431 12279 10457
rect 12305 10431 12306 10457
rect 12278 10425 12306 10431
rect 12726 10458 12754 10463
rect 11886 10402 11914 10407
rect 11718 10401 11914 10402
rect 11718 10375 11719 10401
rect 11745 10375 11887 10401
rect 11913 10375 11914 10401
rect 11718 10374 11914 10375
rect 11718 10369 11746 10374
rect 11886 10369 11914 10374
rect 11662 10257 11690 10262
rect 12670 10066 12698 10071
rect 12670 10019 12698 10038
rect 12726 10065 12754 10430
rect 13174 10458 13202 10766
rect 18830 10794 18858 10799
rect 18830 10747 18858 10766
rect 20006 10794 20034 11215
rect 20006 10761 20034 10766
rect 20006 10681 20034 10687
rect 20006 10655 20007 10681
rect 20033 10655 20034 10681
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 13174 10425 13202 10430
rect 13342 10458 13370 10463
rect 13342 10411 13370 10430
rect 20006 10458 20034 10655
rect 20006 10425 20034 10430
rect 12726 10039 12727 10065
rect 12753 10039 12754 10065
rect 12726 10033 12754 10039
rect 11606 9977 11634 9982
rect 11718 9953 11746 9959
rect 11718 9927 11719 9953
rect 11745 9927 11746 9953
rect 11718 9898 11746 9927
rect 11382 9870 11746 9898
rect 11326 9814 11690 9842
rect 11158 9758 11354 9786
rect 11102 9618 11130 9623
rect 11102 9571 11130 9590
rect 11046 9422 11186 9450
rect 10990 9310 11074 9338
rect 10766 9305 10794 9310
rect 10654 9255 10655 9281
rect 10681 9255 10682 9281
rect 10654 9249 10682 9255
rect 10710 9282 10738 9287
rect 10710 9235 10738 9254
rect 10318 9179 10346 9198
rect 10766 9226 10794 9231
rect 10262 8969 10290 8974
rect 10150 8353 10178 8358
rect 10206 8834 10234 8839
rect 10206 8274 10234 8806
rect 10766 8778 10794 9198
rect 10822 9226 10850 9231
rect 10934 9226 10962 9231
rect 10822 9225 10962 9226
rect 10822 9199 10823 9225
rect 10849 9199 10935 9225
rect 10961 9199 10962 9225
rect 10822 9198 10962 9199
rect 10822 9193 10850 9198
rect 10934 9193 10962 9198
rect 10990 9225 11018 9231
rect 10990 9199 10991 9225
rect 11017 9199 11018 9225
rect 10990 9170 11018 9199
rect 10990 9137 11018 9142
rect 11046 9114 11074 9310
rect 11102 9170 11130 9175
rect 11102 9123 11130 9142
rect 11158 9114 11186 9422
rect 11214 9226 11242 9231
rect 11214 9179 11242 9198
rect 11326 9225 11354 9758
rect 11606 9674 11634 9679
rect 11606 9627 11634 9646
rect 11662 9617 11690 9814
rect 11662 9591 11663 9617
rect 11689 9591 11690 9617
rect 11662 9585 11690 9591
rect 11494 9561 11522 9567
rect 11494 9535 11495 9561
rect 11521 9535 11522 9561
rect 11438 9506 11466 9511
rect 11494 9506 11522 9535
rect 11466 9478 11522 9506
rect 11438 9473 11466 9478
rect 11718 9450 11746 9870
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 12222 9674 12250 9679
rect 12222 9627 12250 9646
rect 13286 9673 13314 9679
rect 13286 9647 13287 9673
rect 13313 9647 13314 9673
rect 11830 9618 11858 9623
rect 11326 9199 11327 9225
rect 11353 9199 11354 9225
rect 11326 9193 11354 9199
rect 11494 9422 11746 9450
rect 11774 9617 11858 9618
rect 11774 9591 11831 9617
rect 11857 9591 11858 9617
rect 11774 9590 11858 9591
rect 11158 9086 11242 9114
rect 11046 9081 11074 9086
rect 10990 8834 11018 8839
rect 10822 8778 10850 8783
rect 10766 8777 10850 8778
rect 10766 8751 10823 8777
rect 10849 8751 10850 8777
rect 10766 8750 10850 8751
rect 10822 8745 10850 8750
rect 10990 8777 11018 8806
rect 10990 8751 10991 8777
rect 11017 8751 11018 8777
rect 10990 8745 11018 8751
rect 10654 8721 10682 8727
rect 10654 8695 10655 8721
rect 10681 8695 10682 8721
rect 10598 8498 10626 8503
rect 10598 8451 10626 8470
rect 9982 7967 9983 7993
rect 10009 7967 10010 7993
rect 9982 7961 10010 7967
rect 10094 8246 10234 8274
rect 9702 7938 9730 7943
rect 9702 7602 9730 7910
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 10094 7769 10122 8246
rect 10654 8162 10682 8695
rect 11158 8721 11186 8727
rect 11158 8695 11159 8721
rect 11185 8695 11186 8721
rect 10262 8161 10682 8162
rect 10262 8135 10655 8161
rect 10681 8135 10682 8161
rect 10262 8134 10682 8135
rect 10206 7994 10234 7999
rect 10206 7947 10234 7966
rect 10094 7743 10095 7769
rect 10121 7743 10122 7769
rect 10094 7737 10122 7743
rect 10206 7714 10234 7719
rect 10262 7714 10290 8134
rect 10654 8129 10682 8134
rect 10934 8498 10962 8503
rect 10374 7994 10402 7999
rect 10374 7947 10402 7966
rect 10710 7994 10738 7999
rect 10710 7947 10738 7966
rect 10206 7713 10290 7714
rect 10206 7687 10207 7713
rect 10233 7687 10290 7713
rect 10206 7686 10290 7687
rect 10206 7681 10234 7686
rect 10934 7657 10962 8470
rect 11158 8050 11186 8695
rect 11158 8003 11186 8022
rect 11214 7937 11242 9086
rect 11494 8441 11522 9422
rect 11774 8890 11802 9590
rect 11830 9585 11858 9590
rect 13286 9618 13314 9647
rect 20006 9673 20034 9679
rect 20006 9647 20007 9673
rect 20033 9647 20034 9673
rect 13286 9585 13314 9590
rect 18830 9618 18858 9623
rect 18830 9571 18858 9590
rect 20006 9450 20034 9647
rect 20006 9417 20034 9422
rect 12950 9282 12978 9287
rect 11550 8862 11802 8890
rect 11886 9170 11914 9175
rect 11886 8889 11914 9142
rect 11886 8863 11887 8889
rect 11913 8863 11914 8889
rect 11550 8833 11578 8862
rect 11886 8857 11914 8863
rect 12950 8890 12978 9254
rect 18830 9225 18858 9231
rect 18830 9199 18831 9225
rect 18857 9199 18858 9225
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 12950 8843 12978 8862
rect 18830 8890 18858 9199
rect 20006 9114 20034 9119
rect 20006 9067 20034 9086
rect 18830 8857 18858 8862
rect 11550 8807 11551 8833
rect 11577 8807 11578 8833
rect 11550 8498 11578 8807
rect 11550 8465 11578 8470
rect 11494 8415 11495 8441
rect 11521 8415 11522 8441
rect 11494 8409 11522 8415
rect 11438 8386 11466 8391
rect 11438 8161 11466 8358
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 11438 8135 11439 8161
rect 11465 8135 11466 8161
rect 11270 8050 11298 8055
rect 11270 8049 11354 8050
rect 11270 8023 11271 8049
rect 11297 8023 11354 8049
rect 11270 8022 11354 8023
rect 11270 8017 11298 8022
rect 11214 7911 11215 7937
rect 11241 7911 11242 7937
rect 11214 7905 11242 7911
rect 11326 7994 11354 8022
rect 11270 7714 11298 7719
rect 11270 7667 11298 7686
rect 10934 7631 10935 7657
rect 10961 7631 10962 7657
rect 10934 7625 10962 7631
rect 9702 7265 9730 7574
rect 10094 7602 10122 7621
rect 10094 7569 10122 7574
rect 9758 7546 9786 7551
rect 9758 7545 10010 7546
rect 9758 7519 9759 7545
rect 9785 7519 10010 7545
rect 9758 7518 10010 7519
rect 9758 7513 9786 7518
rect 9702 7239 9703 7265
rect 9729 7239 9730 7265
rect 9702 7233 9730 7239
rect 9982 7265 10010 7518
rect 9982 7239 9983 7265
rect 10009 7239 10010 7265
rect 9982 7233 10010 7239
rect 10150 7154 10178 7159
rect 10150 7153 10290 7154
rect 10150 7127 10151 7153
rect 10177 7127 10290 7153
rect 10150 7126 10290 7127
rect 10150 7121 10178 7126
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9646 6958 9898 6986
rect 9646 6706 9674 6958
rect 9870 6873 9898 6958
rect 10262 6929 10290 7126
rect 10262 6903 10263 6929
rect 10289 6903 10290 6929
rect 10262 6897 10290 6903
rect 9870 6847 9871 6873
rect 9897 6847 9898 6873
rect 9870 6841 9898 6847
rect 11326 6817 11354 7966
rect 11438 7714 11466 8135
rect 11438 7681 11466 7686
rect 11494 8050 11522 8055
rect 11494 7993 11522 8022
rect 11494 7967 11495 7993
rect 11521 7967 11522 7993
rect 11494 7602 11522 7967
rect 11494 7569 11522 7574
rect 12334 7602 12362 7621
rect 12334 7569 12362 7574
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 11326 6791 11327 6817
rect 11353 6791 11354 6817
rect 11326 6785 11354 6791
rect 9646 6673 9674 6678
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 9646 6370 9674 6375
rect 9814 6370 9842 6375
rect 9366 6369 9730 6370
rect 9366 6343 9647 6369
rect 9673 6343 9730 6369
rect 9366 6342 9730 6343
rect 9366 6089 9394 6342
rect 9646 6337 9674 6342
rect 9366 6063 9367 6089
rect 9393 6063 9394 6089
rect 9366 6057 9394 6063
rect 9478 6145 9506 6151
rect 9478 6119 9479 6145
rect 9505 6119 9506 6145
rect 9478 4214 9506 6119
rect 9478 4186 9562 4214
rect 9366 2618 9394 2623
rect 9366 2571 9394 2590
rect 8862 2535 8863 2561
rect 8889 2535 8890 2561
rect 8862 2529 8890 2535
rect 9366 2226 9394 2231
rect 9366 2225 9506 2226
rect 9366 2199 9367 2225
rect 9393 2199 9506 2225
rect 9366 2198 9506 2199
rect 9366 2193 9394 2198
rect 9422 2058 9450 2063
rect 9086 1833 9114 1839
rect 9086 1807 9087 1833
rect 9113 1807 9114 1833
rect 9086 400 9114 1807
rect 9422 400 9450 2030
rect 9478 1162 9506 2198
rect 9534 2169 9562 4186
rect 9534 2143 9535 2169
rect 9561 2143 9562 2169
rect 9534 2137 9562 2143
rect 9702 1778 9730 6342
rect 9814 6323 9842 6342
rect 10374 6370 10402 6375
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 10038 2058 10066 2063
rect 10038 2011 10066 2030
rect 9870 1778 9898 1783
rect 9702 1777 9898 1778
rect 9702 1751 9871 1777
rect 9897 1751 9898 1777
rect 9702 1750 9898 1751
rect 9870 1745 9898 1750
rect 10374 1777 10402 6342
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 20118 5361 20146 5367
rect 20118 5335 20119 5361
rect 20145 5335 20146 5361
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 20118 5082 20146 5335
rect 20118 5049 20146 5054
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 20118 2449 20146 2455
rect 20118 2423 20119 2449
rect 20145 2423 20146 2449
rect 20118 2394 20146 2423
rect 20118 2361 20146 2366
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 10374 1751 10375 1777
rect 10401 1751 10402 1777
rect 10374 1745 10402 1751
rect 10094 1722 10122 1727
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 9478 1134 9786 1162
rect 9758 400 9786 1134
rect 10094 400 10122 1694
rect 10878 1722 10906 1727
rect 10878 1665 10906 1694
rect 10878 1639 10879 1665
rect 10905 1639 10906 1665
rect 10878 1633 10906 1639
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 9408 0 9464 400
rect 9744 0 9800 400
rect 10080 0 10136 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 8078 18718 8106 18746
rect 9198 18745 9226 18746
rect 9198 18719 9199 18745
rect 9199 18719 9225 18745
rect 9225 18719 9226 18745
rect 9198 18718 9226 18719
rect 854 18494 882 18522
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 2478 13118 2506 13146
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 966 12446 994 12474
rect 2142 12278 2170 12306
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 966 11241 994 11242
rect 966 11215 967 11241
rect 967 11215 993 11241
rect 993 11215 994 11241
rect 966 11214 994 11215
rect 2142 11185 2170 11186
rect 2142 11159 2143 11185
rect 2143 11159 2169 11185
rect 2169 11159 2170 11185
rect 2142 11158 2170 11159
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 7854 13118 7882 13146
rect 7238 13089 7266 13090
rect 7238 13063 7239 13089
rect 7239 13063 7265 13089
rect 7265 13063 7266 13089
rect 7238 13062 7266 13063
rect 8190 13062 8218 13090
rect 7350 12473 7378 12474
rect 7350 12447 7351 12473
rect 7351 12447 7377 12473
rect 7377 12447 7378 12473
rect 7350 12446 7378 12447
rect 7630 12446 7658 12474
rect 5614 12305 5642 12306
rect 5614 12279 5615 12305
rect 5615 12279 5641 12305
rect 5641 12279 5642 12305
rect 5614 12278 5642 12279
rect 6790 12025 6818 12026
rect 6790 11999 6791 12025
rect 6791 11999 6817 12025
rect 6817 11999 6818 12025
rect 6790 11998 6818 11999
rect 7238 12278 7266 12306
rect 7406 11998 7434 12026
rect 7182 11774 7210 11802
rect 6118 11662 6146 11690
rect 4718 11158 4746 11186
rect 6398 11662 6426 11690
rect 6286 11158 6314 11186
rect 6174 10905 6202 10906
rect 6174 10879 6175 10905
rect 6175 10879 6201 10905
rect 6201 10879 6202 10905
rect 6174 10878 6202 10879
rect 5950 10737 5978 10738
rect 5950 10711 5951 10737
rect 5951 10711 5977 10737
rect 5977 10711 5978 10737
rect 5950 10710 5978 10711
rect 5838 10598 5866 10626
rect 6118 10401 6146 10402
rect 6118 10375 6119 10401
rect 6119 10375 6145 10401
rect 6145 10375 6146 10401
rect 6118 10374 6146 10375
rect 6398 10793 6426 10794
rect 6398 10767 6399 10793
rect 6399 10767 6425 10793
rect 6425 10767 6426 10793
rect 6398 10766 6426 10767
rect 6342 10737 6370 10738
rect 6342 10711 6343 10737
rect 6343 10711 6369 10737
rect 6369 10711 6370 10737
rect 6342 10710 6370 10711
rect 7574 12361 7602 12362
rect 7574 12335 7575 12361
rect 7575 12335 7601 12361
rect 7601 12335 7602 12361
rect 7574 12334 7602 12335
rect 7910 13006 7938 13034
rect 8302 13089 8330 13090
rect 8302 13063 8303 13089
rect 8303 13063 8329 13089
rect 8329 13063 8330 13089
rect 8302 13062 8330 13063
rect 7854 12446 7882 12474
rect 7742 11689 7770 11690
rect 7742 11663 7743 11689
rect 7743 11663 7769 11689
rect 7769 11663 7770 11689
rect 7742 11662 7770 11663
rect 7518 11521 7546 11522
rect 7518 11495 7519 11521
rect 7519 11495 7545 11521
rect 7545 11495 7546 11521
rect 7518 11494 7546 11495
rect 8694 13062 8722 13090
rect 8526 11969 8554 11970
rect 8526 11943 8527 11969
rect 8527 11943 8553 11969
rect 8553 11943 8554 11969
rect 8526 11942 8554 11943
rect 9198 13089 9226 13090
rect 9198 13063 9199 13089
rect 9199 13063 9225 13089
rect 9225 13063 9226 13089
rect 9198 13062 9226 13063
rect 9310 12894 9338 12922
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 10430 19110 10458 19138
rect 11046 19137 11074 19138
rect 11046 19111 11047 19137
rect 11047 19111 11073 19137
rect 11073 19111 11074 19137
rect 11046 19110 11074 19111
rect 12446 19110 12474 19138
rect 10094 18718 10122 18746
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 10710 18745 10738 18746
rect 10710 18719 10711 18745
rect 10711 18719 10737 18745
rect 10737 18719 10738 18745
rect 10710 18718 10738 18719
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 10262 13174 10290 13202
rect 9758 13062 9786 13090
rect 9926 13006 9954 13034
rect 10094 12894 10122 12922
rect 10542 13145 10570 13146
rect 10542 13119 10543 13145
rect 10543 13119 10569 13145
rect 10569 13119 10570 13145
rect 10542 13118 10570 13119
rect 9814 12558 9842 12586
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9646 12390 9674 12418
rect 10094 12390 10122 12418
rect 8918 11942 8946 11970
rect 8190 11774 8218 11802
rect 8638 11774 8666 11802
rect 7798 11270 7826 11298
rect 7910 11494 7938 11522
rect 7910 11214 7938 11242
rect 8414 11241 8442 11242
rect 8414 11215 8415 11241
rect 8415 11215 8441 11241
rect 8441 11215 8442 11241
rect 8414 11214 8442 11215
rect 8638 11185 8666 11186
rect 8638 11159 8639 11185
rect 8639 11159 8665 11185
rect 8665 11159 8666 11185
rect 8638 11158 8666 11159
rect 6678 10905 6706 10906
rect 6678 10879 6679 10905
rect 6679 10879 6705 10905
rect 6705 10879 6706 10905
rect 6678 10878 6706 10879
rect 7406 10849 7434 10850
rect 7406 10823 7407 10849
rect 7407 10823 7433 10849
rect 7433 10823 7434 10849
rect 7406 10822 7434 10823
rect 6790 10766 6818 10794
rect 2478 10262 2506 10290
rect 6678 10401 6706 10402
rect 6678 10375 6679 10401
rect 6679 10375 6705 10401
rect 6705 10375 6706 10401
rect 6678 10374 6706 10375
rect 6846 10486 6874 10514
rect 7294 10486 7322 10514
rect 6790 10345 6818 10346
rect 6790 10319 6791 10345
rect 6791 10319 6817 10345
rect 6817 10319 6818 10345
rect 6790 10318 6818 10319
rect 6230 10038 6258 10066
rect 2142 10009 2170 10010
rect 2142 9983 2143 10009
rect 2143 9983 2169 10009
rect 2169 9983 2170 10009
rect 2142 9982 2170 9983
rect 4774 9982 4802 10010
rect 7462 10318 7490 10346
rect 6678 10038 6706 10066
rect 6454 9982 6482 10010
rect 966 9897 994 9898
rect 966 9871 967 9897
rect 967 9871 993 9897
rect 993 9871 994 9897
rect 966 9870 994 9871
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 7350 9814 7378 9842
rect 6958 9646 6986 9674
rect 6510 9534 6538 9562
rect 6790 9534 6818 9562
rect 2142 9225 2170 9226
rect 2142 9199 2143 9225
rect 2143 9199 2169 9225
rect 2169 9199 2170 9225
rect 2142 9198 2170 9199
rect 4886 9198 4914 9226
rect 6342 9225 6370 9226
rect 6342 9199 6343 9225
rect 6343 9199 6369 9225
rect 6369 9199 6370 9225
rect 6342 9198 6370 9199
rect 966 9113 994 9114
rect 966 9087 967 9113
rect 967 9087 993 9113
rect 993 9087 994 9113
rect 966 9086 994 9087
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 5726 8889 5754 8890
rect 5726 8863 5727 8889
rect 5727 8863 5753 8889
rect 5753 8863 5754 8889
rect 5726 8862 5754 8863
rect 6846 9225 6874 9226
rect 6846 9199 6847 9225
rect 6847 9199 6873 9225
rect 6873 9199 6874 9225
rect 6846 9198 6874 9199
rect 6846 8889 6874 8890
rect 6846 8863 6847 8889
rect 6847 8863 6873 8889
rect 6873 8863 6874 8889
rect 6846 8862 6874 8863
rect 4886 8750 4914 8778
rect 7182 9561 7210 9562
rect 7182 9535 7183 9561
rect 7183 9535 7209 9561
rect 7209 9535 7210 9561
rect 7182 9534 7210 9535
rect 6846 8777 6874 8778
rect 6846 8751 6847 8777
rect 6847 8751 6873 8777
rect 6873 8751 6874 8777
rect 6846 8750 6874 8751
rect 6286 8358 6314 8386
rect 5502 8302 5530 8330
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 2142 8049 2170 8050
rect 2142 8023 2143 8049
rect 2143 8023 2169 8049
rect 2169 8023 2170 8049
rect 2142 8022 2170 8023
rect 966 7742 994 7770
rect 2142 7657 2170 7658
rect 2142 7631 2143 7657
rect 2143 7631 2169 7657
rect 2169 7631 2170 7657
rect 2142 7630 2170 7631
rect 7014 9198 7042 9226
rect 6790 8385 6818 8386
rect 6790 8359 6791 8385
rect 6791 8359 6817 8385
rect 6817 8359 6818 8385
rect 6790 8358 6818 8359
rect 6734 8302 6762 8330
rect 5502 7630 5530 7658
rect 966 7545 994 7546
rect 966 7519 967 7545
rect 967 7519 993 7545
rect 993 7519 994 7545
rect 966 7518 994 7519
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 5614 8022 5642 8050
rect 7126 9142 7154 9170
rect 7070 8974 7098 9002
rect 5614 7854 5642 7882
rect 6398 7910 6426 7938
rect 6958 7937 6986 7938
rect 6958 7911 6959 7937
rect 6959 7911 6985 7937
rect 6985 7911 6986 7937
rect 6958 7910 6986 7911
rect 6902 7854 6930 7882
rect 7014 7742 7042 7770
rect 7630 10905 7658 10906
rect 7630 10879 7631 10905
rect 7631 10879 7657 10905
rect 7657 10879 7658 10905
rect 7630 10878 7658 10879
rect 8134 10878 8162 10906
rect 7798 10793 7826 10794
rect 7798 10767 7799 10793
rect 7799 10767 7825 10793
rect 7825 10767 7826 10793
rect 7798 10766 7826 10767
rect 8302 11073 8330 11074
rect 8302 11047 8303 11073
rect 8303 11047 8329 11073
rect 8329 11047 8330 11073
rect 8302 11046 8330 11047
rect 8638 10934 8666 10962
rect 8246 10849 8274 10850
rect 8246 10823 8247 10849
rect 8247 10823 8273 10849
rect 8273 10823 8274 10849
rect 8246 10822 8274 10823
rect 8414 10766 8442 10794
rect 7910 10345 7938 10346
rect 7910 10319 7911 10345
rect 7911 10319 7937 10345
rect 7937 10319 7938 10345
rect 7910 10318 7938 10319
rect 8078 10345 8106 10346
rect 8078 10319 8079 10345
rect 8079 10319 8105 10345
rect 8105 10319 8106 10345
rect 8078 10318 8106 10319
rect 7686 10038 7714 10066
rect 8246 9646 8274 9674
rect 8918 11662 8946 11690
rect 9422 12334 9450 12362
rect 8862 11438 8890 11466
rect 8806 11297 8834 11298
rect 8806 11271 8807 11297
rect 8807 11271 8833 11297
rect 8833 11271 8834 11297
rect 8806 11270 8834 11271
rect 8918 11270 8946 11298
rect 8694 10486 8722 10514
rect 8694 10374 8722 10402
rect 8974 11185 9002 11186
rect 8974 11159 8975 11185
rect 8975 11159 9001 11185
rect 9001 11159 9002 11185
rect 8974 11158 9002 11159
rect 9870 12361 9898 12362
rect 9870 12335 9871 12361
rect 9871 12335 9897 12361
rect 9897 12335 9898 12361
rect 9870 12334 9898 12335
rect 9870 12222 9898 12250
rect 9702 11998 9730 12026
rect 9534 11438 9562 11466
rect 8918 10934 8946 10962
rect 9030 11129 9058 11130
rect 9030 11103 9031 11129
rect 9031 11103 9057 11129
rect 9057 11103 9058 11129
rect 9030 11102 9058 11103
rect 8974 10766 9002 10794
rect 8806 10430 8834 10458
rect 8694 10065 8722 10066
rect 8694 10039 8695 10065
rect 8695 10039 8721 10065
rect 8721 10039 8722 10065
rect 8694 10038 8722 10039
rect 9142 10878 9170 10906
rect 9198 10822 9226 10850
rect 9086 10374 9114 10402
rect 8862 10345 8890 10346
rect 8862 10319 8863 10345
rect 8863 10319 8889 10345
rect 8889 10319 8890 10345
rect 8862 10318 8890 10319
rect 9142 10766 9170 10794
rect 9254 10430 9282 10458
rect 9198 10374 9226 10402
rect 9254 10289 9282 10290
rect 9254 10263 9255 10289
rect 9255 10263 9281 10289
rect 9281 10263 9282 10289
rect 9254 10262 9282 10263
rect 8694 9814 8722 9842
rect 8862 9702 8890 9730
rect 8358 9590 8386 9618
rect 7910 9198 7938 9226
rect 8470 9617 8498 9618
rect 8470 9591 8471 9617
rect 8471 9591 8497 9617
rect 8497 9591 8498 9617
rect 8470 9590 8498 9591
rect 8806 9617 8834 9618
rect 8806 9591 8807 9617
rect 8807 9591 8833 9617
rect 8833 9591 8834 9617
rect 8806 9590 8834 9591
rect 8806 9478 8834 9506
rect 8806 9198 8834 9226
rect 9030 9590 9058 9618
rect 8918 9198 8946 9226
rect 7518 8974 7546 9002
rect 8750 9086 8778 9114
rect 8414 7657 8442 7658
rect 8414 7631 8415 7657
rect 8415 7631 8441 7657
rect 8441 7631 8442 7657
rect 8414 7630 8442 7631
rect 8302 7574 8330 7602
rect 8414 7126 8442 7154
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 7462 6678 7490 6706
rect 8078 6678 8106 6706
rect 2342 6650 2370 6651
rect 8918 7769 8946 7770
rect 8918 7743 8919 7769
rect 8919 7743 8945 7769
rect 8945 7743 8946 7769
rect 8918 7742 8946 7743
rect 9142 9702 9170 9730
rect 8862 7657 8890 7658
rect 8862 7631 8863 7657
rect 8863 7631 8889 7657
rect 8889 7631 8890 7657
rect 8862 7630 8890 7631
rect 9030 7574 9058 7602
rect 9254 9646 9282 9674
rect 9198 9086 9226 9114
rect 9310 9617 9338 9618
rect 9310 9591 9311 9617
rect 9311 9591 9337 9617
rect 9337 9591 9338 9617
rect 9310 9590 9338 9591
rect 9646 11185 9674 11186
rect 9646 11159 9647 11185
rect 9647 11159 9673 11185
rect 9673 11159 9674 11185
rect 9646 11158 9674 11159
rect 9590 10598 9618 10626
rect 9590 10513 9618 10514
rect 9590 10487 9591 10513
rect 9591 10487 9617 10513
rect 9617 10487 9618 10513
rect 9590 10486 9618 10487
rect 9982 12361 10010 12362
rect 9982 12335 9983 12361
rect 9983 12335 10009 12361
rect 10009 12335 10010 12361
rect 9982 12334 10010 12335
rect 9926 12166 9954 12194
rect 9926 12054 9954 12082
rect 9982 11998 10010 12026
rect 10038 12110 10066 12138
rect 10094 12054 10122 12082
rect 10150 12278 10178 12306
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 10766 13201 10794 13202
rect 10766 13175 10767 13201
rect 10767 13175 10793 13201
rect 10793 13175 10794 13201
rect 10766 13174 10794 13175
rect 10822 13145 10850 13146
rect 10822 13119 10823 13145
rect 10823 13119 10849 13145
rect 10849 13119 10850 13145
rect 10822 13118 10850 13119
rect 10766 13033 10794 13034
rect 10766 13007 10767 13033
rect 10767 13007 10793 13033
rect 10793 13007 10794 13033
rect 10766 13006 10794 13007
rect 10710 12305 10738 12306
rect 10710 12279 10711 12305
rect 10711 12279 10737 12305
rect 10737 12279 10738 12305
rect 10710 12278 10738 12279
rect 10766 12446 10794 12474
rect 10206 11718 10234 11746
rect 10150 11662 10178 11690
rect 9926 11129 9954 11130
rect 9926 11103 9927 11129
rect 9927 11103 9953 11129
rect 9953 11103 9954 11129
rect 9926 11102 9954 11103
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 10206 11185 10234 11186
rect 10206 11159 10207 11185
rect 10207 11159 10233 11185
rect 10233 11159 10234 11185
rect 10206 11158 10234 11159
rect 10318 11185 10346 11186
rect 10318 11159 10319 11185
rect 10319 11159 10345 11185
rect 10345 11159 10346 11185
rect 10318 11158 10346 11159
rect 10374 11102 10402 11130
rect 10710 11718 10738 11746
rect 10934 12278 10962 12306
rect 11270 12305 11298 12306
rect 11270 12279 11271 12305
rect 11271 12279 11297 12305
rect 11297 12279 11298 12305
rect 11270 12278 11298 12279
rect 11270 11998 11298 12026
rect 11046 11942 11074 11970
rect 10822 11913 10850 11914
rect 10822 11887 10823 11913
rect 10823 11887 10849 11913
rect 10849 11887 10850 11913
rect 10822 11886 10850 11887
rect 10598 11102 10626 11130
rect 11158 11718 11186 11746
rect 10654 11073 10682 11074
rect 10654 11047 10655 11073
rect 10655 11047 10681 11073
rect 10681 11047 10682 11073
rect 10654 11046 10682 11047
rect 10318 10990 10346 11018
rect 10262 10934 10290 10962
rect 10206 10878 10234 10906
rect 9702 10822 9730 10850
rect 9422 9142 9450 9170
rect 9646 9086 9674 9114
rect 9646 8470 9674 8498
rect 9590 8078 9618 8106
rect 9198 7937 9226 7938
rect 9198 7911 9199 7937
rect 9199 7911 9225 7937
rect 9225 7911 9226 7937
rect 9198 7910 9226 7911
rect 8750 7070 8778 7098
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 8750 2590 8778 2618
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9478 7742 9506 7770
rect 9198 7153 9226 7154
rect 9198 7127 9199 7153
rect 9199 7127 9225 7153
rect 9225 7127 9226 7153
rect 9198 7126 9226 7127
rect 9590 7070 9618 7098
rect 9814 10262 9842 10290
rect 10094 10401 10122 10402
rect 10094 10375 10095 10401
rect 10095 10375 10121 10401
rect 10121 10375 10122 10401
rect 10094 10374 10122 10375
rect 10766 10878 10794 10906
rect 10878 11129 10906 11130
rect 10878 11103 10879 11129
rect 10879 11103 10905 11129
rect 10905 11103 10906 11129
rect 10878 11102 10906 11103
rect 10318 10822 10346 10850
rect 10318 10457 10346 10458
rect 10318 10431 10319 10457
rect 10319 10431 10345 10457
rect 10345 10431 10346 10457
rect 10318 10430 10346 10431
rect 10374 10374 10402 10402
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9982 10094 10010 10122
rect 9814 9646 9842 9674
rect 10262 9534 10290 9562
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 10038 8806 10066 8834
rect 10206 9225 10234 9226
rect 10206 9199 10207 9225
rect 10207 9199 10233 9225
rect 10233 9199 10234 9225
rect 10206 9198 10234 9199
rect 10150 9142 10178 9170
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 9982 8358 10010 8386
rect 9814 8078 9842 8106
rect 9870 7993 9898 7994
rect 9870 7967 9871 7993
rect 9871 7967 9897 7993
rect 9897 7967 9898 7993
rect 9870 7966 9898 7967
rect 10822 10793 10850 10794
rect 10822 10767 10823 10793
rect 10823 10767 10849 10793
rect 10849 10767 10850 10793
rect 10822 10766 10850 10767
rect 10542 10262 10570 10290
rect 10934 10654 10962 10682
rect 11158 10766 11186 10794
rect 11046 10598 11074 10626
rect 10990 10486 11018 10514
rect 11214 10430 11242 10458
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 13062 19137 13090 19138
rect 13062 19111 13063 19137
rect 13063 19111 13089 19137
rect 13089 19111 13090 19137
rect 13062 19110 13090 19111
rect 12782 18718 12810 18746
rect 13398 18745 13426 18746
rect 13398 18719 13399 18745
rect 13399 18719 13425 18745
rect 13425 18719 13426 18745
rect 13398 18718 13426 18719
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 11886 12278 11914 12306
rect 11774 12222 11802 12250
rect 11662 11998 11690 12026
rect 11326 11969 11354 11970
rect 11326 11943 11327 11969
rect 11327 11943 11353 11969
rect 11353 11943 11354 11969
rect 11326 11942 11354 11943
rect 11550 11969 11578 11970
rect 11550 11943 11551 11969
rect 11551 11943 11577 11969
rect 11577 11943 11578 11969
rect 11550 11942 11578 11943
rect 11718 11774 11746 11802
rect 11326 11185 11354 11186
rect 11326 11159 11327 11185
rect 11327 11159 11353 11185
rect 11353 11159 11354 11185
rect 11326 11158 11354 11159
rect 11326 10681 11354 10682
rect 11326 10655 11327 10681
rect 11327 10655 11353 10681
rect 11353 10655 11354 10681
rect 11326 10654 11354 10655
rect 10878 10289 10906 10290
rect 10878 10263 10879 10289
rect 10879 10263 10905 10289
rect 10905 10263 10906 10289
rect 10878 10262 10906 10263
rect 10766 10150 10794 10178
rect 10766 10038 10794 10066
rect 10654 9814 10682 9842
rect 10598 9617 10626 9618
rect 10598 9591 10599 9617
rect 10599 9591 10625 9617
rect 10625 9591 10626 9617
rect 10598 9590 10626 9591
rect 10374 9337 10402 9338
rect 10374 9311 10375 9337
rect 10375 9311 10401 9337
rect 10401 9311 10402 9337
rect 10374 9310 10402 9311
rect 10766 9561 10794 9562
rect 10766 9535 10767 9561
rect 10767 9535 10793 9561
rect 10793 9535 10794 9561
rect 10766 9534 10794 9535
rect 10822 9505 10850 9506
rect 10822 9479 10823 9505
rect 10823 9479 10849 9505
rect 10849 9479 10850 9505
rect 10822 9478 10850 9479
rect 10766 9310 10794 9338
rect 11270 10038 11298 10066
rect 12334 12222 12362 12250
rect 12390 12446 12418 12474
rect 12054 11998 12082 12026
rect 11942 11886 11970 11914
rect 12614 12473 12642 12474
rect 12614 12447 12615 12473
rect 12615 12447 12641 12473
rect 12641 12447 12642 12473
rect 12614 12446 12642 12447
rect 12950 12473 12978 12474
rect 12950 12447 12951 12473
rect 12951 12447 12977 12473
rect 12977 12447 12978 12473
rect 12950 12446 12978 12447
rect 13118 12502 13146 12530
rect 18830 12502 18858 12530
rect 20006 12446 20034 12474
rect 12782 12417 12810 12418
rect 12782 12391 12783 12417
rect 12783 12391 12809 12417
rect 12809 12391 12810 12417
rect 12782 12390 12810 12391
rect 18830 12361 18858 12362
rect 18830 12335 18831 12361
rect 18831 12335 18857 12361
rect 18857 12335 18858 12361
rect 18830 12334 18858 12335
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 20006 12110 20034 12138
rect 12446 11969 12474 11970
rect 12446 11943 12447 11969
rect 12447 11943 12473 11969
rect 12473 11943 12474 11969
rect 12446 11942 12474 11943
rect 12278 11774 12306 11802
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 11438 10822 11466 10850
rect 11494 10737 11522 10738
rect 11494 10711 11495 10737
rect 11495 10711 11521 10737
rect 11521 10711 11522 10737
rect 11494 10710 11522 10711
rect 11550 10038 11578 10066
rect 11718 10878 11746 10906
rect 18830 10878 18858 10906
rect 11774 10822 11802 10850
rect 13342 10849 13370 10850
rect 13342 10823 13343 10849
rect 13343 10823 13369 10849
rect 13369 10823 13370 10849
rect 13342 10822 13370 10823
rect 13174 10793 13202 10794
rect 13174 10767 13175 10793
rect 13175 10767 13201 10793
rect 13201 10767 13202 10793
rect 13174 10766 13202 10767
rect 12278 10710 12306 10738
rect 12726 10430 12754 10458
rect 11662 10262 11690 10290
rect 12670 10065 12698 10066
rect 12670 10039 12671 10065
rect 12671 10039 12697 10065
rect 12697 10039 12698 10065
rect 12670 10038 12698 10039
rect 18830 10793 18858 10794
rect 18830 10767 18831 10793
rect 18831 10767 18857 10793
rect 18857 10767 18858 10793
rect 18830 10766 18858 10767
rect 20006 10766 20034 10794
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 13174 10430 13202 10458
rect 13342 10457 13370 10458
rect 13342 10431 13343 10457
rect 13343 10431 13369 10457
rect 13369 10431 13370 10457
rect 13342 10430 13370 10431
rect 20006 10430 20034 10458
rect 11606 9982 11634 10010
rect 11102 9617 11130 9618
rect 11102 9591 11103 9617
rect 11103 9591 11129 9617
rect 11129 9591 11130 9617
rect 11102 9590 11130 9591
rect 10710 9281 10738 9282
rect 10710 9255 10711 9281
rect 10711 9255 10737 9281
rect 10737 9255 10738 9281
rect 10710 9254 10738 9255
rect 10318 9225 10346 9226
rect 10318 9199 10319 9225
rect 10319 9199 10345 9225
rect 10345 9199 10346 9225
rect 10318 9198 10346 9199
rect 10766 9198 10794 9226
rect 10262 8974 10290 9002
rect 10150 8358 10178 8386
rect 10206 8806 10234 8834
rect 10990 9142 11018 9170
rect 11102 9169 11130 9170
rect 11102 9143 11103 9169
rect 11103 9143 11129 9169
rect 11129 9143 11130 9169
rect 11102 9142 11130 9143
rect 11046 9086 11074 9114
rect 11214 9225 11242 9226
rect 11214 9199 11215 9225
rect 11215 9199 11241 9225
rect 11241 9199 11242 9225
rect 11214 9198 11242 9199
rect 11606 9673 11634 9674
rect 11606 9647 11607 9673
rect 11607 9647 11633 9673
rect 11633 9647 11634 9673
rect 11606 9646 11634 9647
rect 11438 9478 11466 9506
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 12222 9673 12250 9674
rect 12222 9647 12223 9673
rect 12223 9647 12249 9673
rect 12249 9647 12250 9673
rect 12222 9646 12250 9647
rect 10990 8806 11018 8834
rect 10598 8497 10626 8498
rect 10598 8471 10599 8497
rect 10599 8471 10625 8497
rect 10625 8471 10626 8497
rect 10598 8470 10626 8471
rect 9702 7910 9730 7938
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 10206 7993 10234 7994
rect 10206 7967 10207 7993
rect 10207 7967 10233 7993
rect 10233 7967 10234 7993
rect 10206 7966 10234 7967
rect 10934 8470 10962 8498
rect 10374 7993 10402 7994
rect 10374 7967 10375 7993
rect 10375 7967 10401 7993
rect 10401 7967 10402 7993
rect 10374 7966 10402 7967
rect 10710 7993 10738 7994
rect 10710 7967 10711 7993
rect 10711 7967 10737 7993
rect 10737 7967 10738 7993
rect 10710 7966 10738 7967
rect 11158 8049 11186 8050
rect 11158 8023 11159 8049
rect 11159 8023 11185 8049
rect 11185 8023 11186 8049
rect 11158 8022 11186 8023
rect 13286 9590 13314 9618
rect 18830 9617 18858 9618
rect 18830 9591 18831 9617
rect 18831 9591 18857 9617
rect 18857 9591 18858 9617
rect 18830 9590 18858 9591
rect 20006 9422 20034 9450
rect 12950 9254 12978 9282
rect 11886 9142 11914 9170
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 12950 8889 12978 8890
rect 12950 8863 12951 8889
rect 12951 8863 12977 8889
rect 12977 8863 12978 8889
rect 12950 8862 12978 8863
rect 20006 9113 20034 9114
rect 20006 9087 20007 9113
rect 20007 9087 20033 9113
rect 20033 9087 20034 9113
rect 20006 9086 20034 9087
rect 18830 8862 18858 8890
rect 11550 8470 11578 8498
rect 11438 8358 11466 8386
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 11326 7966 11354 7994
rect 11270 7713 11298 7714
rect 11270 7687 11271 7713
rect 11271 7687 11297 7713
rect 11297 7687 11298 7713
rect 11270 7686 11298 7687
rect 9702 7574 9730 7602
rect 10094 7601 10122 7602
rect 10094 7575 10095 7601
rect 10095 7575 10121 7601
rect 10121 7575 10122 7601
rect 10094 7574 10122 7575
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 11438 7686 11466 7714
rect 11494 8022 11522 8050
rect 11494 7574 11522 7602
rect 12334 7601 12362 7602
rect 12334 7575 12335 7601
rect 12335 7575 12361 7601
rect 12361 7575 12362 7601
rect 12334 7574 12362 7575
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 9646 6678 9674 6706
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 9366 2617 9394 2618
rect 9366 2591 9367 2617
rect 9367 2591 9393 2617
rect 9393 2591 9394 2617
rect 9366 2590 9394 2591
rect 9422 2030 9450 2058
rect 9814 6369 9842 6370
rect 9814 6343 9815 6369
rect 9815 6343 9841 6369
rect 9841 6343 9842 6369
rect 9814 6342 9842 6343
rect 10374 6342 10402 6370
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 10038 2057 10066 2058
rect 10038 2031 10039 2057
rect 10039 2031 10065 2057
rect 10065 2031 10066 2057
rect 10038 2030 10066 2031
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 20118 5054 20146 5082
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 20118 2366 20146 2394
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 10094 1694 10122 1722
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 10878 1694 10906 1722
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 10425 19110 10430 19138
rect 10458 19110 11046 19138
rect 11074 19110 11079 19138
rect 12441 19110 12446 19138
rect 12474 19110 13062 19138
rect 13090 19110 13095 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 8073 18718 8078 18746
rect 8106 18718 9198 18746
rect 9226 18718 9231 18746
rect 10089 18718 10094 18746
rect 10122 18718 10710 18746
rect 10738 18718 10743 18746
rect 12777 18718 12782 18746
rect 12810 18718 13398 18746
rect 13426 18718 13431 18746
rect 0 18522 400 18536
rect 0 18494 854 18522
rect 882 18494 887 18522
rect 0 18480 400 18494
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 10257 13174 10262 13202
rect 10290 13174 10766 13202
rect 10794 13174 10799 13202
rect 0 13146 400 13160
rect 0 13118 2478 13146
rect 2506 13118 2511 13146
rect 7849 13118 7854 13146
rect 7882 13118 10542 13146
rect 10570 13118 10822 13146
rect 10850 13118 10855 13146
rect 0 13104 400 13118
rect 7233 13062 7238 13090
rect 7266 13062 8190 13090
rect 8218 13062 8223 13090
rect 8297 13062 8302 13090
rect 8330 13062 8694 13090
rect 8722 13062 8727 13090
rect 9193 13062 9198 13090
rect 9226 13062 9758 13090
rect 9786 13062 9791 13090
rect 8302 13034 8330 13062
rect 7905 13006 7910 13034
rect 7938 13006 8330 13034
rect 9921 13006 9926 13034
rect 9954 13006 10766 13034
rect 10794 13006 10799 13034
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 9305 12894 9310 12922
rect 9338 12894 10094 12922
rect 10122 12894 10127 12922
rect 9809 12558 9814 12586
rect 9842 12558 9847 12586
rect 0 12474 400 12488
rect 9814 12474 9842 12558
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 13113 12502 13118 12530
rect 13146 12502 18830 12530
rect 18858 12502 18863 12530
rect 20600 12474 21000 12488
rect 0 12446 966 12474
rect 994 12446 999 12474
rect 7345 12446 7350 12474
rect 7378 12446 7630 12474
rect 7658 12446 7854 12474
rect 7882 12446 7887 12474
rect 9814 12446 10766 12474
rect 10794 12446 10799 12474
rect 12385 12446 12390 12474
rect 12418 12446 12614 12474
rect 12642 12446 12950 12474
rect 12978 12446 12983 12474
rect 20001 12446 20006 12474
rect 20034 12446 21000 12474
rect 0 12432 400 12446
rect 20600 12432 21000 12446
rect 9641 12390 9646 12418
rect 9674 12390 10094 12418
rect 10122 12390 10127 12418
rect 12777 12390 12782 12418
rect 12810 12390 15974 12418
rect 15946 12362 15974 12390
rect 7569 12334 7574 12362
rect 7602 12334 9422 12362
rect 9450 12334 9870 12362
rect 9898 12334 9903 12362
rect 9977 12334 9982 12362
rect 10010 12334 10015 12362
rect 15946 12334 18830 12362
rect 18858 12334 18863 12362
rect 2137 12278 2142 12306
rect 2170 12278 5614 12306
rect 5642 12278 7238 12306
rect 7266 12278 7271 12306
rect 9982 12250 10010 12334
rect 10145 12278 10150 12306
rect 10178 12278 10710 12306
rect 10738 12278 10934 12306
rect 10962 12278 10967 12306
rect 11265 12278 11270 12306
rect 11298 12278 11886 12306
rect 11914 12278 11919 12306
rect 9865 12222 9870 12250
rect 9898 12222 10010 12250
rect 11769 12222 11774 12250
rect 11802 12222 12334 12250
rect 12362 12222 12367 12250
rect 9921 12166 9926 12194
rect 9954 12166 9959 12194
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 9926 12138 9954 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 20600 12138 21000 12152
rect 9926 12110 10038 12138
rect 10066 12110 10071 12138
rect 20001 12110 20006 12138
rect 20034 12110 21000 12138
rect 20600 12096 21000 12110
rect 9921 12054 9926 12082
rect 9954 12054 10094 12082
rect 10122 12054 10127 12082
rect 6785 11998 6790 12026
rect 6818 11998 7406 12026
rect 7434 11998 7439 12026
rect 9697 11998 9702 12026
rect 9730 11998 9982 12026
rect 10010 11998 10015 12026
rect 11265 11998 11270 12026
rect 11298 11998 11662 12026
rect 11690 11998 12054 12026
rect 12082 11998 12087 12026
rect 8521 11942 8526 11970
rect 8554 11942 8918 11970
rect 8946 11942 8951 11970
rect 11041 11942 11046 11970
rect 11074 11942 11326 11970
rect 11354 11942 11359 11970
rect 11545 11942 11550 11970
rect 11578 11942 12446 11970
rect 12474 11942 12479 11970
rect 10817 11886 10822 11914
rect 10850 11886 11942 11914
rect 11970 11886 11975 11914
rect 7177 11774 7182 11802
rect 7210 11774 7215 11802
rect 8185 11774 8190 11802
rect 8218 11774 8638 11802
rect 8666 11774 8671 11802
rect 11713 11774 11718 11802
rect 11746 11774 12278 11802
rect 12306 11774 12311 11802
rect 7182 11690 7210 11774
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 10201 11718 10206 11746
rect 10234 11718 10710 11746
rect 10738 11718 11158 11746
rect 11186 11718 11191 11746
rect 6113 11662 6118 11690
rect 6146 11662 6398 11690
rect 6426 11662 7742 11690
rect 7770 11662 8918 11690
rect 8946 11662 10150 11690
rect 10178 11662 10183 11690
rect 7513 11494 7518 11522
rect 7546 11494 7910 11522
rect 7938 11494 7943 11522
rect 8857 11438 8862 11466
rect 8890 11438 9534 11466
rect 9562 11438 9567 11466
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 7793 11270 7798 11298
rect 7826 11270 8806 11298
rect 8834 11270 8918 11298
rect 8946 11270 8951 11298
rect 961 11214 966 11242
rect 994 11214 999 11242
rect 7905 11214 7910 11242
rect 7938 11214 8414 11242
rect 8442 11214 8447 11242
rect 0 11130 400 11144
rect 966 11130 994 11214
rect 2137 11158 2142 11186
rect 2170 11158 4718 11186
rect 4746 11158 6286 11186
rect 6314 11158 6319 11186
rect 8633 11158 8638 11186
rect 8666 11158 8974 11186
rect 9002 11158 9007 11186
rect 9641 11158 9646 11186
rect 9674 11158 10206 11186
rect 10234 11158 10239 11186
rect 10313 11158 10318 11186
rect 10346 11158 11326 11186
rect 11354 11158 11359 11186
rect 0 11102 994 11130
rect 9025 11102 9030 11130
rect 9058 11102 9926 11130
rect 9954 11102 9959 11130
rect 10369 11102 10374 11130
rect 10402 11102 10598 11130
rect 10626 11102 10878 11130
rect 10906 11102 10911 11130
rect 0 11088 400 11102
rect 8297 11046 8302 11074
rect 8330 11046 10654 11074
rect 10682 11046 10687 11074
rect 10094 10990 10318 11018
rect 10346 10990 10351 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 8633 10934 8638 10962
rect 8666 10934 8918 10962
rect 8946 10934 8951 10962
rect 10094 10906 10122 10990
rect 10257 10934 10262 10962
rect 10290 10934 10906 10962
rect 10878 10906 10906 10934
rect 6169 10878 6174 10906
rect 6202 10878 6678 10906
rect 6706 10878 7630 10906
rect 7658 10878 8134 10906
rect 8162 10878 8167 10906
rect 9137 10878 9142 10906
rect 9170 10878 10122 10906
rect 10201 10878 10206 10906
rect 10234 10878 10766 10906
rect 10794 10878 10799 10906
rect 10878 10878 11718 10906
rect 11746 10878 11751 10906
rect 15946 10878 18830 10906
rect 18858 10878 18863 10906
rect 15946 10850 15974 10878
rect 7401 10822 7406 10850
rect 7434 10822 8246 10850
rect 8274 10822 9198 10850
rect 9226 10822 9231 10850
rect 9697 10822 9702 10850
rect 9730 10822 10318 10850
rect 10346 10822 11438 10850
rect 11466 10822 11774 10850
rect 11802 10822 11807 10850
rect 13337 10822 13342 10850
rect 13370 10822 15974 10850
rect 20600 10794 21000 10808
rect 6393 10766 6398 10794
rect 6426 10766 6790 10794
rect 6818 10766 6823 10794
rect 7793 10766 7798 10794
rect 7826 10766 8414 10794
rect 8442 10766 8447 10794
rect 8969 10766 8974 10794
rect 9002 10766 9142 10794
rect 9170 10766 10822 10794
rect 10850 10766 11158 10794
rect 11186 10766 11191 10794
rect 13169 10766 13174 10794
rect 13202 10766 18830 10794
rect 18858 10766 18863 10794
rect 20001 10766 20006 10794
rect 20034 10766 21000 10794
rect 20600 10752 21000 10766
rect 5945 10710 5950 10738
rect 5978 10710 6342 10738
rect 6370 10710 6375 10738
rect 11489 10710 11494 10738
rect 11522 10710 12278 10738
rect 12306 10710 12311 10738
rect 10929 10654 10934 10682
rect 10962 10654 11326 10682
rect 11354 10654 11359 10682
rect 5833 10598 5838 10626
rect 5866 10598 9590 10626
rect 9618 10598 11046 10626
rect 11074 10598 11079 10626
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 6841 10486 6846 10514
rect 6874 10486 7294 10514
rect 7322 10486 8694 10514
rect 8722 10486 9590 10514
rect 9618 10486 9623 10514
rect 10206 10486 10990 10514
rect 11018 10486 11023 10514
rect 10206 10458 10234 10486
rect 20600 10458 21000 10472
rect 8801 10430 8806 10458
rect 8834 10430 9254 10458
rect 9282 10430 10234 10458
rect 10313 10430 10318 10458
rect 10346 10430 11214 10458
rect 11242 10430 11247 10458
rect 12721 10430 12726 10458
rect 12754 10430 13174 10458
rect 13202 10430 13342 10458
rect 13370 10430 13375 10458
rect 20001 10430 20006 10458
rect 20034 10430 21000 10458
rect 20600 10416 21000 10430
rect 6113 10374 6118 10402
rect 6146 10374 6678 10402
rect 6706 10374 6711 10402
rect 8689 10374 8694 10402
rect 8722 10374 9086 10402
rect 9114 10374 9119 10402
rect 9193 10374 9198 10402
rect 9226 10374 10094 10402
rect 10122 10374 10374 10402
rect 10402 10374 10407 10402
rect 9086 10346 9114 10374
rect 6785 10318 6790 10346
rect 6818 10318 7462 10346
rect 7490 10318 7910 10346
rect 7938 10318 7943 10346
rect 8073 10318 8078 10346
rect 8106 10318 8862 10346
rect 8890 10318 8895 10346
rect 9086 10318 9842 10346
rect 9814 10290 9842 10318
rect 2473 10262 2478 10290
rect 2506 10262 9254 10290
rect 9282 10262 9287 10290
rect 9809 10262 9814 10290
rect 9842 10262 9847 10290
rect 10537 10262 10542 10290
rect 10570 10262 10878 10290
rect 10906 10262 11662 10290
rect 11690 10262 11695 10290
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 10094 10150 10766 10178
rect 10794 10150 10799 10178
rect 10094 10122 10122 10150
rect 9977 10094 9982 10122
rect 10010 10094 10122 10122
rect 6225 10038 6230 10066
rect 6258 10038 6678 10066
rect 6706 10038 6711 10066
rect 7681 10038 7686 10066
rect 7714 10038 8694 10066
rect 8722 10038 8727 10066
rect 10761 10038 10766 10066
rect 10794 10038 11270 10066
rect 11298 10038 11303 10066
rect 11545 10038 11550 10066
rect 11578 10038 12670 10066
rect 12698 10038 12703 10066
rect 11270 10010 11298 10038
rect 2137 9982 2142 10010
rect 2170 9982 4774 10010
rect 4802 9982 6454 10010
rect 6482 9982 6487 10010
rect 11270 9982 11606 10010
rect 11634 9982 11639 10010
rect 961 9870 966 9898
rect 994 9870 999 9898
rect 0 9786 400 9800
rect 966 9786 994 9870
rect 7345 9814 7350 9842
rect 7378 9814 8694 9842
rect 8722 9814 10654 9842
rect 10682 9814 10687 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 0 9758 994 9786
rect 0 9744 400 9758
rect 8857 9702 8862 9730
rect 8890 9702 9142 9730
rect 9170 9702 9175 9730
rect 6953 9646 6958 9674
rect 6986 9646 8246 9674
rect 8274 9646 9254 9674
rect 9282 9646 9814 9674
rect 9842 9646 9847 9674
rect 11601 9646 11606 9674
rect 11634 9646 12222 9674
rect 12250 9646 12255 9674
rect 13426 9646 15974 9674
rect 13426 9618 13454 9646
rect 8353 9590 8358 9618
rect 8386 9590 8470 9618
rect 8498 9590 8806 9618
rect 8834 9590 9030 9618
rect 9058 9590 9063 9618
rect 9305 9590 9310 9618
rect 9338 9590 10598 9618
rect 10626 9590 10631 9618
rect 11097 9590 11102 9618
rect 11130 9590 13286 9618
rect 13314 9590 13454 9618
rect 15946 9618 15974 9646
rect 15946 9590 18830 9618
rect 18858 9590 18863 9618
rect 6505 9534 6510 9562
rect 6538 9534 6790 9562
rect 6818 9534 7182 9562
rect 7210 9534 7215 9562
rect 9310 9506 9338 9590
rect 10257 9534 10262 9562
rect 10290 9534 10766 9562
rect 10794 9534 10799 9562
rect 8801 9478 8806 9506
rect 8834 9478 9338 9506
rect 10817 9478 10822 9506
rect 10850 9478 11438 9506
rect 11466 9478 11471 9506
rect 20600 9450 21000 9464
rect 20001 9422 20006 9450
rect 20034 9422 21000 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 20600 9408 21000 9422
rect 10369 9310 10374 9338
rect 10402 9310 10766 9338
rect 10794 9310 10799 9338
rect 10705 9254 10710 9282
rect 10738 9254 12950 9282
rect 12978 9254 12983 9282
rect 2137 9198 2142 9226
rect 2170 9198 4886 9226
rect 4914 9198 4919 9226
rect 6337 9198 6342 9226
rect 6370 9198 6846 9226
rect 6874 9198 7014 9226
rect 7042 9198 7047 9226
rect 7905 9198 7910 9226
rect 7938 9198 8806 9226
rect 8834 9198 8839 9226
rect 8913 9198 8918 9226
rect 8946 9198 10206 9226
rect 10234 9198 10239 9226
rect 10313 9198 10318 9226
rect 10346 9198 10766 9226
rect 10794 9198 11214 9226
rect 11242 9198 11247 9226
rect 7121 9142 7126 9170
rect 7154 9142 9422 9170
rect 9450 9142 9455 9170
rect 10145 9142 10150 9170
rect 10178 9142 10990 9170
rect 11018 9142 11023 9170
rect 11097 9142 11102 9170
rect 11130 9142 11886 9170
rect 11914 9142 11919 9170
rect 0 9114 400 9128
rect 20600 9114 21000 9128
rect 0 9086 966 9114
rect 994 9086 999 9114
rect 8745 9086 8750 9114
rect 8778 9086 9198 9114
rect 9226 9086 9646 9114
rect 9674 9086 11046 9114
rect 11074 9086 11079 9114
rect 20001 9086 20006 9114
rect 20034 9086 21000 9114
rect 0 9072 400 9086
rect 20600 9072 21000 9086
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 7065 8974 7070 9002
rect 7098 8974 7518 9002
rect 7546 8974 10262 9002
rect 10290 8974 10295 9002
rect 5721 8862 5726 8890
rect 5754 8862 6846 8890
rect 6874 8862 6879 8890
rect 12945 8862 12950 8890
rect 12978 8862 18830 8890
rect 18858 8862 18863 8890
rect 10033 8806 10038 8834
rect 10066 8806 10206 8834
rect 10234 8806 10990 8834
rect 11018 8806 11023 8834
rect 4881 8750 4886 8778
rect 4914 8750 6846 8778
rect 6874 8750 6879 8778
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 9641 8470 9646 8498
rect 9674 8470 10598 8498
rect 10626 8470 10934 8498
rect 10962 8470 11550 8498
rect 11578 8470 11583 8498
rect 6281 8358 6286 8386
rect 6314 8358 6790 8386
rect 6818 8358 6823 8386
rect 9977 8358 9982 8386
rect 10010 8358 10150 8386
rect 10178 8358 11438 8386
rect 11466 8358 11471 8386
rect 5497 8302 5502 8330
rect 5530 8302 6734 8330
rect 6762 8302 6767 8330
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 9585 8078 9590 8106
rect 9618 8078 9814 8106
rect 9842 8078 9847 8106
rect 2137 8022 2142 8050
rect 2170 8022 5614 8050
rect 5642 8022 5647 8050
rect 11153 8022 11158 8050
rect 11186 8022 11494 8050
rect 11522 8022 11527 8050
rect 9865 7966 9870 7994
rect 9898 7966 10206 7994
rect 10234 7966 10239 7994
rect 10369 7966 10374 7994
rect 10402 7966 10710 7994
rect 10738 7966 11326 7994
rect 11354 7966 11359 7994
rect 6393 7910 6398 7938
rect 6426 7910 6958 7938
rect 6986 7910 6991 7938
rect 9193 7910 9198 7938
rect 9226 7910 9702 7938
rect 9730 7910 9735 7938
rect 5609 7854 5614 7882
rect 5642 7854 6902 7882
rect 6930 7854 6935 7882
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 0 7770 400 7784
rect 0 7742 966 7770
rect 994 7742 999 7770
rect 7009 7742 7014 7770
rect 7042 7742 8918 7770
rect 8946 7742 9478 7770
rect 9506 7742 9511 7770
rect 0 7728 400 7742
rect 11265 7686 11270 7714
rect 11298 7686 11438 7714
rect 11466 7686 11471 7714
rect 2137 7630 2142 7658
rect 2170 7630 5502 7658
rect 5530 7630 5535 7658
rect 8409 7630 8414 7658
rect 8442 7630 8862 7658
rect 8890 7630 8895 7658
rect 8297 7574 8302 7602
rect 8330 7574 9030 7602
rect 9058 7574 9063 7602
rect 9697 7574 9702 7602
rect 9730 7574 10094 7602
rect 10122 7574 10127 7602
rect 11489 7574 11494 7602
rect 11522 7574 12334 7602
rect 12362 7574 12367 7602
rect 961 7518 966 7546
rect 994 7518 999 7546
rect 0 7434 400 7448
rect 966 7434 994 7518
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 0 7406 994 7434
rect 0 7392 400 7406
rect 8409 7126 8414 7154
rect 8442 7126 9198 7154
rect 9226 7126 9231 7154
rect 8745 7070 8750 7098
rect 8778 7070 9590 7098
rect 9618 7070 9623 7098
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 7457 6678 7462 6706
rect 7490 6678 8078 6706
rect 8106 6678 9646 6706
rect 9674 6678 9679 6706
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9809 6342 9814 6370
rect 9842 6342 10374 6370
rect 10402 6342 10407 6370
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 20600 5082 21000 5096
rect 20113 5054 20118 5082
rect 20146 5054 21000 5082
rect 20600 5040 21000 5054
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 8745 2590 8750 2618
rect 8778 2590 9366 2618
rect 9394 2590 9399 2618
rect 20600 2394 21000 2408
rect 20113 2366 20118 2394
rect 20146 2366 21000 2394
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 20600 2352 21000 2366
rect 9417 2030 9422 2058
rect 9450 2030 10038 2058
rect 10066 2030 10071 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 10089 1694 10094 1722
rect 10122 1694 10878 1722
rect 10906 1694 10911 1722
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _085_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10808 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _086_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10304 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _087_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9856 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _088_
timestamp 1698175906
transform -1 0 10472 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _089_
timestamp 1698175906
transform 1 0 9800 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _090_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _091_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9912 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _092_
timestamp 1698175906
transform -1 0 7896 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _093_
timestamp 1698175906
transform -1 0 8176 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _094_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9968 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _095_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 6944 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _096_
timestamp 1698175906
transform -1 0 8512 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _097_
timestamp 1698175906
transform -1 0 7504 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _098_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6496 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _099_
timestamp 1698175906
transform 1 0 8456 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _101_
timestamp 1698175906
transform 1 0 7280 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _102_
timestamp 1698175906
transform 1 0 8680 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8904 0 1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _104_
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1698175906
transform 1 0 8960 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _106_
timestamp 1698175906
transform -1 0 9240 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9128 0 -1 7840
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _108_
timestamp 1698175906
transform -1 0 8512 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _109_
timestamp 1698175906
transform -1 0 9912 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _110_
timestamp 1698175906
transform -1 0 6496 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _111_
timestamp 1698175906
transform -1 0 6048 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11536 0 1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _113_
timestamp 1698175906
transform -1 0 10640 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _114_
timestamp 1698175906
transform -1 0 10304 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform -1 0 7448 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _116_
timestamp 1698175906
transform -1 0 6608 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _117_
timestamp 1698175906
transform 1 0 6048 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8680 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _119_
timestamp 1698175906
transform -1 0 7056 0 -1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _120_
timestamp 1698175906
transform 1 0 6216 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _122_
timestamp 1698175906
transform 1 0 9744 0 1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _123_
timestamp 1698175906
transform -1 0 10920 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _124_
timestamp 1698175906
transform -1 0 10024 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _125_
timestamp 1698175906
transform -1 0 7168 0 1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _126_
timestamp 1698175906
transform 1 0 5656 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _127_
timestamp 1698175906
transform -1 0 9520 0 1 7840
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _128_
timestamp 1698175906
transform -1 0 9688 0 -1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9408 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _130_
timestamp 1698175906
transform 1 0 7784 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _131_
timestamp 1698175906
transform 1 0 8064 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _132_
timestamp 1698175906
transform -1 0 7224 0 1 7840
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _133_
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _134_
timestamp 1698175906
transform 1 0 10584 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10864 0 -1 9408
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _136_
timestamp 1698175906
transform -1 0 12824 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10920 0 -1 10976
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _138_
timestamp 1698175906
transform 1 0 9688 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _139_
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _140_
timestamp 1698175906
transform -1 0 11088 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _141_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11032 0 -1 10976
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform 1 0 12208 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _143_
timestamp 1698175906
transform 1 0 8064 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _144_
timestamp 1698175906
transform 1 0 9856 0 1 10976
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _145_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _146_
timestamp 1698175906
transform 1 0 11088 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _147_
timestamp 1698175906
transform 1 0 11312 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _148_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9912 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _149_
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _150_
timestamp 1698175906
transform 1 0 11424 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _151_
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _152_
timestamp 1698175906
transform 1 0 11648 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _153_
timestamp 1698175906
transform 1 0 11760 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _154_
timestamp 1698175906
transform -1 0 10248 0 -1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _155_
timestamp 1698175906
transform 1 0 9408 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _156_
timestamp 1698175906
transform -1 0 11368 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _157_
timestamp 1698175906
transform -1 0 11872 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _158_
timestamp 1698175906
transform 1 0 7896 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _159_
timestamp 1698175906
transform -1 0 8064 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _160_
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _161_
timestamp 1698175906
transform 1 0 9184 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _162_
timestamp 1698175906
transform 1 0 8792 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _163_
timestamp 1698175906
transform 1 0 8344 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _164_
timestamp 1698175906
transform 1 0 8568 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _165_
timestamp 1698175906
transform -1 0 7896 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _166_
timestamp 1698175906
transform 1 0 7168 0 -1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _167_
timestamp 1698175906
transform -1 0 6888 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _168_
timestamp 1698175906
transform -1 0 11592 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _169_
timestamp 1698175906
transform -1 0 11256 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _170_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7168 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _171_
timestamp 1698175906
transform 1 0 10808 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _172_
timestamp 1698175906
transform 1 0 9800 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _173_
timestamp 1698175906
transform 1 0 5992 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _174_
timestamp 1698175906
transform 1 0 6776 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _175_
timestamp 1698175906
transform 1 0 7336 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _176_
timestamp 1698175906
transform -1 0 6272 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _177_
timestamp 1698175906
transform 1 0 8848 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _178_
timestamp 1698175906
transform -1 0 6328 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _179_
timestamp 1698175906
transform -1 0 7056 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _180_
timestamp 1698175906
transform 1 0 8736 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _181_
timestamp 1698175906
transform -1 0 6440 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _182_
timestamp 1698175906
transform 1 0 7952 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _183_
timestamp 1698175906
transform 1 0 6776 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _184_
timestamp 1698175906
transform -1 0 7168 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _185_
timestamp 1698175906
transform 1 0 11424 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _186_
timestamp 1698175906
transform 1 0 11816 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _187_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11256 0 1 12544
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _188_
timestamp 1698175906
transform 1 0 11760 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _189_
timestamp 1698175906
transform 1 0 10808 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _190_
timestamp 1698175906
transform 1 0 8400 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _195_
timestamp 1698175906
transform 1 0 9576 0 1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _196_
timestamp 1698175906
transform 1 0 9240 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _197_
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _198_
timestamp 1698175906
transform 1 0 12880 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _199_
timestamp 1698175906
transform 1 0 13104 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__170__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7168 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__173__CLK
timestamp 1698175906
transform 1 0 7728 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__CLK
timestamp 1698175906
transform 1 0 6384 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__CLK
timestamp 1698175906
transform 1 0 10696 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__CLK
timestamp 1698175906
transform 1 0 6720 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__CLK
timestamp 1698175906
transform 1 0 11032 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__CLK
timestamp 1698175906
transform 1 0 8400 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__CLK
timestamp 1698175906
transform 1 0 11704 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__CLK
timestamp 1698175906
transform 1 0 11144 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__CLK
timestamp 1698175906
transform 1 0 10696 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__CLK
timestamp 1698175906
transform 1 0 10136 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 9240 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9240 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 11704 0 -1 8624
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform -1 0 11480 0 -1 11760
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_198
timestamp 1698175906
transform 1 0 11760 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_202
timestamp 1698175906
transform 1 0 11984 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_150
timestamp 1698175906
transform 1 0 9072 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_152
timestamp 1698175906
transform 1 0 9184 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_183 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10920 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_199
timestamp 1698175906
transform 1 0 11816 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 12264 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 16128 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_139
timestamp 1698175906
transform 1 0 8456 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_143
timestamp 1698175906
transform 1 0 8680 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_333
timestamp 1698175906
transform 1 0 19320 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_341
timestamp 1698175906
transform 1 0 19768 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_314
timestamp 1698175906
transform 1 0 18256 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_330
timestamp 1698175906
transform 1 0 19152 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_338
timestamp 1698175906
transform 1 0 19600 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_342
timestamp 1698175906
transform 1 0 19824 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_344
timestamp 1698175906
transform 1 0 19936 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_150
timestamp 1698175906
transform 1 0 9072 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_152
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_159
timestamp 1698175906
transform 1 0 9576 0 -1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_191
timestamp 1698175906
transform 1 0 11368 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_207
timestamp 1698175906
transform 1 0 12264 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698175906
transform 1 0 12376 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_123
timestamp 1698175906
transform 1 0 7560 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_127
timestamp 1698175906
transform 1 0 7784 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_129
timestamp 1698175906
transform 1 0 7896 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_165
timestamp 1698175906
transform 1 0 9912 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698175906
transform 1 0 10360 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_80
timestamp 1698175906
transform 1 0 5152 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_84
timestamp 1698175906
transform 1 0 5376 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_114
timestamp 1698175906
transform 1 0 7056 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_130
timestamp 1698175906
transform 1 0 7952 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_138
timestamp 1698175906
transform 1 0 8400 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_150
timestamp 1698175906
transform 1 0 9072 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_154
timestamp 1698175906
transform 1 0 9296 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_161
timestamp 1698175906
transform 1 0 9688 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_192
timestamp 1698175906
transform 1 0 11424 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698175906
transform 1 0 12320 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_115
timestamp 1698175906
transform 1 0 7112 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_156
timestamp 1698175906
transform 1 0 9408 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_164
timestamp 1698175906
transform 1 0 9856 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698175906
transform 1 0 10248 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 14168 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_28
timestamp 1698175906
transform 1 0 2240 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_60
timestamp 1698175906
transform 1 0 4032 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_68
timestamp 1698175906
transform 1 0 4480 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_80
timestamp 1698175906
transform 1 0 5152 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_84
timestamp 1698175906
transform 1 0 5376 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_86
timestamp 1698175906
transform 1 0 5488 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_116
timestamp 1698175906
transform 1 0 7168 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_132
timestamp 1698175906
transform 1 0 8064 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_151
timestamp 1698175906
transform 1 0 9128 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_155
timestamp 1698175906
transform 1 0 9352 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_164
timestamp 1698175906
transform 1 0 9856 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_172
timestamp 1698175906
transform 1 0 10304 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_180
timestamp 1698175906
transform 1 0 10752 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 16128 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_28
timestamp 1698175906
transform 1 0 2240 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698175906
transform 1 0 2464 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_69
timestamp 1698175906
transform 1 0 4536 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_85
timestamp 1698175906
transform 1 0 5432 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_93
timestamp 1698175906
transform 1 0 5880 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_97
timestamp 1698175906
transform 1 0 6104 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_103
timestamp 1698175906
transform 1 0 6440 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_117
timestamp 1698175906
transform 1 0 7224 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_158
timestamp 1698175906
transform 1 0 9520 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_162
timestamp 1698175906
transform 1 0 9744 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_195
timestamp 1698175906
transform 1 0 11592 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_227
timestamp 1698175906
transform 1 0 13384 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 14280 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_104
timestamp 1698175906
transform 1 0 6496 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_114
timestamp 1698175906
transform 1 0 7056 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_130
timestamp 1698175906
transform 1 0 7952 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698175906
transform 1 0 8400 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_146
timestamp 1698175906
transform 1 0 8848 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_197
timestamp 1698175906
transform 1 0 11704 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_205
timestamp 1698175906
transform 1 0 12152 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 12376 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 16128 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 20048 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 20160 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_69
timestamp 1698175906
transform 1 0 4536 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_85
timestamp 1698175906
transform 1 0 5432 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_93
timestamp 1698175906
transform 1 0 5880 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_116
timestamp 1698175906
transform 1 0 7168 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_148
timestamp 1698175906
transform 1 0 8960 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_156
timestamp 1698175906
transform 1 0 9408 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_158
timestamp 1698175906
transform 1 0 9520 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_165
timestamp 1698175906
transform 1 0 9912 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698175906
transform 1 0 10360 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_189
timestamp 1698175906
transform 1 0 11256 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_191
timestamp 1698175906
transform 1 0 11368 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_221
timestamp 1698175906
transform 1 0 13048 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_237
timestamp 1698175906
transform 1 0 13944 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 2240 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 4032 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 4480 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_103
timestamp 1698175906
transform 1 0 6440 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_107
timestamp 1698175906
transform 1 0 6664 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698175906
transform 1 0 8400 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_154
timestamp 1698175906
transform 1 0 9296 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_162
timestamp 1698175906
transform 1 0 9744 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_164
timestamp 1698175906
transform 1 0 9856 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_175
timestamp 1698175906
transform 1 0 10472 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_193
timestamp 1698175906
transform 1 0 11480 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 12376 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698175906
transform 1 0 16128 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 18256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 18704 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_121
timestamp 1698175906
transform 1 0 7448 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_149
timestamp 1698175906
transform 1 0 9016 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_151
timestamp 1698175906
transform 1 0 9128 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_158
timestamp 1698175906
transform 1 0 9520 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_188
timestamp 1698175906
transform 1 0 11200 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_227
timestamp 1698175906
transform 1 0 13384 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698175906
transform 1 0 14280 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 2240 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 4032 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 4480 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_106
timestamp 1698175906
transform 1 0 6608 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_110
timestamp 1698175906
transform 1 0 6832 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_126
timestamp 1698175906
transform 1 0 7728 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_134
timestamp 1698175906
transform 1 0 8176 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_138
timestamp 1698175906
transform 1 0 8400 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_203
timestamp 1698175906
transform 1 0 12040 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_207
timestamp 1698175906
transform 1 0 12264 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 12376 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_212
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_217
timestamp 1698175906
transform 1 0 12824 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_249
timestamp 1698175906
transform 1 0 14616 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_265
timestamp 1698175906
transform 1 0 15512 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_273
timestamp 1698175906
transform 1 0 15960 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698175906
transform 1 0 16184 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 16296 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 20048 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 20160 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_69
timestamp 1698175906
transform 1 0 4536 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_85
timestamp 1698175906
transform 1 0 5432 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_93
timestamp 1698175906
transform 1 0 5880 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_95
timestamp 1698175906
transform 1 0 5992 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698175906
transform 1 0 6496 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_112
timestamp 1698175906
transform 1 0 6944 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_134
timestamp 1698175906
transform 1 0 8176 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_138
timestamp 1698175906
transform 1 0 8400 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_151
timestamp 1698175906
transform 1 0 9128 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_155
timestamp 1698175906
transform 1 0 9352 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_157
timestamp 1698175906
transform 1 0 9464 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_166
timestamp 1698175906
transform 1 0 9968 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_177
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_192
timestamp 1698175906
transform 1 0 11424 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_196
timestamp 1698175906
transform 1 0 11648 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_228
timestamp 1698175906
transform 1 0 13440 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 14336 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_88
timestamp 1698175906
transform 1 0 5600 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_112
timestamp 1698175906
transform 1 0 6944 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_122
timestamp 1698175906
transform 1 0 7504 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_129
timestamp 1698175906
transform 1 0 7896 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_133
timestamp 1698175906
transform 1 0 8120 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_155
timestamp 1698175906
transform 1 0 9352 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_159
timestamp 1698175906
transform 1 0 9576 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_167
timestamp 1698175906
transform 1 0 10024 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_169
timestamp 1698175906
transform 1 0 10136 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_183
timestamp 1698175906
transform 1 0 10920 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_196
timestamp 1698175906
transform 1 0 11648 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_204
timestamp 1698175906
transform 1 0 12096 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698175906
transform 1 0 12320 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_220
timestamp 1698175906
transform 1 0 12992 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_228
timestamp 1698175906
transform 1 0 13440 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_260
timestamp 1698175906
transform 1 0 15232 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698175906
transform 1 0 16128 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 2240 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 2464 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_69
timestamp 1698175906
transform 1 0 4536 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_100
timestamp 1698175906
transform 1 0 6272 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_104
timestamp 1698175906
transform 1 0 6496 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_123
timestamp 1698175906
transform 1 0 7560 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_125
timestamp 1698175906
transform 1 0 7672 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_200
timestamp 1698175906
transform 1 0 11872 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_232
timestamp 1698175906
transform 1 0 13664 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_240
timestamp 1698175906
transform 1 0 14112 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 14336 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_88
timestamp 1698175906
transform 1 0 5600 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_92
timestamp 1698175906
transform 1 0 5824 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_94
timestamp 1698175906
transform 1 0 5936 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_124
timestamp 1698175906
transform 1 0 7616 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_128
timestamp 1698175906
transform 1 0 7840 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698175906
transform 1 0 8288 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_193
timestamp 1698175906
transform 1 0 11480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_195
timestamp 1698175906
transform 1 0 11592 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_201
timestamp 1698175906
transform 1 0 11928 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698175906
transform 1 0 16128 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 20048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 20160 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_111
timestamp 1698175906
transform 1 0 6888 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_115
timestamp 1698175906
transform 1 0 7112 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_118
timestamp 1698175906
transform 1 0 7280 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_122
timestamp 1698175906
transform 1 0 7504 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_129
timestamp 1698175906
transform 1 0 7896 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_137
timestamp 1698175906
transform 1 0 8344 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_167
timestamp 1698175906
transform 1 0 10024 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698175906
transform 1 0 10248 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_182
timestamp 1698175906
transform 1 0 10864 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_211
timestamp 1698175906
transform 1 0 12488 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 14280 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698175906
transform 1 0 5152 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_84
timestamp 1698175906
transform 1 0 5376 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_86
timestamp 1698175906
transform 1 0 5488 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_125
timestamp 1698175906
transform 1 0 7672 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_133
timestamp 1698175906
transform 1 0 8120 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_137
timestamp 1698175906
transform 1 0 8344 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 8456 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_158
timestamp 1698175906
transform 1 0 9520 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_171
timestamp 1698175906
transform 1 0 10248 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_224
timestamp 1698175906
transform 1 0 13216 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_256
timestamp 1698175906
transform 1 0 15008 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_272
timestamp 1698175906
transform 1 0 15904 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 18256 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 18704 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 2240 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 2464 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_123
timestamp 1698175906
transform 1 0 7560 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_137
timestamp 1698175906
transform 1 0 8344 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_153
timestamp 1698175906
transform 1 0 9240 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_161
timestamp 1698175906
transform 1 0 9688 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698175906
transform 1 0 10304 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 10416 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_185
timestamp 1698175906
transform 1 0 11032 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_220
timestamp 1698175906
transform 1 0 12992 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_236
timestamp 1698175906
transform 1 0 13888 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 14336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 18648 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_104
timestamp 1698175906
transform 1 0 6496 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_108
timestamp 1698175906
transform 1 0 6720 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698175906
transform 1 0 8400 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_183
timestamp 1698175906
transform 1 0 10920 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_187
timestamp 1698175906
transform 1 0 11144 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_203
timestamp 1698175906
transform 1 0 12040 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698175906
transform 1 0 12264 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 12376 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 16128 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 20048 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 20160 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_123
timestamp 1698175906
transform 1 0 7560 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_131
timestamp 1698175906
transform 1 0 8008 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_135
timestamp 1698175906
transform 1 0 8232 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_137
timestamp 1698175906
transform 1 0 8344 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_140
timestamp 1698175906
transform 1 0 8512 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_144
timestamp 1698175906
transform 1 0 8736 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_181
timestamp 1698175906
transform 1 0 10808 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698175906
transform 1 0 12208 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_6
timestamp 1698175906
transform 1 0 1008 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_168
timestamp 1698175906
transform 1 0 10080 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_195
timestamp 1698175906
transform 1 0 11592 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698175906
transform 1 0 12040 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 12768 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_243
timestamp 1698175906
transform 1 0 14280 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698175906
transform 1 0 16072 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 16296 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698175906
transform 1 0 10416 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_201
timestamp 1698175906
transform 1 0 11928 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_203
timestamp 1698175906
transform 1 0 12040 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_206
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_210
timestamp 1698175906
transform 1 0 12432 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_237
timestamp 1698175906
transform 1 0 13944 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita23_23 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 1008 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita23_24
timestamp 1698175906
transform 1 0 9240 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita23_25
timestamp 1698175906
transform 1 0 19992 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita23_26
timestamp 1698175906
transform 1 0 19992 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10192 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 12488 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 9464 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 18760 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18760 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 12824 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform -1 0 2240 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 2240 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 18760 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 10136 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform -1 0 2240 0 -1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 2240 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 10472 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform -1 0 2240 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 8792 0 1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 2240 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 10192 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13104 400 13160 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 18480 400 18536 0 FreeSans 224 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 20600 9408 21000 9464 0 FreeSans 224 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 20600 10416 21000 10472 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 12432 20600 12488 21000 0 FreeSans 224 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 10080 0 10136 400 0 FreeSans 224 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 9744 0 9800 400 0 FreeSans 224 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 20600 2352 21000 2408 0 FreeSans 224 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 9408 0 9464 400 0 FreeSans 224 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 20600 5040 21000 5096 0 FreeSans 224 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 20600 12096 21000 12152 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 20600 12432 21000 12488 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 20600 10752 21000 10808 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 12768 20600 12824 21000 0 FreeSans 224 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 9072 400 9128 0 FreeSans 224 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 7728 400 7784 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 20600 9072 21000 9128 0 FreeSans 224 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 10080 20600 10136 21000 0 FreeSans 224 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 0 7392 400 7448 0 FreeSans 224 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 0 9744 400 9800 0 FreeSans 224 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 10416 20600 10472 21000 0 FreeSans 224 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 11088 400 11144 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 8736 0 8792 400 0 FreeSans 224 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 8064 20600 8120 21000 0 FreeSans 224 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 0 12432 400 12488 0 FreeSans 224 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 9744 20600 9800 21000 0 FreeSans 224 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 6748 12180 6748 12180 0 _000_
rlabel metal2 11004 9184 11004 9184 0 _001_
rlabel metal2 10276 7028 10276 7028 0 _002_
rlabel metal2 6636 11200 6636 11200 0 _003_
rlabel metal2 7252 9380 7252 9380 0 _004_
rlabel metal2 7812 7420 7812 7420 0 _005_
rlabel metal2 5796 10920 5796 10920 0 _006_
rlabel metal2 10164 12880 10164 12880 0 _007_
rlabel metal2 5852 10080 5852 10080 0 _008_
rlabel metal2 6580 7000 6580 7000 0 _009_
rlabel metal2 9772 12908 9772 12908 0 _010_
rlabel metal2 5796 9044 5796 9044 0 _011_
rlabel metal2 8428 6832 8428 6832 0 _012_
rlabel metal2 8204 12964 8204 12964 0 _013_
rlabel metal2 6468 7462 6468 7462 0 _014_
rlabel metal2 11900 9016 11900 9016 0 _015_
rlabel metal2 12292 10584 12292 10584 0 _016_
rlabel metal2 11452 12348 11452 12348 0 _017_
rlabel metal3 11928 9660 11928 9660 0 _018_
rlabel metal2 11900 12152 11900 12152 0 _019_
rlabel metal2 9548 11340 9548 11340 0 _020_
rlabel metal2 9436 7112 9436 7112 0 _021_
rlabel metal2 8092 12684 8092 12684 0 _022_
rlabel metal3 6692 7924 6692 7924 0 _023_
rlabel metal2 10892 9212 10892 9212 0 _024_
rlabel metal3 12124 10052 12124 10052 0 _025_
rlabel metal2 10332 10780 10332 10780 0 _026_
rlabel metal2 10080 11172 10080 11172 0 _027_
rlabel metal3 10780 10444 10780 10444 0 _028_
rlabel metal2 10948 10556 10948 10556 0 _029_
rlabel metal3 12012 11956 12012 11956 0 _030_
rlabel metal3 9492 11060 9492 11060 0 _031_
rlabel metal3 10640 11116 10640 11116 0 _032_
rlabel metal2 11060 11592 11060 11592 0 _033_
rlabel metal2 11676 11984 11676 11984 0 _034_
rlabel metal2 10892 9464 10892 9464 0 _035_
rlabel metal3 11144 9492 11144 9492 0 _036_
rlabel metal2 11956 11928 11956 11928 0 _037_
rlabel metal2 11872 11676 11872 11676 0 _038_
rlabel metal2 9800 11172 9800 11172 0 _039_
rlabel metal2 10892 10248 10892 10248 0 _040_
rlabel metal3 10528 9548 10528 9548 0 _041_
rlabel metal3 8484 10332 8484 10332 0 _042_
rlabel metal2 8428 9576 8428 9576 0 _043_
rlabel metal3 9968 9604 9968 9604 0 _044_
rlabel metal2 9436 9324 9436 9324 0 _045_
rlabel metal3 11004 10780 11004 10780 0 _046_
rlabel metal3 8820 11172 8820 11172 0 _047_
rlabel metal3 8876 11284 8876 11284 0 _048_
rlabel metal3 10696 13132 10696 13132 0 _049_
rlabel metal3 7112 12012 7112 12012 0 _050_
rlabel metal2 10052 9520 10052 9520 0 _051_
rlabel metal2 10668 8428 10668 8428 0 _052_
rlabel metal3 9464 7924 9464 7924 0 _053_
rlabel metal2 9576 7196 9576 7196 0 _054_
rlabel metal3 10052 7980 10052 7980 0 _055_
rlabel metal2 9884 8092 9884 8092 0 _056_
rlabel metal2 9996 7392 9996 7392 0 _057_
rlabel metal2 8148 11004 8148 11004 0 _058_
rlabel metal2 7924 10444 7924 10444 0 _059_
rlabel metal2 8708 10640 8708 10640 0 _060_
rlabel metal2 6692 10500 6692 10500 0 _061_
rlabel metal2 9184 10052 9184 10052 0 _062_
rlabel metal2 7140 10752 7140 10752 0 _063_
rlabel metal3 10836 11172 10836 11172 0 _064_
rlabel metal2 8736 10892 8736 10892 0 _065_
rlabel metal2 8932 9352 8932 9352 0 _066_
rlabel metal2 8792 10052 8792 10052 0 _067_
rlabel metal2 9044 7406 9044 7406 0 _068_
rlabel metal2 9604 7000 9604 7000 0 _069_
rlabel metal2 9100 8988 9100 8988 0 _070_
rlabel metal3 8652 7644 8652 7644 0 _071_
rlabel metal2 11060 10696 11060 10696 0 _072_
rlabel metal3 6160 10724 6160 10724 0 _073_
rlabel metal2 10724 11788 10724 11788 0 _074_
rlabel metal2 10276 12740 10276 12740 0 _075_
rlabel metal3 6860 9548 6860 9548 0 _076_
rlabel metal2 6356 10192 6356 10192 0 _077_
rlabel metal2 8260 9688 8260 9688 0 _078_
rlabel metal2 6300 8232 6300 8232 0 _079_
rlabel metal2 10360 9548 10360 9548 0 _080_
rlabel metal2 10836 11172 10836 11172 0 _081_
rlabel metal2 9940 12880 9940 12880 0 _082_
rlabel metal3 6300 8876 6300 8876 0 _083_
rlabel metal2 9240 7812 9240 7812 0 _084_
rlabel metal2 9296 10276 9296 10276 0 clk
rlabel metal2 11732 9688 11732 9688 0 clknet_0_clk
rlabel metal2 9884 6916 9884 6916 0 clknet_1_0__leaf_clk
rlabel metal2 11816 10388 11816 10388 0 clknet_1_1__leaf_clk
rlabel metal2 11508 7784 11508 7784 0 dut23.count\[0\]
rlabel metal2 11312 8036 11312 8036 0 dut23.count\[1\]
rlabel metal2 7924 11340 7924 11340 0 dut23.count\[2\]
rlabel metal3 8932 9604 8932 9604 0 dut23.count\[3\]
rlabel metal2 9800 1764 9800 1764 0 net1
rlabel metal2 12908 16030 12908 16030 0 net10
rlabel metal2 4900 9184 4900 9184 0 net11
rlabel metal2 5628 7812 5628 7812 0 net12
rlabel metal2 18844 9044 18844 9044 0 net13
rlabel metal2 10444 17948 10444 17948 0 net14
rlabel metal3 3836 7644 3836 7644 0 net15
rlabel metal2 4788 9968 4788 9968 0 net16
rlabel metal2 10444 13580 10444 13580 0 net17
rlabel metal2 4732 11200 4732 11200 0 net18
rlabel metal2 8848 7308 8848 7308 0 net19
rlabel metal3 15960 9632 15960 9632 0 net2
rlabel metal3 8512 13076 8512 13076 0 net20
rlabel metal3 3892 12292 3892 12292 0 net21
rlabel metal2 9772 19012 9772 19012 0 net22
rlabel metal3 623 18508 623 18508 0 net23
rlabel metal2 9772 763 9772 763 0 net24
rlabel metal2 20132 2408 20132 2408 0 net25
rlabel metal2 20132 5208 20132 5208 0 net26
rlabel metal3 13048 10444 13048 10444 0 net3
rlabel metal2 12348 12432 12348 12432 0 net4
rlabel metal2 10388 4060 10388 4060 0 net5
rlabel metal2 9548 3178 9548 3178 0 net6
rlabel metal3 15960 12376 15960 12376 0 net7
rlabel metal2 18844 12628 18844 12628 0 net8
rlabel metal3 15960 10864 15960 10864 0 net9
rlabel metal2 9100 1099 9100 1099 0 segm[10]
rlabel metal2 20020 9548 20020 9548 0 segm[11]
rlabel metal2 20020 10556 20020 10556 0 segm[12]
rlabel metal2 12460 19873 12460 19873 0 segm[13]
rlabel metal2 10108 1043 10108 1043 0 segm[1]
rlabel metal2 9436 1211 9436 1211 0 segm[4]
rlabel metal2 20020 12180 20020 12180 0 segm[6]
rlabel metal2 20020 12628 20020 12628 0 segm[7]
rlabel metal2 20020 11004 20020 11004 0 segm[8]
rlabel metal2 12796 19677 12796 19677 0 segm[9]
rlabel metal3 679 9100 679 9100 0 sel[0]
rlabel metal3 679 7756 679 7756 0 sel[10]
rlabel metal3 20321 9100 20321 9100 0 sel[11]
rlabel metal2 10108 19677 10108 19677 0 sel[1]
rlabel metal3 679 7420 679 7420 0 sel[2]
rlabel metal3 679 9772 679 9772 0 sel[3]
rlabel metal2 10444 19873 10444 19873 0 sel[4]
rlabel metal3 679 11116 679 11116 0 sel[5]
rlabel metal2 8764 1491 8764 1491 0 sel[6]
rlabel metal2 8092 19677 8092 19677 0 sel[7]
rlabel metal3 679 12460 679 12460 0 sel[8]
rlabel metal2 9772 19873 9772 19873 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
