magic
tech gf180mcuD
magscale 1 5
timestamp 1699641640
<< obsm1 >>
rect 672 1538 20328 19238
<< metal2 >>
rect 7728 20600 7784 21000
rect 8064 20600 8120 21000
rect 9408 20600 9464 21000
rect 10416 20600 10472 21000
rect 12096 20600 12152 21000
rect 13104 20600 13160 21000
rect 8400 0 8456 400
rect 10752 0 10808 400
rect 11760 0 11816 400
rect 12432 0 12488 400
rect 12768 0 12824 400
<< obsm2 >>
rect 966 20570 7698 20600
rect 7814 20570 8034 20600
rect 8150 20570 9378 20600
rect 9494 20570 10386 20600
rect 10502 20570 12066 20600
rect 12182 20570 13074 20600
rect 13190 20570 20034 20600
rect 966 430 20034 20570
rect 966 400 8370 430
rect 8486 400 10722 430
rect 10838 400 11730 430
rect 11846 400 12402 430
rect 12518 400 12738 430
rect 12854 400 20034 430
<< metal3 >>
rect 20600 13776 21000 13832
rect 0 13440 400 13496
rect 0 12432 400 12488
rect 20600 12432 21000 12488
rect 0 12096 400 12152
rect 0 11760 400 11816
rect 20600 11760 21000 11816
rect 0 11424 400 11480
rect 20600 10752 21000 10808
rect 0 10416 400 10472
rect 20600 10080 21000 10136
rect 0 9744 400 9800
rect 20600 8736 21000 8792
rect 0 8400 400 8456
rect 20600 8400 21000 8456
rect 20600 7392 21000 7448
<< obsm3 >>
rect 400 13862 20600 19222
rect 400 13746 20570 13862
rect 400 13526 20600 13746
rect 430 13410 20600 13526
rect 400 12518 20600 13410
rect 430 12402 20570 12518
rect 400 12182 20600 12402
rect 430 12066 20600 12182
rect 400 11846 20600 12066
rect 430 11730 20570 11846
rect 400 11510 20600 11730
rect 430 11394 20600 11510
rect 400 10838 20600 11394
rect 400 10722 20570 10838
rect 400 10502 20600 10722
rect 430 10386 20600 10502
rect 400 10166 20600 10386
rect 400 10050 20570 10166
rect 400 9830 20600 10050
rect 430 9714 20600 9830
rect 400 8822 20600 9714
rect 400 8706 20570 8822
rect 400 8486 20600 8706
rect 430 8370 20570 8486
rect 400 7478 20600 8370
rect 400 7362 20570 7478
rect 400 1554 20600 7362
<< metal4 >>
rect 2224 1538 2384 19238
rect 9904 1538 10064 19238
rect 17584 1538 17744 19238
<< labels >>
rlabel metal3 s 0 13440 400 13496 6 clk
port 1 nsew signal input
rlabel metal2 s 7728 20600 7784 21000 6 segm[0]
port 2 nsew signal output
rlabel metal3 s 0 12432 400 12488 6 segm[10]
port 3 nsew signal output
rlabel metal2 s 12432 0 12488 400 6 segm[11]
port 4 nsew signal output
rlabel metal3 s 20600 11760 21000 11816 6 segm[12]
port 5 nsew signal output
rlabel metal2 s 10416 20600 10472 21000 6 segm[13]
port 6 nsew signal output
rlabel metal3 s 0 10416 400 10472 6 segm[1]
port 7 nsew signal output
rlabel metal3 s 20600 8400 21000 8456 6 segm[2]
port 8 nsew signal output
rlabel metal3 s 20600 13776 21000 13832 6 segm[3]
port 9 nsew signal output
rlabel metal3 s 0 9744 400 9800 6 segm[4]
port 10 nsew signal output
rlabel metal3 s 20600 8736 21000 8792 6 segm[5]
port 11 nsew signal output
rlabel metal3 s 20600 10080 21000 10136 6 segm[6]
port 12 nsew signal output
rlabel metal3 s 0 11424 400 11480 6 segm[7]
port 13 nsew signal output
rlabel metal3 s 0 12096 400 12152 6 segm[8]
port 14 nsew signal output
rlabel metal3 s 0 11760 400 11816 6 segm[9]
port 15 nsew signal output
rlabel metal2 s 8400 0 8456 400 6 sel[0]
port 16 nsew signal output
rlabel metal2 s 10752 0 10808 400 6 sel[10]
port 17 nsew signal output
rlabel metal2 s 8064 20600 8120 21000 6 sel[11]
port 18 nsew signal output
rlabel metal3 s 20600 12432 21000 12488 6 sel[1]
port 19 nsew signal output
rlabel metal2 s 13104 20600 13160 21000 6 sel[2]
port 20 nsew signal output
rlabel metal3 s 20600 10752 21000 10808 6 sel[3]
port 21 nsew signal output
rlabel metal2 s 12096 20600 12152 21000 6 sel[4]
port 22 nsew signal output
rlabel metal3 s 0 8400 400 8456 6 sel[5]
port 23 nsew signal output
rlabel metal2 s 9408 20600 9464 21000 6 sel[6]
port 24 nsew signal output
rlabel metal3 s 20600 7392 21000 7448 6 sel[7]
port 25 nsew signal output
rlabel metal2 s 11760 0 11816 400 6 sel[8]
port 26 nsew signal output
rlabel metal2 s 12768 0 12824 400 6 sel[9]
port 27 nsew signal output
rlabel metal4 s 2224 1538 2384 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 19238 6 vss
port 29 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 21000 21000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 525342
string GDS_FILE /home/urielcho/Proyectos_caravel/ITA23_GFMPW1b/openlane/ita21/runs/23_11_10_12_38/results/signoff/ita21.magic.gds
string GDS_START 168910
<< end >>

