* NGSPICE file created from ita24.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

.subckt ita24 clk segm[10] segm[11] segm[12] segm[13] segm[1] segm[2] segm[4] segm[5]
+ segm[6] segm[7] segm[8] segm[9] sel[0] sel[10] sel[11] sel[1] sel[2] sel[3] sel[4]
+ sel[5] sel[6] sel[7] sel[8] sel[9] vdd vss segm[3] segm[0]
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_15_Left_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_37_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_14_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_0_Left_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_42_Left_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_131_ _082_ _086_ _087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_200_ _102_ _051_ _058_ _095_ _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_31_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_114_ _071_ _072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__224__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput20 net20 sel[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput7 net7 segm[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_9_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_130_ _071_ _086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_31_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_113_ dut24.count\[2\] _071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput8 net8 segm[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput10 net10 segm[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput21 net21 sel[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__214__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_9_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_28_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_189_ _068_ _069_ _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_112_ _001_ _069_ _070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_18_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput11 net11 segm[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput22 net22 sel[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput9 net9 segm[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_41_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_17_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_19_Left_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__227__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_4_Left_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_188_ _050_ _016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_111_ dut24.count\[1\] _069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_7_Left_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput23 net23 sel[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_33_Left_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput12 net12 segm[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_1_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_36_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_34_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Left_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_187_ _038_ _048_ _049_ _050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_0_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__217__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_110_ _068_ _001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput24 net24 sel[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput13 net13 sel[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_17_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_8_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_186_ _086_ _070_ _033_ _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_30_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_169_ _032_ _034_ _036_ _011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__207__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput14 net14 sel[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_17_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_8_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_185_ net4 _074_ _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_42_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_44_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_168_ _035_ _093_ _036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput15 net15 sel[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_184_ _045_ _046_ _047_ _041_ _015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_24_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_167_ _088_ _062_ _096_ _033_ _035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_7_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_27_Left_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_11_Left_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_219_ _011_ clknet_1_0__leaf_clk net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__230__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput16 net16 sel[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_34_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_clk clk clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_42_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_25_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_183_ net1 _074_ _047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_41_Left_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_30_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_235_ net8 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_166_ _062_ _030_ _033_ net12 _034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_21_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_149_ _073_ _100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_218_ _010_ clknet_1_1__leaf_clk net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput17 net17 sel[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__220__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_42_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_10_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_182_ _035_ _097_ _046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_234_ net10 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_165_ dut24.count\[3\] _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_217_ _009_ clknet_1_0__leaf_clk net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_148_ net19 _085_ _099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput18 net18 sel[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_20_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_42_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_10_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__210__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_181_ _039_ _078_ _043_ _045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_0_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_164_ _062_ _066_ _032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_233_ net7 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_147_ _097_ _098_ _005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_216_ _008_ clknet_1_0__leaf_clk net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput19 net19 sel[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_22_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_27_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_180_ _041_ _042_ _043_ _044_ _014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XPHY_EDGE_ROW_18_Left_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_3_Left_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_163_ _101_ _031_ _087_ _010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__223__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_146_ net20 _080_ _098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_215_ _007_ clknet_1_0__leaf_clk net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_6_Left_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_129_ _082_ _085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_16_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_32_Left_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_22_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_10_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_35_Left_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_162_ net13 _030_ _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_0_clk_I clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_145_ _088_ _089_ _094_ _096_ _097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_214_ _006_ clknet_1_1__leaf_clk net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__213__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_128_ _083_ _077_ _084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_16_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_39_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xita24_25 segm[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_32_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_230_ _022_ clknet_1_1__leaf_clk net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_161_ _096_ _030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_213_ _005_ clknet_1_1__leaf_clk net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_144_ _065_ _096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_127_ _082_ _072_ _083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__226__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xita24_26 segm[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_1_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_160_ _029_ _009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_143_ _095_ _076_ _078_ _004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_212_ _004_ clknet_1_1__leaf_clk dut24.count\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_126_ dut24.count\[3\] _082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_7_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_109_ dut24.count\[0\] _068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_13_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_24_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_39_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__216__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_23_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_211_ _003_ clknet_1_0__leaf_clk dut24.count\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_142_ _094_ _095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_19_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_125_ _078_ _081_ _024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_26_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_10_Left_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_36_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_108_ _066_ _067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_13_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_40_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_141_ _063_ _094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_210_ _002_ clknet_1_0__leaf_clk dut24.count\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_19_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_124_ net22 _080_ _081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__206__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__229__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_107_ _064_ _065_ _066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_13_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_140_ _067_ _093_ _003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_123_ _079_ _080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_106_ dut24.count\[2\] _065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_13_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_4_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__219__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_199_ net15 _102_ _058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_122_ _064_ _071_ _079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_105_ _063_ _064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_14_Left_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_27_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_32_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_17_Left_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__209__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_2_Left_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_198_ _088_ _032_ _057_ _019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_44_Left_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_121_ _077_ _078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_1_0__f_clk clknet_0_clk clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_104_ dut24.count\[3\] _063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_5_Left_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_31_Left_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_197_ net14 _085_ _030_ _057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_42_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_120_ _064_ _065_ _076_ _077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_16_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_103_ dut24.count\[1\] _062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_44_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_4_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_196_ _083_ _078_ _043_ _056_ _018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_179_ _087_ _092_ _044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_16_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_35_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_23_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__222__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_195_ net3 _085_ _056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_178_ _002_ _025_ _043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_7_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_12_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_9_Left_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_38_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_22_Left_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_194_ _095_ _054_ _055_ _084_ _017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_177_ net10 _074_ _042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__212__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_44_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_229_ _021_ clknet_1_1__leaf_clk net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_25_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_193_ net7 _094_ _055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_18_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_176_ _083_ _100_ _041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_7_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_159_ net16 _079_ _025_ _070_ _029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_228_ _020_ clknet_1_1__leaf_clk net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_26_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__225__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_192_ _052_ _053_ _054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_175_ _039_ _040_ _013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_158_ _027_ _028_ _008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_227_ _019_ clknet_1_0__leaf_clk net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_43_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_1_1__f_clk clknet_0_clk clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_25_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__215__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_191_ _096_ _092_ _053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_174_ net8 _080_ _040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_15_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_157_ net17 _080_ _028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_226_ _018_ clknet_1_1__leaf_clk net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_43_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_29_Left_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_13_Left_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_209_ _001_ clknet_1_0__leaf_clk dut24.count\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_16_Left_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_190_ _086_ _051_ _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_173_ _082_ _086_ _073_ _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_1_Left_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_43_Left_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_156_ _090_ _025_ _027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_225_ _017_ clknet_1_1__leaf_clk net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__228__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_139_ _072_ _076_ _093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_208_ _000_ clknet_1_1__leaf_clk net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_30_Left_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_172_ _027_ _037_ _038_ _012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_23_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_224_ _016_ clknet_1_0__leaf_clk net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_155_ _026_ _007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_6_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_26_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_207_ _024_ clknet_1_1__leaf_clk net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_138_ _092_ _002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__218__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_171_ _083_ _100_ _038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_38_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_223_ _015_ clknet_1_1__leaf_clk net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_154_ net18 _079_ _025_ _076_ _026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_40_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_206_ _023_ clknet_1_0__leaf_clk net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_137_ dut24.count\[0\] dut24.count\[1\] _092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_43_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__208__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput1 net1 segm[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_170_ net6 _033_ _067_ _100_ _037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_29_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_222_ _014_ clknet_1_1__leaf_clk net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_153_ dut24.count\[3\] _065_ _025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_20_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_40_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_136_ _084_ _091_ _000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_205_ _049_ _053_ _060_ _061_ _022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_8_Left_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_119_ _068_ dut24.count\[1\] _076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_34_Left_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput2 net2 segm[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_37_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_21_Left_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_29_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_221_ _013_ clknet_1_1__leaf_clk net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_152_ _099_ _101_ _102_ _006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_34_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_204_ net2 _030_ _061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_40_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_135_ net21 _085_ _087_ _090_ _091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_118_ _062_ _067_ _075_ _023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_24_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput3 net3 segm[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_18_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_220_ _012_ clknet_1_1__leaf_clk net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_151_ _072_ _102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_6_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_134_ _088_ _089_ _090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_203_ _102_ _051_ _095_ _060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_117_ _067_ _070_ _074_ net24 _075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_39_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput4 net4 segm[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__221__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_150_ _094_ _100_ _101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_40_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_202_ _052_ _044_ _059_ _021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_25_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_133_ _069_ _089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_31_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_116_ _072_ _073_ _064_ _074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_0_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput5 net5 segm[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_37_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_14_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__211__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_201_ net11 _079_ _059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_25_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_132_ dut24.count\[0\] _088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_31_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_115_ _068_ _069_ _073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_12_Left_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput6 net6 segm[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_26_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
.ends

