magic
tech gf180mcuD
magscale 1 5
timestamp 1699641280
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9311 19137 9337 19143
rect 9311 19105 9337 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 11097 19055 11103 19081
rect 11129 19055 11135 19081
rect 9025 18999 9031 19025
rect 9057 18999 9063 19025
rect 11769 18999 11775 19025
rect 11801 18999 11807 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 10599 18913 10625 18919
rect 10599 18881 10625 18887
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 9927 18745 9953 18751
rect 9927 18713 9953 18719
rect 11383 18745 11409 18751
rect 11383 18713 11409 18719
rect 20119 18689 20145 18695
rect 20119 18657 20145 18663
rect 9417 18607 9423 18633
rect 9449 18607 9455 18633
rect 10985 18607 10991 18633
rect 11017 18607 11023 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 9031 18353 9057 18359
rect 9031 18321 9057 18327
rect 8521 18215 8527 18241
rect 8553 18215 8559 18241
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 7911 14041 7937 14047
rect 7911 14009 7937 14015
rect 8359 14041 8385 14047
rect 8359 14009 8385 14015
rect 10151 14041 10177 14047
rect 10151 14009 10177 14015
rect 7967 13929 7993 13935
rect 8129 13903 8135 13929
rect 8161 13903 8167 13929
rect 8241 13903 8247 13929
rect 8273 13903 8279 13929
rect 10257 13903 10263 13929
rect 10289 13903 10295 13929
rect 7967 13897 7993 13903
rect 8191 13873 8217 13879
rect 10649 13847 10655 13873
rect 10681 13847 10687 13873
rect 11713 13847 11719 13873
rect 11745 13847 11751 13873
rect 8191 13841 8217 13847
rect 7911 13817 7937 13823
rect 7911 13785 7937 13791
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 11047 13649 11073 13655
rect 11047 13617 11073 13623
rect 20007 13593 20033 13599
rect 9081 13567 9087 13593
rect 9113 13567 9119 13593
rect 13673 13567 13679 13593
rect 13705 13567 13711 13593
rect 20007 13561 20033 13567
rect 11103 13537 11129 13543
rect 7625 13511 7631 13537
rect 7657 13511 7663 13537
rect 12273 13511 12279 13537
rect 12305 13511 12311 13537
rect 18825 13511 18831 13537
rect 18857 13511 18863 13537
rect 11103 13505 11129 13511
rect 8017 13455 8023 13481
rect 8049 13455 8055 13481
rect 12609 13455 12615 13481
rect 12641 13455 12647 13481
rect 9311 13425 9337 13431
rect 9311 13393 9337 13399
rect 13903 13425 13929 13431
rect 13903 13393 13929 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 8919 13257 8945 13263
rect 8919 13225 8945 13231
rect 9143 13257 9169 13263
rect 9143 13225 9169 13231
rect 11383 13257 11409 13263
rect 11383 13225 11409 13231
rect 11439 13257 11465 13263
rect 11439 13225 11465 13231
rect 13231 13257 13257 13263
rect 13231 13225 13257 13231
rect 11495 13201 11521 13207
rect 7345 13175 7351 13201
rect 7377 13175 7383 13201
rect 11495 13169 11521 13175
rect 11327 13145 11353 13151
rect 13119 13145 13145 13151
rect 2137 13119 2143 13145
rect 2169 13119 2175 13145
rect 7009 13119 7015 13145
rect 7041 13119 7047 13145
rect 8689 13119 8695 13145
rect 8721 13119 8727 13145
rect 8801 13119 8807 13145
rect 8833 13119 8839 13145
rect 9641 13119 9647 13145
rect 9673 13119 9679 13145
rect 11713 13119 11719 13145
rect 11745 13119 11751 13145
rect 11327 13113 11353 13119
rect 13119 13113 13145 13119
rect 13287 13145 13313 13151
rect 13897 13119 13903 13145
rect 13929 13119 13935 13145
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 13287 13113 13313 13119
rect 15583 13089 15609 13095
rect 8409 13063 8415 13089
rect 8441 13063 8447 13089
rect 9977 13063 9983 13089
rect 10009 13063 10015 13089
rect 11041 13063 11047 13089
rect 11073 13063 11079 13089
rect 14289 13063 14295 13089
rect 14321 13063 14327 13089
rect 15353 13063 15359 13089
rect 15385 13063 15391 13089
rect 19945 13063 19951 13089
rect 19977 13063 19983 13089
rect 15583 13057 15609 13063
rect 967 13033 993 13039
rect 967 13001 993 13007
rect 8751 13033 8777 13039
rect 8751 13001 8777 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 10655 12865 10681 12871
rect 10655 12833 10681 12839
rect 14127 12865 14153 12871
rect 14127 12833 14153 12839
rect 7687 12809 7713 12815
rect 7687 12777 7713 12783
rect 11159 12809 11185 12815
rect 11159 12777 11185 12783
rect 12783 12809 12809 12815
rect 12783 12777 12809 12783
rect 20007 12809 20033 12815
rect 20007 12777 20033 12783
rect 7799 12753 7825 12759
rect 7799 12721 7825 12727
rect 8415 12753 8441 12759
rect 8415 12721 8441 12727
rect 8583 12753 8609 12759
rect 8583 12721 8609 12727
rect 13119 12753 13145 12759
rect 13119 12721 13145 12727
rect 14239 12753 14265 12759
rect 14239 12721 14265 12727
rect 14743 12753 14769 12759
rect 18825 12727 18831 12753
rect 18857 12727 18863 12753
rect 14743 12721 14769 12727
rect 10711 12697 10737 12703
rect 10711 12665 10737 12671
rect 12839 12697 12865 12703
rect 12839 12665 12865 12671
rect 12951 12697 12977 12703
rect 12951 12665 12977 12671
rect 14575 12697 14601 12703
rect 14575 12665 14601 12671
rect 14631 12697 14657 12703
rect 14631 12665 14657 12671
rect 7519 12641 7545 12647
rect 7519 12609 7545 12615
rect 7631 12641 7657 12647
rect 7631 12609 7657 12615
rect 8527 12641 8553 12647
rect 8527 12609 8553 12615
rect 13063 12641 13089 12647
rect 13063 12609 13089 12615
rect 13959 12641 13985 12647
rect 13959 12609 13985 12615
rect 14071 12641 14097 12647
rect 14071 12609 14097 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 8975 12473 9001 12479
rect 8689 12447 8695 12473
rect 8721 12447 8727 12473
rect 8975 12441 9001 12447
rect 10767 12473 10793 12479
rect 11321 12447 11327 12473
rect 11353 12447 11359 12473
rect 10767 12441 10793 12447
rect 9087 12417 9113 12423
rect 11159 12417 11185 12423
rect 11041 12391 11047 12417
rect 11073 12391 11079 12417
rect 9087 12385 9113 12391
rect 11159 12385 11185 12391
rect 8863 12361 8889 12367
rect 7569 12335 7575 12361
rect 7601 12335 7607 12361
rect 8863 12329 8889 12335
rect 9143 12361 9169 12367
rect 9143 12329 9169 12335
rect 10711 12361 10737 12367
rect 11433 12335 11439 12361
rect 11465 12335 11471 12361
rect 12665 12335 12671 12361
rect 12697 12335 12703 12361
rect 14289 12335 14295 12361
rect 14321 12335 14327 12361
rect 10711 12329 10737 12335
rect 7799 12305 7825 12311
rect 6113 12279 6119 12305
rect 6145 12279 6151 12305
rect 7177 12279 7183 12305
rect 7209 12279 7215 12305
rect 7799 12273 7825 12279
rect 10823 12305 10849 12311
rect 15919 12305 15945 12311
rect 13001 12279 13007 12305
rect 13033 12279 13039 12305
rect 14065 12279 14071 12305
rect 14097 12279 14103 12305
rect 14625 12279 14631 12305
rect 14657 12279 14663 12305
rect 15689 12279 15695 12305
rect 15721 12279 15727 12305
rect 10823 12273 10849 12279
rect 15919 12273 15945 12279
rect 10935 12249 10961 12255
rect 10935 12217 10961 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 7631 12081 7657 12087
rect 7631 12049 7657 12055
rect 10991 12081 11017 12087
rect 10991 12049 11017 12055
rect 13343 12081 13369 12087
rect 13343 12049 13369 12055
rect 14183 12081 14209 12087
rect 14183 12049 14209 12055
rect 7351 12025 7377 12031
rect 13847 12025 13873 12031
rect 13001 11999 13007 12025
rect 13033 11999 13039 12025
rect 7351 11993 7377 11999
rect 13847 11993 13873 11999
rect 20007 12025 20033 12031
rect 20007 11993 20033 11999
rect 7239 11969 7265 11975
rect 6729 11943 6735 11969
rect 6761 11943 6767 11969
rect 7239 11937 7265 11943
rect 7575 11969 7601 11975
rect 7575 11937 7601 11943
rect 10823 11969 10849 11975
rect 12279 11969 12305 11975
rect 11265 11943 11271 11969
rect 11297 11943 11303 11969
rect 11601 11943 11607 11969
rect 11633 11943 11639 11969
rect 10823 11937 10849 11943
rect 12279 11937 12305 11943
rect 12839 11969 12865 11975
rect 12839 11937 12865 11943
rect 14295 11969 14321 11975
rect 14295 11937 14321 11943
rect 14575 11969 14601 11975
rect 14575 11937 14601 11943
rect 14743 11969 14769 11975
rect 18825 11943 18831 11969
rect 18857 11943 18863 11969
rect 14743 11937 14769 11943
rect 6903 11913 6929 11919
rect 6903 11881 6929 11887
rect 9199 11913 9225 11919
rect 9199 11881 9225 11887
rect 10711 11913 10737 11919
rect 12447 11913 12473 11919
rect 11153 11887 11159 11913
rect 11185 11887 11191 11913
rect 10711 11881 10737 11887
rect 12447 11881 12473 11887
rect 13119 11913 13145 11919
rect 13119 11881 13145 11887
rect 13287 11913 13313 11919
rect 13287 11881 13313 11887
rect 14015 11913 14041 11919
rect 14015 11881 14041 11887
rect 14631 11913 14657 11919
rect 14631 11881 14657 11887
rect 6847 11857 6873 11863
rect 6847 11825 6873 11831
rect 7183 11857 7209 11863
rect 12391 11857 12417 11863
rect 9025 11831 9031 11857
rect 9057 11831 9063 11857
rect 11489 11831 11495 11857
rect 11521 11831 11527 11857
rect 7183 11825 7209 11831
rect 12391 11825 12417 11831
rect 13007 11857 13033 11863
rect 13007 11825 13033 11831
rect 13343 11857 13369 11863
rect 13343 11825 13369 11831
rect 14127 11857 14153 11863
rect 14127 11825 14153 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 9255 11689 9281 11695
rect 9255 11657 9281 11663
rect 12055 11689 12081 11695
rect 12055 11657 12081 11663
rect 12839 11689 12865 11695
rect 12839 11657 12865 11663
rect 8863 11633 8889 11639
rect 8863 11601 8889 11607
rect 12895 11633 12921 11639
rect 12895 11601 12921 11607
rect 7575 11577 7601 11583
rect 2137 11551 2143 11577
rect 2169 11551 2175 11577
rect 7289 11551 7295 11577
rect 7321 11551 7327 11577
rect 7457 11551 7463 11577
rect 7489 11551 7495 11577
rect 7575 11545 7601 11551
rect 7687 11577 7713 11583
rect 8639 11577 8665 11583
rect 7793 11551 7799 11577
rect 7825 11551 7831 11577
rect 7687 11545 7713 11551
rect 8639 11545 8665 11551
rect 8919 11577 8945 11583
rect 8919 11545 8945 11551
rect 9143 11577 9169 11583
rect 9143 11545 9169 11551
rect 9199 11577 9225 11583
rect 9199 11545 9225 11551
rect 9479 11577 9505 11583
rect 11607 11577 11633 11583
rect 11321 11551 11327 11577
rect 11353 11551 11359 11577
rect 11489 11551 11495 11577
rect 11521 11551 11527 11577
rect 9479 11545 9505 11551
rect 11607 11545 11633 11551
rect 11719 11577 11745 11583
rect 11719 11545 11745 11551
rect 11775 11577 11801 11583
rect 11775 11545 11801 11551
rect 12783 11577 12809 11583
rect 13001 11551 13007 11577
rect 13033 11551 13039 11577
rect 13169 11551 13175 11577
rect 13201 11551 13207 11577
rect 12783 11545 12809 11551
rect 7631 11521 7657 11527
rect 5833 11495 5839 11521
rect 5865 11495 5871 11521
rect 6897 11495 6903 11521
rect 6929 11495 6935 11521
rect 7631 11489 7657 11495
rect 8023 11521 8049 11527
rect 8023 11489 8049 11495
rect 8751 11521 8777 11527
rect 11663 11521 11689 11527
rect 9865 11495 9871 11521
rect 9897 11495 9903 11521
rect 10929 11495 10935 11521
rect 10961 11495 10967 11521
rect 8751 11489 8777 11495
rect 11663 11489 11689 11495
rect 967 11465 993 11471
rect 967 11433 993 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 6903 11297 6929 11303
rect 6903 11265 6929 11271
rect 13119 11297 13145 11303
rect 13119 11265 13145 11271
rect 967 11241 993 11247
rect 7519 11241 7545 11247
rect 9759 11241 9785 11247
rect 6785 11215 6791 11241
rect 6817 11215 6823 11241
rect 8465 11215 8471 11241
rect 8497 11215 8503 11241
rect 9529 11215 9535 11241
rect 9561 11215 9567 11241
rect 967 11209 993 11215
rect 7519 11209 7545 11215
rect 9759 11209 9785 11215
rect 10935 11241 10961 11247
rect 20007 11241 20033 11247
rect 13617 11215 13623 11241
rect 13649 11215 13655 11241
rect 10935 11209 10961 11215
rect 20007 11209 20033 11215
rect 7407 11185 7433 11191
rect 2137 11159 2143 11185
rect 2169 11159 2175 11185
rect 7407 11153 7433 11159
rect 7575 11185 7601 11191
rect 10879 11185 10905 11191
rect 7681 11159 7687 11185
rect 7713 11159 7719 11185
rect 8073 11159 8079 11185
rect 8105 11159 8111 11185
rect 7575 11153 7601 11159
rect 10879 11153 10905 11159
rect 11159 11185 11185 11191
rect 11159 11153 11185 11159
rect 11551 11185 11577 11191
rect 11551 11153 11577 11159
rect 11719 11185 11745 11191
rect 11719 11153 11745 11159
rect 13063 11185 13089 11191
rect 13063 11153 13089 11159
rect 13847 11185 13873 11191
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 13847 11153 13873 11159
rect 11047 11129 11073 11135
rect 10089 11103 10095 11129
rect 10121 11103 10127 11129
rect 11047 11097 11073 11103
rect 13567 11129 13593 11135
rect 13567 11097 13593 11103
rect 6791 11073 6817 11079
rect 6791 11041 6817 11047
rect 7463 11073 7489 11079
rect 7463 11041 7489 11047
rect 10263 11073 10289 11079
rect 10263 11041 10289 11047
rect 11439 11073 11465 11079
rect 11439 11041 11465 11047
rect 11607 11073 11633 11079
rect 11607 11041 11633 11047
rect 11999 11073 12025 11079
rect 12671 11073 12697 11079
rect 13119 11073 13145 11079
rect 12161 11047 12167 11073
rect 12193 11047 12199 11073
rect 12833 11047 12839 11073
rect 12865 11047 12871 11073
rect 11999 11041 12025 11047
rect 12671 11041 12697 11047
rect 13119 11041 13145 11047
rect 13679 11073 13705 11079
rect 13679 11041 13705 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 7799 10905 7825 10911
rect 7799 10873 7825 10879
rect 11719 10905 11745 10911
rect 11719 10873 11745 10879
rect 13455 10905 13481 10911
rect 13455 10873 13481 10879
rect 12895 10849 12921 10855
rect 6841 10823 6847 10849
rect 6873 10823 6879 10849
rect 7625 10823 7631 10849
rect 7657 10823 7663 10849
rect 9753 10823 9759 10849
rect 9785 10823 9791 10849
rect 12895 10817 12921 10823
rect 12951 10849 12977 10855
rect 12951 10817 12977 10823
rect 13511 10849 13537 10855
rect 14401 10823 14407 10849
rect 14433 10823 14439 10849
rect 13511 10817 13537 10823
rect 7463 10793 7489 10799
rect 11663 10793 11689 10799
rect 7233 10767 7239 10793
rect 7265 10767 7271 10793
rect 11489 10767 11495 10793
rect 11521 10767 11527 10793
rect 7463 10761 7489 10767
rect 11663 10761 11689 10767
rect 11831 10793 11857 10799
rect 11831 10761 11857 10767
rect 11943 10793 11969 10799
rect 11943 10761 11969 10767
rect 12783 10793 12809 10799
rect 13343 10793 13369 10799
rect 13113 10767 13119 10793
rect 13145 10767 13151 10793
rect 13673 10767 13679 10793
rect 13705 10767 13711 10793
rect 14009 10767 14015 10793
rect 14041 10767 14047 10793
rect 12783 10761 12809 10767
rect 13343 10761 13369 10767
rect 15695 10737 15721 10743
rect 5777 10711 5783 10737
rect 5809 10711 5815 10737
rect 13169 10711 13175 10737
rect 13201 10711 13207 10737
rect 13729 10711 13735 10737
rect 13761 10711 13767 10737
rect 15465 10711 15471 10737
rect 15497 10711 15503 10737
rect 15695 10705 15721 10711
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 967 10457 993 10463
rect 967 10425 993 10431
rect 20007 10457 20033 10463
rect 20007 10425 20033 10431
rect 7911 10401 7937 10407
rect 2137 10375 2143 10401
rect 2169 10375 2175 10401
rect 7911 10369 7937 10375
rect 9759 10401 9785 10407
rect 13455 10401 13481 10407
rect 10257 10375 10263 10401
rect 10289 10375 10295 10401
rect 10649 10375 10655 10401
rect 10681 10375 10687 10401
rect 13841 10375 13847 10401
rect 13873 10375 13879 10401
rect 18825 10375 18831 10401
rect 18857 10375 18863 10401
rect 9759 10369 9785 10375
rect 13455 10369 13481 10375
rect 6735 10345 6761 10351
rect 6735 10313 6761 10319
rect 7631 10345 7657 10351
rect 7631 10313 7657 10319
rect 7743 10345 7769 10351
rect 8807 10345 8833 10351
rect 8409 10319 8415 10345
rect 8441 10319 8447 10345
rect 7743 10313 7769 10319
rect 8807 10313 8833 10319
rect 9871 10345 9897 10351
rect 9871 10313 9897 10319
rect 10039 10345 10065 10351
rect 13567 10345 13593 10351
rect 10369 10319 10375 10345
rect 10401 10319 10407 10345
rect 12553 10319 12559 10345
rect 12585 10319 12591 10345
rect 10039 10313 10065 10319
rect 13567 10313 13593 10319
rect 13623 10345 13649 10351
rect 13623 10313 13649 10319
rect 6791 10289 6817 10295
rect 6791 10257 6817 10263
rect 6847 10289 6873 10295
rect 6847 10257 6873 10263
rect 7799 10289 7825 10295
rect 7799 10257 7825 10263
rect 8583 10289 8609 10295
rect 8583 10257 8609 10263
rect 8975 10289 9001 10295
rect 8975 10257 9001 10263
rect 13511 10289 13537 10295
rect 13511 10257 13537 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 10823 10121 10849 10127
rect 10823 10089 10849 10095
rect 11159 10121 11185 10127
rect 11159 10089 11185 10095
rect 12223 10121 12249 10127
rect 12223 10089 12249 10095
rect 9031 10065 9057 10071
rect 10151 10065 10177 10071
rect 6337 10039 6343 10065
rect 6369 10039 6375 10065
rect 7289 10039 7295 10065
rect 7321 10039 7327 10065
rect 9473 10039 9479 10065
rect 9505 10039 9511 10065
rect 9031 10033 9057 10039
rect 10151 10033 10177 10039
rect 10207 10065 10233 10071
rect 10207 10033 10233 10039
rect 12279 10065 12305 10071
rect 12279 10033 12305 10039
rect 15415 10065 15441 10071
rect 15415 10033 15441 10039
rect 9647 10009 9673 10015
rect 6729 9983 6735 10009
rect 6761 9983 6767 10009
rect 6953 9983 6959 10009
rect 6985 9983 6991 10009
rect 9647 9977 9673 9983
rect 10095 10009 10121 10015
rect 10095 9977 10121 9983
rect 10431 10009 10457 10015
rect 10431 9977 10457 9983
rect 10655 10009 10681 10015
rect 10655 9977 10681 9983
rect 10767 10009 10793 10015
rect 10767 9977 10793 9983
rect 10991 10009 11017 10015
rect 10991 9977 11017 9983
rect 11103 10009 11129 10015
rect 11103 9977 11129 9983
rect 11271 10009 11297 10015
rect 11937 9983 11943 10009
rect 11969 9983 11975 10009
rect 12609 9983 12615 10009
rect 12641 9983 12647 10009
rect 11271 9977 11297 9983
rect 8751 9953 8777 9959
rect 15471 9953 15497 9959
rect 5273 9927 5279 9953
rect 5305 9927 5311 9953
rect 8353 9927 8359 9953
rect 8385 9927 8391 9953
rect 11825 9927 11831 9953
rect 11857 9927 11863 9953
rect 14625 9927 14631 9953
rect 14657 9927 14663 9953
rect 8751 9921 8777 9927
rect 15471 9921 15497 9927
rect 8807 9897 8833 9903
rect 11713 9871 11719 9897
rect 11745 9871 11751 9897
rect 8807 9865 8833 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 6735 9729 6761 9735
rect 6735 9697 6761 9703
rect 6903 9729 6929 9735
rect 6903 9697 6929 9703
rect 9983 9729 10009 9735
rect 9983 9697 10009 9703
rect 10151 9729 10177 9735
rect 10151 9697 10177 9703
rect 7127 9673 7153 9679
rect 8751 9673 8777 9679
rect 7625 9647 7631 9673
rect 7657 9647 7663 9673
rect 8073 9647 8079 9673
rect 8105 9647 8111 9673
rect 9809 9647 9815 9673
rect 9841 9647 9847 9673
rect 16025 9647 16031 9673
rect 16057 9647 16063 9673
rect 7127 9641 7153 9647
rect 8751 9641 8777 9647
rect 8639 9617 8665 9623
rect 7569 9591 7575 9617
rect 7601 9591 7607 9617
rect 8297 9591 8303 9617
rect 8329 9591 8335 9617
rect 8639 9585 8665 9591
rect 9143 9617 9169 9623
rect 9143 9585 9169 9591
rect 9647 9617 9673 9623
rect 11047 9617 11073 9623
rect 12559 9617 12585 9623
rect 13399 9617 13425 9623
rect 10649 9591 10655 9617
rect 10681 9591 10687 9617
rect 11825 9591 11831 9617
rect 11857 9591 11863 9617
rect 12273 9591 12279 9617
rect 12305 9591 12311 9617
rect 12777 9591 12783 9617
rect 12809 9591 12815 9617
rect 13113 9591 13119 9617
rect 13145 9591 13151 9617
rect 13281 9591 13287 9617
rect 13313 9591 13319 9617
rect 14625 9591 14631 9617
rect 14657 9591 14663 9617
rect 9647 9585 9673 9591
rect 11047 9585 11073 9591
rect 12559 9585 12585 9591
rect 13399 9585 13425 9591
rect 6791 9561 6817 9567
rect 6791 9529 6817 9535
rect 7743 9561 7769 9567
rect 7743 9529 7769 9535
rect 8023 9561 8049 9567
rect 8023 9529 8049 9535
rect 8079 9561 8105 9567
rect 10207 9561 10233 9567
rect 9473 9535 9479 9561
rect 9505 9535 9511 9561
rect 8079 9529 8105 9535
rect 10207 9529 10233 9535
rect 10823 9561 10849 9567
rect 10823 9529 10849 9535
rect 11271 9561 11297 9567
rect 11271 9529 11297 9535
rect 12615 9561 12641 9567
rect 12615 9529 12641 9535
rect 12895 9561 12921 9567
rect 12895 9529 12921 9535
rect 13455 9561 13481 9567
rect 13959 9561 13985 9567
rect 13673 9535 13679 9561
rect 13705 9535 13711 9561
rect 13455 9529 13481 9535
rect 13959 9529 13985 9535
rect 14127 9561 14153 9567
rect 14961 9535 14967 9561
rect 14993 9535 14999 9561
rect 14127 9529 14153 9535
rect 7911 9505 7937 9511
rect 9871 9505 9897 9511
rect 8465 9479 8471 9505
rect 8497 9479 8503 9505
rect 9305 9479 9311 9505
rect 9337 9479 9343 9505
rect 7911 9473 7937 9479
rect 9871 9473 9897 9479
rect 10767 9505 10793 9511
rect 10767 9473 10793 9479
rect 11103 9505 11129 9511
rect 11103 9473 11129 9479
rect 11159 9505 11185 9511
rect 12951 9505 12977 9511
rect 11937 9479 11943 9505
rect 11969 9479 11975 9505
rect 11159 9473 11185 9479
rect 12951 9473 12977 9479
rect 13007 9505 13033 9511
rect 13007 9473 13033 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 7295 9337 7321 9343
rect 9703 9337 9729 9343
rect 7681 9311 7687 9337
rect 7713 9311 7719 9337
rect 12665 9311 12671 9337
rect 12697 9311 12703 9337
rect 7295 9305 7321 9311
rect 9703 9305 9729 9311
rect 9591 9281 9617 9287
rect 9591 9249 9617 9255
rect 10879 9281 10905 9287
rect 10879 9249 10905 9255
rect 10991 9281 11017 9287
rect 10991 9249 11017 9255
rect 11047 9281 11073 9287
rect 11047 9249 11073 9255
rect 11831 9281 11857 9287
rect 11831 9249 11857 9255
rect 11887 9281 11913 9287
rect 13735 9281 13761 9287
rect 13057 9255 13063 9281
rect 13089 9255 13095 9281
rect 11887 9249 11913 9255
rect 13735 9249 13761 9255
rect 13791 9281 13817 9287
rect 13791 9249 13817 9255
rect 7183 9225 7209 9231
rect 7183 9193 7209 9199
rect 7407 9225 7433 9231
rect 7407 9193 7433 9199
rect 7855 9225 7881 9231
rect 7855 9193 7881 9199
rect 10095 9225 10121 9231
rect 10095 9193 10121 9199
rect 10375 9225 10401 9231
rect 13567 9225 13593 9231
rect 12609 9199 12615 9225
rect 12641 9199 12647 9225
rect 13169 9199 13175 9225
rect 13201 9199 13207 9225
rect 13449 9199 13455 9225
rect 13481 9199 13487 9225
rect 13673 9199 13679 9225
rect 13705 9199 13711 9225
rect 14009 9199 14015 9225
rect 14041 9199 14047 9225
rect 14345 9199 14351 9225
rect 14377 9199 14383 9225
rect 18825 9199 18831 9225
rect 18857 9199 18863 9225
rect 10375 9193 10401 9199
rect 13567 9193 13593 9199
rect 7351 9169 7377 9175
rect 7351 9137 7377 9143
rect 9647 9169 9673 9175
rect 15639 9169 15665 9175
rect 15409 9143 15415 9169
rect 15441 9143 15447 9169
rect 9647 9137 9673 9143
rect 15639 9137 15665 9143
rect 7071 9113 7097 9119
rect 7071 9081 7097 9087
rect 11831 9113 11857 9119
rect 11831 9081 11857 9087
rect 20007 9113 20033 9119
rect 20007 9081 20033 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 8023 8945 8049 8951
rect 8023 8913 8049 8919
rect 14855 8945 14881 8951
rect 14855 8913 14881 8919
rect 967 8889 993 8895
rect 8359 8889 8385 8895
rect 12503 8889 12529 8895
rect 8185 8863 8191 8889
rect 8217 8863 8223 8889
rect 10873 8863 10879 8889
rect 10905 8863 10911 8889
rect 967 8857 993 8863
rect 8359 8857 8385 8863
rect 12503 8857 12529 8863
rect 14911 8889 14937 8895
rect 14911 8857 14937 8863
rect 20007 8889 20033 8895
rect 20007 8857 20033 8863
rect 10823 8833 10849 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 8521 8807 8527 8833
rect 8553 8807 8559 8833
rect 10823 8801 10849 8807
rect 11271 8833 11297 8839
rect 11271 8801 11297 8807
rect 11943 8833 11969 8839
rect 11943 8801 11969 8807
rect 12223 8833 12249 8839
rect 12223 8801 12249 8807
rect 12951 8833 12977 8839
rect 12951 8801 12977 8807
rect 13007 8833 13033 8839
rect 13007 8801 13033 8807
rect 13063 8833 13089 8839
rect 13063 8801 13089 8807
rect 13287 8833 13313 8839
rect 13505 8807 13511 8833
rect 13537 8807 13543 8833
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 13287 8801 13313 8807
rect 8135 8777 8161 8783
rect 8135 8745 8161 8751
rect 11327 8777 11353 8783
rect 11327 8745 11353 8751
rect 11439 8777 11465 8783
rect 11439 8745 11465 8751
rect 12055 8777 12081 8783
rect 13393 8751 13399 8777
rect 13425 8751 13431 8777
rect 12055 8745 12081 8751
rect 8415 8721 8441 8727
rect 8415 8689 8441 8695
rect 10991 8721 11017 8727
rect 10991 8689 11017 8695
rect 12167 8721 12193 8727
rect 12167 8689 12193 8695
rect 12783 8721 12809 8727
rect 12783 8689 12809 8695
rect 14631 8721 14657 8727
rect 14631 8689 14657 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 7351 8553 7377 8559
rect 11153 8527 11159 8553
rect 11185 8527 11191 8553
rect 12161 8527 12167 8553
rect 12193 8527 12199 8553
rect 7351 8521 7377 8527
rect 9591 8497 9617 8503
rect 6729 8471 6735 8497
rect 6761 8471 6767 8497
rect 9591 8465 9617 8471
rect 9647 8497 9673 8503
rect 9647 8465 9673 8471
rect 12335 8497 12361 8503
rect 13001 8471 13007 8497
rect 13033 8471 13039 8497
rect 12335 8465 12361 8471
rect 9535 8441 9561 8447
rect 7121 8415 7127 8441
rect 7153 8415 7159 8441
rect 9305 8415 9311 8441
rect 9337 8415 9343 8441
rect 9535 8409 9561 8415
rect 10543 8441 10569 8447
rect 10543 8409 10569 8415
rect 10599 8441 10625 8447
rect 10599 8409 10625 8415
rect 10711 8441 10737 8447
rect 10711 8409 10737 8415
rect 10767 8441 10793 8447
rect 10767 8409 10793 8415
rect 10991 8441 11017 8447
rect 14295 8441 14321 8447
rect 12665 8415 12671 8441
rect 12697 8415 12703 8441
rect 10991 8409 11017 8415
rect 14295 8409 14321 8415
rect 10655 8385 10681 8391
rect 5665 8359 5671 8385
rect 5697 8359 5703 8385
rect 14065 8359 14071 8385
rect 14097 8359 14103 8385
rect 10655 8353 10681 8359
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 6791 8161 6817 8167
rect 6791 8129 6817 8135
rect 10319 8161 10345 8167
rect 10319 8129 10345 8135
rect 10823 8161 10849 8167
rect 10823 8129 10849 8135
rect 6735 8105 6761 8111
rect 9255 8105 9281 8111
rect 7961 8079 7967 8105
rect 7993 8079 7999 8105
rect 9025 8079 9031 8105
rect 9057 8079 9063 8105
rect 6735 8073 6761 8079
rect 9255 8073 9281 8079
rect 11943 8105 11969 8111
rect 12161 8079 12167 8105
rect 12193 8079 12199 8105
rect 11943 8073 11969 8079
rect 9927 8049 9953 8055
rect 7625 8023 7631 8049
rect 7657 8023 7663 8049
rect 9927 8017 9953 8023
rect 10095 8049 10121 8055
rect 10095 8017 10121 8023
rect 10375 8049 10401 8055
rect 11047 8049 11073 8055
rect 10649 8023 10655 8049
rect 10681 8023 10687 8049
rect 10929 8023 10935 8049
rect 10961 8023 10967 8049
rect 12217 8023 12223 8049
rect 12249 8023 12255 8049
rect 12889 8023 12895 8049
rect 12921 8023 12927 8049
rect 13113 8023 13119 8049
rect 13145 8023 13151 8049
rect 10375 8017 10401 8023
rect 11047 8017 11073 8023
rect 13505 7967 13511 7993
rect 13537 7967 13543 7993
rect 10039 7937 10065 7943
rect 10039 7905 10065 7911
rect 10319 7937 10345 7943
rect 10319 7905 10345 7911
rect 10655 7937 10681 7943
rect 10655 7905 10681 7911
rect 12839 7937 12865 7943
rect 12839 7905 12865 7911
rect 13343 7937 13369 7943
rect 13343 7905 13369 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 11551 7769 11577 7775
rect 11551 7737 11577 7743
rect 12671 7769 12697 7775
rect 12889 7743 12895 7769
rect 12921 7743 12927 7769
rect 12671 7737 12697 7743
rect 8695 7713 8721 7719
rect 8695 7681 8721 7687
rect 8863 7713 8889 7719
rect 11103 7713 11129 7719
rect 9697 7687 9703 7713
rect 9729 7687 9735 7713
rect 8863 7681 8889 7687
rect 11103 7681 11129 7687
rect 11383 7713 11409 7719
rect 11383 7681 11409 7687
rect 11439 7713 11465 7719
rect 11439 7681 11465 7687
rect 12615 7713 12641 7719
rect 12615 7681 12641 7687
rect 10879 7657 10905 7663
rect 9305 7631 9311 7657
rect 9337 7631 9343 7657
rect 10879 7625 10905 7631
rect 11159 7657 11185 7663
rect 11159 7625 11185 7631
rect 10991 7601 11017 7607
rect 10761 7575 10767 7601
rect 10793 7575 10799 7601
rect 10991 7569 11017 7575
rect 13175 7601 13201 7607
rect 13175 7569 13201 7575
rect 13063 7545 13089 7551
rect 13063 7513 13089 7519
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 8353 7295 8359 7321
rect 8385 7295 8391 7321
rect 9417 7295 9423 7321
rect 9449 7295 9455 7321
rect 10655 7265 10681 7271
rect 8017 7239 8023 7265
rect 8049 7239 8055 7265
rect 10655 7233 10681 7239
rect 10823 7265 10849 7271
rect 13343 7265 13369 7271
rect 13225 7239 13231 7265
rect 13257 7239 13263 7265
rect 10823 7233 10849 7239
rect 13343 7233 13369 7239
rect 12559 7209 12585 7215
rect 12559 7177 12585 7183
rect 12727 7209 12753 7215
rect 12727 7177 12753 7183
rect 12895 7209 12921 7215
rect 13561 7183 13567 7209
rect 13593 7183 13599 7209
rect 12895 7177 12921 7183
rect 9647 7153 9673 7159
rect 9647 7121 9673 7127
rect 10711 7153 10737 7159
rect 10711 7121 10737 7127
rect 10991 7153 11017 7159
rect 10991 7121 11017 7127
rect 13735 7153 13761 7159
rect 13735 7121 13761 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 9199 6985 9225 6991
rect 9199 6953 9225 6959
rect 11831 6985 11857 6991
rect 11831 6953 11857 6959
rect 10201 6903 10207 6929
rect 10233 6903 10239 6929
rect 11601 6903 11607 6929
rect 11633 6903 11639 6929
rect 13001 6903 13007 6929
rect 13033 6903 13039 6929
rect 11439 6873 11465 6879
rect 9809 6847 9815 6873
rect 9841 6847 9847 6873
rect 12609 6847 12615 6873
rect 12641 6847 12647 6873
rect 11439 6841 11465 6847
rect 9143 6817 9169 6823
rect 14295 6817 14321 6823
rect 11265 6791 11271 6817
rect 11297 6791 11303 6817
rect 14065 6791 14071 6817
rect 14097 6791 14103 6817
rect 9143 6785 9169 6791
rect 14295 6785 14321 6791
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 13735 6537 13761 6543
rect 12385 6511 12391 6537
rect 12417 6511 12423 6537
rect 13449 6511 13455 6537
rect 13481 6511 13487 6537
rect 13735 6505 13761 6511
rect 12049 6455 12055 6481
rect 12081 6455 12087 6481
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 11159 2617 11185 2623
rect 11159 2585 11185 2591
rect 10649 2535 10655 2561
rect 10681 2535 10687 2561
rect 855 2449 881 2455
rect 855 2417 881 2423
rect 20119 2449 20145 2455
rect 20119 2417 20145 2423
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 9417 2143 9423 2169
rect 9449 2143 9455 2169
rect 11097 2143 11103 2169
rect 11129 2143 11135 2169
rect 9927 2057 9953 2063
rect 9927 2025 9953 2031
rect 11383 2057 11409 2063
rect 11383 2025 11409 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 11769 1751 11775 1777
rect 11801 1751 11807 1777
rect 11097 1695 11103 1721
rect 11129 1695 11135 1721
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9311 19111 9337 19137
rect 12783 19111 12809 19137
rect 11103 19055 11129 19081
rect 9031 18999 9057 19025
rect 11775 18999 11801 19025
rect 12279 18999 12305 19025
rect 10599 18887 10625 18913
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 9927 18719 9953 18745
rect 11383 18719 11409 18745
rect 20119 18663 20145 18689
rect 9423 18607 9449 18633
rect 10991 18607 11017 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9031 18327 9057 18353
rect 8527 18215 8553 18241
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 7911 14015 7937 14041
rect 8359 14015 8385 14041
rect 10151 14015 10177 14041
rect 7967 13903 7993 13929
rect 8135 13903 8161 13929
rect 8247 13903 8273 13929
rect 10263 13903 10289 13929
rect 8191 13847 8217 13873
rect 10655 13847 10681 13873
rect 11719 13847 11745 13873
rect 7911 13791 7937 13817
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 11047 13623 11073 13649
rect 9087 13567 9113 13593
rect 13679 13567 13705 13593
rect 20007 13567 20033 13593
rect 7631 13511 7657 13537
rect 11103 13511 11129 13537
rect 12279 13511 12305 13537
rect 18831 13511 18857 13537
rect 8023 13455 8049 13481
rect 12615 13455 12641 13481
rect 9311 13399 9337 13425
rect 13903 13399 13929 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 8919 13231 8945 13257
rect 9143 13231 9169 13257
rect 11383 13231 11409 13257
rect 11439 13231 11465 13257
rect 13231 13231 13257 13257
rect 7351 13175 7377 13201
rect 11495 13175 11521 13201
rect 2143 13119 2169 13145
rect 7015 13119 7041 13145
rect 8695 13119 8721 13145
rect 8807 13119 8833 13145
rect 9647 13119 9673 13145
rect 11327 13119 11353 13145
rect 11719 13119 11745 13145
rect 13119 13119 13145 13145
rect 13287 13119 13313 13145
rect 13903 13119 13929 13145
rect 18831 13119 18857 13145
rect 8415 13063 8441 13089
rect 9983 13063 10009 13089
rect 11047 13063 11073 13089
rect 14295 13063 14321 13089
rect 15359 13063 15385 13089
rect 15583 13063 15609 13089
rect 19951 13063 19977 13089
rect 967 13007 993 13033
rect 8751 13007 8777 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 10655 12839 10681 12865
rect 14127 12839 14153 12865
rect 7687 12783 7713 12809
rect 11159 12783 11185 12809
rect 12783 12783 12809 12809
rect 20007 12783 20033 12809
rect 7799 12727 7825 12753
rect 8415 12727 8441 12753
rect 8583 12727 8609 12753
rect 13119 12727 13145 12753
rect 14239 12727 14265 12753
rect 14743 12727 14769 12753
rect 18831 12727 18857 12753
rect 10711 12671 10737 12697
rect 12839 12671 12865 12697
rect 12951 12671 12977 12697
rect 14575 12671 14601 12697
rect 14631 12671 14657 12697
rect 7519 12615 7545 12641
rect 7631 12615 7657 12641
rect 8527 12615 8553 12641
rect 13063 12615 13089 12641
rect 13959 12615 13985 12641
rect 14071 12615 14097 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 8695 12447 8721 12473
rect 8975 12447 9001 12473
rect 10767 12447 10793 12473
rect 11327 12447 11353 12473
rect 9087 12391 9113 12417
rect 11047 12391 11073 12417
rect 11159 12391 11185 12417
rect 7575 12335 7601 12361
rect 8863 12335 8889 12361
rect 9143 12335 9169 12361
rect 10711 12335 10737 12361
rect 11439 12335 11465 12361
rect 12671 12335 12697 12361
rect 14295 12335 14321 12361
rect 6119 12279 6145 12305
rect 7183 12279 7209 12305
rect 7799 12279 7825 12305
rect 10823 12279 10849 12305
rect 13007 12279 13033 12305
rect 14071 12279 14097 12305
rect 14631 12279 14657 12305
rect 15695 12279 15721 12305
rect 15919 12279 15945 12305
rect 10935 12223 10961 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 7631 12055 7657 12081
rect 10991 12055 11017 12081
rect 13343 12055 13369 12081
rect 14183 12055 14209 12081
rect 7351 11999 7377 12025
rect 13007 11999 13033 12025
rect 13847 11999 13873 12025
rect 20007 11999 20033 12025
rect 6735 11943 6761 11969
rect 7239 11943 7265 11969
rect 7575 11943 7601 11969
rect 10823 11943 10849 11969
rect 11271 11943 11297 11969
rect 11607 11943 11633 11969
rect 12279 11943 12305 11969
rect 12839 11943 12865 11969
rect 14295 11943 14321 11969
rect 14575 11943 14601 11969
rect 14743 11943 14769 11969
rect 18831 11943 18857 11969
rect 6903 11887 6929 11913
rect 9199 11887 9225 11913
rect 10711 11887 10737 11913
rect 11159 11887 11185 11913
rect 12447 11887 12473 11913
rect 13119 11887 13145 11913
rect 13287 11887 13313 11913
rect 14015 11887 14041 11913
rect 14631 11887 14657 11913
rect 6847 11831 6873 11857
rect 7183 11831 7209 11857
rect 9031 11831 9057 11857
rect 11495 11831 11521 11857
rect 12391 11831 12417 11857
rect 13007 11831 13033 11857
rect 13343 11831 13369 11857
rect 14127 11831 14153 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 9255 11663 9281 11689
rect 12055 11663 12081 11689
rect 12839 11663 12865 11689
rect 8863 11607 8889 11633
rect 12895 11607 12921 11633
rect 2143 11551 2169 11577
rect 7295 11551 7321 11577
rect 7463 11551 7489 11577
rect 7575 11551 7601 11577
rect 7687 11551 7713 11577
rect 7799 11551 7825 11577
rect 8639 11551 8665 11577
rect 8919 11551 8945 11577
rect 9143 11551 9169 11577
rect 9199 11551 9225 11577
rect 9479 11551 9505 11577
rect 11327 11551 11353 11577
rect 11495 11551 11521 11577
rect 11607 11551 11633 11577
rect 11719 11551 11745 11577
rect 11775 11551 11801 11577
rect 12783 11551 12809 11577
rect 13007 11551 13033 11577
rect 13175 11551 13201 11577
rect 5839 11495 5865 11521
rect 6903 11495 6929 11521
rect 7631 11495 7657 11521
rect 8023 11495 8049 11521
rect 8751 11495 8777 11521
rect 9871 11495 9897 11521
rect 10935 11495 10961 11521
rect 11663 11495 11689 11521
rect 967 11439 993 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 6903 11271 6929 11297
rect 13119 11271 13145 11297
rect 967 11215 993 11241
rect 6791 11215 6817 11241
rect 7519 11215 7545 11241
rect 8471 11215 8497 11241
rect 9535 11215 9561 11241
rect 9759 11215 9785 11241
rect 10935 11215 10961 11241
rect 13623 11215 13649 11241
rect 20007 11215 20033 11241
rect 2143 11159 2169 11185
rect 7407 11159 7433 11185
rect 7575 11159 7601 11185
rect 7687 11159 7713 11185
rect 8079 11159 8105 11185
rect 10879 11159 10905 11185
rect 11159 11159 11185 11185
rect 11551 11159 11577 11185
rect 11719 11159 11745 11185
rect 13063 11159 13089 11185
rect 13847 11159 13873 11185
rect 18831 11159 18857 11185
rect 10095 11103 10121 11129
rect 11047 11103 11073 11129
rect 13567 11103 13593 11129
rect 6791 11047 6817 11073
rect 7463 11047 7489 11073
rect 10263 11047 10289 11073
rect 11439 11047 11465 11073
rect 11607 11047 11633 11073
rect 11999 11047 12025 11073
rect 12167 11047 12193 11073
rect 12671 11047 12697 11073
rect 12839 11047 12865 11073
rect 13119 11047 13145 11073
rect 13679 11047 13705 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 7799 10879 7825 10905
rect 11719 10879 11745 10905
rect 13455 10879 13481 10905
rect 6847 10823 6873 10849
rect 7631 10823 7657 10849
rect 9759 10823 9785 10849
rect 12895 10823 12921 10849
rect 12951 10823 12977 10849
rect 13511 10823 13537 10849
rect 14407 10823 14433 10849
rect 7239 10767 7265 10793
rect 7463 10767 7489 10793
rect 11495 10767 11521 10793
rect 11663 10767 11689 10793
rect 11831 10767 11857 10793
rect 11943 10767 11969 10793
rect 12783 10767 12809 10793
rect 13119 10767 13145 10793
rect 13343 10767 13369 10793
rect 13679 10767 13705 10793
rect 14015 10767 14041 10793
rect 5783 10711 5809 10737
rect 13175 10711 13201 10737
rect 13735 10711 13761 10737
rect 15471 10711 15497 10737
rect 15695 10711 15721 10737
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 967 10431 993 10457
rect 20007 10431 20033 10457
rect 2143 10375 2169 10401
rect 7911 10375 7937 10401
rect 9759 10375 9785 10401
rect 10263 10375 10289 10401
rect 10655 10375 10681 10401
rect 13455 10375 13481 10401
rect 13847 10375 13873 10401
rect 18831 10375 18857 10401
rect 6735 10319 6761 10345
rect 7631 10319 7657 10345
rect 7743 10319 7769 10345
rect 8415 10319 8441 10345
rect 8807 10319 8833 10345
rect 9871 10319 9897 10345
rect 10039 10319 10065 10345
rect 10375 10319 10401 10345
rect 12559 10319 12585 10345
rect 13567 10319 13593 10345
rect 13623 10319 13649 10345
rect 6791 10263 6817 10289
rect 6847 10263 6873 10289
rect 7799 10263 7825 10289
rect 8583 10263 8609 10289
rect 8975 10263 9001 10289
rect 13511 10263 13537 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 10823 10095 10849 10121
rect 11159 10095 11185 10121
rect 12223 10095 12249 10121
rect 6343 10039 6369 10065
rect 7295 10039 7321 10065
rect 9031 10039 9057 10065
rect 9479 10039 9505 10065
rect 10151 10039 10177 10065
rect 10207 10039 10233 10065
rect 12279 10039 12305 10065
rect 15415 10039 15441 10065
rect 6735 9983 6761 10009
rect 6959 9983 6985 10009
rect 9647 9983 9673 10009
rect 10095 9983 10121 10009
rect 10431 9983 10457 10009
rect 10655 9983 10681 10009
rect 10767 9983 10793 10009
rect 10991 9983 11017 10009
rect 11103 9983 11129 10009
rect 11271 9983 11297 10009
rect 11943 9983 11969 10009
rect 12615 9983 12641 10009
rect 5279 9927 5305 9953
rect 8359 9927 8385 9953
rect 8751 9927 8777 9953
rect 11831 9927 11857 9953
rect 14631 9927 14657 9953
rect 15471 9927 15497 9953
rect 8807 9871 8833 9897
rect 11719 9871 11745 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 6735 9703 6761 9729
rect 6903 9703 6929 9729
rect 9983 9703 10009 9729
rect 10151 9703 10177 9729
rect 7127 9647 7153 9673
rect 7631 9647 7657 9673
rect 8079 9647 8105 9673
rect 8751 9647 8777 9673
rect 9815 9647 9841 9673
rect 16031 9647 16057 9673
rect 7575 9591 7601 9617
rect 8303 9591 8329 9617
rect 8639 9591 8665 9617
rect 9143 9591 9169 9617
rect 9647 9591 9673 9617
rect 10655 9591 10681 9617
rect 11047 9591 11073 9617
rect 11831 9591 11857 9617
rect 12279 9591 12305 9617
rect 12559 9591 12585 9617
rect 12783 9591 12809 9617
rect 13119 9591 13145 9617
rect 13287 9591 13313 9617
rect 13399 9591 13425 9617
rect 14631 9591 14657 9617
rect 6791 9535 6817 9561
rect 7743 9535 7769 9561
rect 8023 9535 8049 9561
rect 8079 9535 8105 9561
rect 9479 9535 9505 9561
rect 10207 9535 10233 9561
rect 10823 9535 10849 9561
rect 11271 9535 11297 9561
rect 12615 9535 12641 9561
rect 12895 9535 12921 9561
rect 13455 9535 13481 9561
rect 13679 9535 13705 9561
rect 13959 9535 13985 9561
rect 14127 9535 14153 9561
rect 14967 9535 14993 9561
rect 7911 9479 7937 9505
rect 8471 9479 8497 9505
rect 9311 9479 9337 9505
rect 9871 9479 9897 9505
rect 10767 9479 10793 9505
rect 11103 9479 11129 9505
rect 11159 9479 11185 9505
rect 11943 9479 11969 9505
rect 12951 9479 12977 9505
rect 13007 9479 13033 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 7295 9311 7321 9337
rect 7687 9311 7713 9337
rect 9703 9311 9729 9337
rect 12671 9311 12697 9337
rect 9591 9255 9617 9281
rect 10879 9255 10905 9281
rect 10991 9255 11017 9281
rect 11047 9255 11073 9281
rect 11831 9255 11857 9281
rect 11887 9255 11913 9281
rect 13063 9255 13089 9281
rect 13735 9255 13761 9281
rect 13791 9255 13817 9281
rect 7183 9199 7209 9225
rect 7407 9199 7433 9225
rect 7855 9199 7881 9225
rect 10095 9199 10121 9225
rect 10375 9199 10401 9225
rect 12615 9199 12641 9225
rect 13175 9199 13201 9225
rect 13455 9199 13481 9225
rect 13567 9199 13593 9225
rect 13679 9199 13705 9225
rect 14015 9199 14041 9225
rect 14351 9199 14377 9225
rect 18831 9199 18857 9225
rect 7351 9143 7377 9169
rect 9647 9143 9673 9169
rect 15415 9143 15441 9169
rect 15639 9143 15665 9169
rect 7071 9087 7097 9113
rect 11831 9087 11857 9113
rect 20007 9087 20033 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 8023 8919 8049 8945
rect 14855 8919 14881 8945
rect 967 8863 993 8889
rect 8191 8863 8217 8889
rect 8359 8863 8385 8889
rect 10879 8863 10905 8889
rect 12503 8863 12529 8889
rect 14911 8863 14937 8889
rect 20007 8863 20033 8889
rect 2143 8807 2169 8833
rect 8527 8807 8553 8833
rect 10823 8807 10849 8833
rect 11271 8807 11297 8833
rect 11943 8807 11969 8833
rect 12223 8807 12249 8833
rect 12951 8807 12977 8833
rect 13007 8807 13033 8833
rect 13063 8807 13089 8833
rect 13287 8807 13313 8833
rect 13511 8807 13537 8833
rect 18831 8807 18857 8833
rect 8135 8751 8161 8777
rect 11327 8751 11353 8777
rect 11439 8751 11465 8777
rect 12055 8751 12081 8777
rect 13399 8751 13425 8777
rect 8415 8695 8441 8721
rect 10991 8695 11017 8721
rect 12167 8695 12193 8721
rect 12783 8695 12809 8721
rect 14631 8695 14657 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7351 8527 7377 8553
rect 11159 8527 11185 8553
rect 12167 8527 12193 8553
rect 6735 8471 6761 8497
rect 9591 8471 9617 8497
rect 9647 8471 9673 8497
rect 12335 8471 12361 8497
rect 13007 8471 13033 8497
rect 7127 8415 7153 8441
rect 9311 8415 9337 8441
rect 9535 8415 9561 8441
rect 10543 8415 10569 8441
rect 10599 8415 10625 8441
rect 10711 8415 10737 8441
rect 10767 8415 10793 8441
rect 10991 8415 11017 8441
rect 12671 8415 12697 8441
rect 14295 8415 14321 8441
rect 5671 8359 5697 8385
rect 10655 8359 10681 8385
rect 14071 8359 14097 8385
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 6791 8135 6817 8161
rect 10319 8135 10345 8161
rect 10823 8135 10849 8161
rect 6735 8079 6761 8105
rect 7967 8079 7993 8105
rect 9031 8079 9057 8105
rect 9255 8079 9281 8105
rect 11943 8079 11969 8105
rect 12167 8079 12193 8105
rect 7631 8023 7657 8049
rect 9927 8023 9953 8049
rect 10095 8023 10121 8049
rect 10375 8023 10401 8049
rect 10655 8023 10681 8049
rect 10935 8023 10961 8049
rect 11047 8023 11073 8049
rect 12223 8023 12249 8049
rect 12895 8023 12921 8049
rect 13119 8023 13145 8049
rect 13511 7967 13537 7993
rect 10039 7911 10065 7937
rect 10319 7911 10345 7937
rect 10655 7911 10681 7937
rect 12839 7911 12865 7937
rect 13343 7911 13369 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 11551 7743 11577 7769
rect 12671 7743 12697 7769
rect 12895 7743 12921 7769
rect 8695 7687 8721 7713
rect 8863 7687 8889 7713
rect 9703 7687 9729 7713
rect 11103 7687 11129 7713
rect 11383 7687 11409 7713
rect 11439 7687 11465 7713
rect 12615 7687 12641 7713
rect 9311 7631 9337 7657
rect 10879 7631 10905 7657
rect 11159 7631 11185 7657
rect 10767 7575 10793 7601
rect 10991 7575 11017 7601
rect 13175 7575 13201 7601
rect 13063 7519 13089 7545
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 8359 7295 8385 7321
rect 9423 7295 9449 7321
rect 8023 7239 8049 7265
rect 10655 7239 10681 7265
rect 10823 7239 10849 7265
rect 13231 7239 13257 7265
rect 13343 7239 13369 7265
rect 12559 7183 12585 7209
rect 12727 7183 12753 7209
rect 12895 7183 12921 7209
rect 13567 7183 13593 7209
rect 9647 7127 9673 7153
rect 10711 7127 10737 7153
rect 10991 7127 11017 7153
rect 13735 7127 13761 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 9199 6959 9225 6985
rect 11831 6959 11857 6985
rect 10207 6903 10233 6929
rect 11607 6903 11633 6929
rect 13007 6903 13033 6929
rect 9815 6847 9841 6873
rect 11439 6847 11465 6873
rect 12615 6847 12641 6873
rect 9143 6791 9169 6817
rect 11271 6791 11297 6817
rect 14071 6791 14097 6817
rect 14295 6791 14321 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 12391 6511 12417 6537
rect 13455 6511 13481 6537
rect 13735 6511 13761 6537
rect 12055 6455 12081 6481
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 11159 2591 11185 2617
rect 10655 2535 10681 2561
rect 855 2423 881 2449
rect 20119 2423 20145 2449
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 9423 2143 9449 2169
rect 11103 2143 11129 2169
rect 9927 2031 9953 2057
rect 11383 2031 11409 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 11775 1751 11801 1777
rect 11103 1695 11129 1721
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8400 20600 8456 21000
rect 9072 20600 9128 21000
rect 9408 20600 9464 21000
rect 10752 20600 10808 21000
rect 11088 20600 11144 21000
rect 11424 20600 11480 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 8414 18354 8442 20600
rect 9086 19138 9114 20600
rect 9310 19138 9338 19143
rect 9086 19137 9338 19138
rect 9086 19111 9311 19137
rect 9337 19111 9338 19137
rect 9086 19110 9338 19111
rect 9310 19105 9338 19110
rect 9030 19026 9058 19031
rect 9030 19025 9114 19026
rect 9030 18999 9031 19025
rect 9057 18999 9114 19025
rect 9030 18998 9114 18999
rect 9030 18993 9058 18998
rect 8414 18321 8442 18326
rect 9030 18354 9058 18359
rect 9030 18307 9058 18326
rect 8526 18241 8554 18247
rect 8526 18215 8527 18241
rect 8553 18215 8554 18241
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 8526 15974 8554 18215
rect 8414 15946 8554 15974
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 7910 14042 7938 14047
rect 8358 14042 8386 14047
rect 8414 14042 8442 15946
rect 7910 14041 8218 14042
rect 7910 14015 7911 14041
rect 7937 14015 8218 14041
rect 7910 14014 8218 14015
rect 7910 14009 7938 14014
rect 7966 13929 7994 13935
rect 7966 13903 7967 13929
rect 7993 13903 7994 13929
rect 7350 13818 7378 13823
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 2086 13482 2114 13487
rect 966 13033 994 13039
rect 966 13007 967 13033
rect 993 13007 994 13033
rect 966 12810 994 13007
rect 966 12777 994 12782
rect 966 11466 994 11471
rect 966 11419 994 11438
rect 966 11242 994 11247
rect 966 11195 994 11214
rect 966 10457 994 10463
rect 966 10431 967 10457
rect 993 10431 994 10457
rect 966 10122 994 10431
rect 2086 10402 2114 13454
rect 7350 13201 7378 13790
rect 7910 13818 7938 13823
rect 7910 13771 7938 13790
rect 7630 13537 7658 13543
rect 7630 13511 7631 13537
rect 7657 13511 7658 13537
rect 7630 13482 7658 13511
rect 7350 13175 7351 13201
rect 7377 13175 7378 13201
rect 7350 13169 7378 13175
rect 7518 13454 7658 13482
rect 2142 13146 2170 13151
rect 2142 13099 2170 13118
rect 6118 13146 6146 13151
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 6118 12698 6146 13118
rect 6118 12305 6146 12670
rect 7014 13145 7042 13151
rect 7014 13119 7015 13145
rect 7041 13119 7042 13145
rect 7014 12642 7042 13119
rect 7518 12754 7546 13454
rect 7798 13146 7826 13151
rect 7686 12809 7714 12815
rect 7686 12783 7687 12809
rect 7713 12783 7714 12809
rect 7518 12726 7602 12754
rect 7406 12698 7434 12703
rect 7406 12642 7434 12670
rect 7518 12642 7546 12647
rect 7406 12641 7546 12642
rect 7406 12615 7519 12641
rect 7545 12615 7546 12641
rect 7406 12614 7546 12615
rect 7014 12609 7042 12614
rect 7518 12609 7546 12614
rect 7574 12586 7602 12726
rect 7574 12361 7602 12558
rect 7574 12335 7575 12361
rect 7601 12335 7602 12361
rect 7574 12329 7602 12335
rect 7630 12641 7658 12647
rect 7630 12615 7631 12641
rect 7657 12615 7658 12641
rect 7630 12474 7658 12615
rect 6118 12279 6119 12305
rect 6145 12279 6146 12305
rect 6118 12273 6146 12279
rect 7182 12305 7210 12311
rect 7182 12279 7183 12305
rect 7209 12279 7210 12305
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 6734 11970 6762 11975
rect 2142 11578 2170 11583
rect 2142 11531 2170 11550
rect 5838 11578 5866 11583
rect 5838 11521 5866 11550
rect 5838 11495 5839 11521
rect 5865 11495 5866 11521
rect 5838 11489 5866 11495
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 2142 11186 2170 11191
rect 2142 11139 2170 11158
rect 5782 11186 5810 11191
rect 5782 11074 5810 11158
rect 6734 11074 6762 11942
rect 6902 11914 6930 11919
rect 6902 11867 6930 11886
rect 6846 11857 6874 11863
rect 6846 11831 6847 11857
rect 6873 11831 6874 11857
rect 6846 11634 6874 11831
rect 7182 11857 7210 12279
rect 7630 12250 7658 12446
rect 7574 12222 7658 12250
rect 7350 12026 7378 12031
rect 7294 12025 7378 12026
rect 7294 11999 7351 12025
rect 7377 11999 7378 12025
rect 7294 11998 7378 11999
rect 7182 11831 7183 11857
rect 7209 11831 7210 11857
rect 7182 11825 7210 11831
rect 7238 11969 7266 11975
rect 7238 11943 7239 11969
rect 7265 11943 7266 11969
rect 7238 11746 7266 11943
rect 7294 11970 7322 11998
rect 7350 11993 7378 11998
rect 7294 11937 7322 11942
rect 7574 11969 7602 12222
rect 7630 12082 7658 12087
rect 7686 12082 7714 12783
rect 7798 12753 7826 13118
rect 7798 12727 7799 12753
rect 7825 12727 7826 12753
rect 7798 12721 7826 12727
rect 7630 12081 7714 12082
rect 7630 12055 7631 12081
rect 7657 12055 7714 12081
rect 7630 12054 7714 12055
rect 7798 12642 7826 12647
rect 7798 12305 7826 12614
rect 7798 12279 7799 12305
rect 7825 12279 7826 12305
rect 7630 12049 7658 12054
rect 7798 12026 7826 12279
rect 7574 11943 7575 11969
rect 7601 11943 7602 11969
rect 7574 11937 7602 11943
rect 7742 11998 7826 12026
rect 7406 11914 7434 11919
rect 7434 11886 7546 11914
rect 7406 11881 7434 11886
rect 7238 11713 7266 11718
rect 7462 11690 7490 11695
rect 6846 11606 6986 11634
rect 6902 11522 6930 11527
rect 6790 11521 6930 11522
rect 6790 11495 6903 11521
rect 6929 11495 6930 11521
rect 6790 11494 6930 11495
rect 6790 11241 6818 11494
rect 6902 11489 6930 11494
rect 6902 11410 6930 11415
rect 6902 11297 6930 11382
rect 6902 11271 6903 11297
rect 6929 11271 6930 11297
rect 6902 11265 6930 11271
rect 6790 11215 6791 11241
rect 6817 11215 6818 11241
rect 6790 11209 6818 11215
rect 6790 11074 6818 11079
rect 6734 11073 6818 11074
rect 6734 11047 6791 11073
rect 6817 11047 6818 11073
rect 6734 11046 6818 11047
rect 5782 10737 5810 11046
rect 6790 10794 6818 11046
rect 6846 10850 6874 10855
rect 6958 10850 6986 11606
rect 6846 10849 6986 10850
rect 6846 10823 6847 10849
rect 6873 10823 6986 10849
rect 6846 10822 6986 10823
rect 7294 11578 7322 11583
rect 6846 10817 6874 10822
rect 7238 10794 7266 10799
rect 7294 10794 7322 11550
rect 7462 11577 7490 11662
rect 7462 11551 7463 11577
rect 7489 11551 7490 11577
rect 7406 11186 7434 11191
rect 7462 11186 7490 11551
rect 7518 11241 7546 11886
rect 7574 11577 7602 11583
rect 7574 11551 7575 11577
rect 7601 11551 7602 11577
rect 7574 11522 7602 11551
rect 7686 11577 7714 11583
rect 7686 11551 7687 11577
rect 7713 11551 7714 11577
rect 7574 11489 7602 11494
rect 7630 11521 7658 11527
rect 7630 11495 7631 11521
rect 7657 11495 7658 11521
rect 7630 11410 7658 11495
rect 7630 11377 7658 11382
rect 7686 11298 7714 11551
rect 7742 11578 7770 11998
rect 7910 11746 7938 11751
rect 7742 11545 7770 11550
rect 7798 11577 7826 11583
rect 7798 11551 7799 11577
rect 7825 11551 7826 11577
rect 7798 11522 7826 11551
rect 7798 11489 7826 11494
rect 7518 11215 7519 11241
rect 7545 11215 7546 11241
rect 7518 11209 7546 11215
rect 7574 11270 7714 11298
rect 7742 11354 7770 11359
rect 7406 11185 7490 11186
rect 7406 11159 7407 11185
rect 7433 11159 7490 11185
rect 7406 11158 7490 11159
rect 7574 11185 7602 11270
rect 7574 11159 7575 11185
rect 7601 11159 7602 11185
rect 7406 11153 7434 11158
rect 7462 11074 7490 11079
rect 7462 11027 7490 11046
rect 7462 10794 7490 10799
rect 6790 10761 6818 10766
rect 6958 10793 7490 10794
rect 6958 10767 7239 10793
rect 7265 10767 7463 10793
rect 7489 10767 7490 10793
rect 6958 10766 7490 10767
rect 5782 10711 5783 10737
rect 5809 10711 5810 10737
rect 5782 10705 5810 10711
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 2086 10369 2114 10374
rect 2142 10401 2170 10407
rect 2142 10375 2143 10401
rect 2169 10375 2170 10401
rect 966 10089 994 10094
rect 2142 9954 2170 10375
rect 6734 10345 6762 10351
rect 6734 10319 6735 10345
rect 6761 10319 6762 10345
rect 6342 10290 6370 10295
rect 6342 10065 6370 10262
rect 6734 10122 6762 10319
rect 6790 10290 6818 10295
rect 6790 10243 6818 10262
rect 6846 10289 6874 10295
rect 6846 10263 6847 10289
rect 6873 10263 6874 10289
rect 6846 10178 6874 10263
rect 6846 10145 6874 10150
rect 6342 10039 6343 10065
rect 6369 10039 6370 10065
rect 6342 10033 6370 10039
rect 6678 10094 6762 10122
rect 2142 9921 2170 9926
rect 5278 9954 5306 9959
rect 5278 9907 5306 9926
rect 6678 9898 6706 10094
rect 6958 10066 6986 10766
rect 6734 10038 6986 10066
rect 6734 10009 6762 10038
rect 6734 9983 6735 10009
rect 6761 9983 6762 10009
rect 6734 9977 6762 9983
rect 6958 10009 6986 10038
rect 6958 9983 6959 10009
rect 6985 9983 6986 10009
rect 6958 9977 6986 9983
rect 6790 9898 6818 9903
rect 6678 9870 6762 9898
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 6734 9729 6762 9870
rect 6734 9703 6735 9729
rect 6761 9703 6762 9729
rect 6734 9697 6762 9703
rect 6790 9561 6818 9870
rect 6902 9730 6930 9735
rect 6902 9683 6930 9702
rect 6790 9535 6791 9561
rect 6817 9535 6818 9561
rect 6790 9529 6818 9535
rect 7126 9673 7154 10766
rect 7238 10761 7266 10766
rect 7462 10761 7490 10766
rect 7294 10178 7322 10183
rect 7126 9647 7127 9673
rect 7153 9647 7154 9673
rect 6734 9170 6762 9175
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 966 8890 994 8895
rect 966 8843 994 8862
rect 2142 8834 2170 8839
rect 2142 8787 2170 8806
rect 5670 8834 5698 8839
rect 5670 8385 5698 8806
rect 6734 8497 6762 9142
rect 7070 9114 7098 9119
rect 6734 8471 6735 8497
rect 6761 8471 6762 8497
rect 6734 8465 6762 8471
rect 6790 9113 7098 9114
rect 6790 9087 7071 9113
rect 7097 9087 7098 9113
rect 6790 9086 7098 9087
rect 5670 8359 5671 8385
rect 5697 8359 5698 8385
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 5670 8106 5698 8359
rect 6790 8161 6818 9086
rect 7070 9081 7098 9086
rect 7126 8554 7154 9647
rect 7182 10066 7210 10071
rect 7182 9562 7210 10038
rect 7294 10065 7322 10150
rect 7294 10039 7295 10065
rect 7321 10039 7322 10065
rect 7294 10033 7322 10039
rect 7574 9618 7602 11159
rect 7686 11186 7714 11191
rect 7742 11186 7770 11326
rect 7686 11185 7770 11186
rect 7686 11159 7687 11185
rect 7713 11159 7770 11185
rect 7686 11158 7770 11159
rect 7686 11153 7714 11158
rect 7798 10906 7826 10911
rect 7798 10859 7826 10878
rect 7630 10849 7658 10855
rect 7630 10823 7631 10849
rect 7657 10823 7658 10849
rect 7630 10794 7658 10823
rect 7630 10761 7658 10766
rect 7910 10402 7938 11718
rect 7966 11074 7994 13903
rect 8134 13929 8162 13935
rect 8134 13903 8135 13929
rect 8161 13903 8162 13929
rect 8022 13481 8050 13487
rect 8022 13455 8023 13481
rect 8049 13455 8050 13481
rect 8022 12866 8050 13455
rect 8134 13146 8162 13903
rect 8190 13873 8218 14014
rect 8358 14041 8442 14042
rect 8358 14015 8359 14041
rect 8385 14015 8442 14041
rect 8358 14014 8442 14015
rect 8358 14009 8386 14014
rect 8190 13847 8191 13873
rect 8217 13847 8218 13873
rect 8190 13841 8218 13847
rect 8246 13929 8274 13935
rect 8246 13903 8247 13929
rect 8273 13903 8274 13929
rect 8134 13113 8162 13118
rect 8022 12833 8050 12838
rect 8246 12474 8274 13903
rect 8414 13089 8442 14014
rect 9086 13594 9114 18998
rect 9422 18746 9450 20600
rect 10598 18914 10626 18919
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 9422 18713 9450 18718
rect 9926 18746 9954 18751
rect 9926 18699 9954 18718
rect 9422 18633 9450 18639
rect 9422 18607 9423 18633
rect 9449 18607 9450 18633
rect 9422 15974 9450 18607
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 8918 13593 9114 13594
rect 8918 13567 9087 13593
rect 9113 13567 9114 13593
rect 8918 13566 9114 13567
rect 8918 13257 8946 13566
rect 9086 13561 9114 13566
rect 9254 15946 9450 15974
rect 8918 13231 8919 13257
rect 8945 13231 8946 13257
rect 8918 13225 8946 13231
rect 9142 13426 9170 13431
rect 9142 13257 9170 13398
rect 9142 13231 9143 13257
rect 9169 13231 9170 13257
rect 9142 13225 9170 13231
rect 8694 13146 8722 13151
rect 8694 13099 8722 13118
rect 8806 13145 8834 13151
rect 8806 13119 8807 13145
rect 8833 13119 8834 13145
rect 8414 13063 8415 13089
rect 8441 13063 8442 13089
rect 8414 13057 8442 13063
rect 8750 13034 8778 13039
rect 8582 13033 8778 13034
rect 8582 13007 8751 13033
rect 8777 13007 8778 13033
rect 8582 13006 8778 13007
rect 8414 12866 8442 12871
rect 8414 12753 8442 12838
rect 8414 12727 8415 12753
rect 8441 12727 8442 12753
rect 8414 12721 8442 12727
rect 8582 12753 8610 13006
rect 8750 13001 8778 13006
rect 8806 12810 8834 13119
rect 8582 12727 8583 12753
rect 8609 12727 8610 12753
rect 8582 12721 8610 12727
rect 8750 12782 8834 12810
rect 8526 12642 8554 12647
rect 8526 12641 8666 12642
rect 8526 12615 8527 12641
rect 8553 12615 8666 12641
rect 8526 12614 8666 12615
rect 8526 12609 8554 12614
rect 8246 12441 8274 12446
rect 8638 12362 8666 12614
rect 8694 12474 8722 12479
rect 8750 12474 8778 12782
rect 8974 12474 9002 12479
rect 8722 12446 8778 12474
rect 8806 12473 9002 12474
rect 8806 12447 8975 12473
rect 9001 12447 9002 12473
rect 8806 12446 9002 12447
rect 8694 12427 8722 12446
rect 8806 12362 8834 12446
rect 8974 12441 9002 12446
rect 9086 12417 9114 12423
rect 9086 12391 9087 12417
rect 9113 12391 9114 12417
rect 8638 12334 8834 12362
rect 8862 12361 8890 12367
rect 8862 12335 8863 12361
rect 8889 12335 8890 12361
rect 8862 11914 8890 12335
rect 8862 11881 8890 11886
rect 9030 11857 9058 11863
rect 9030 11831 9031 11857
rect 9057 11831 9058 11857
rect 9030 11802 9058 11831
rect 8806 11774 9058 11802
rect 9086 11858 9114 12391
rect 8806 11634 8834 11774
rect 9086 11746 9114 11830
rect 8806 11601 8834 11606
rect 8862 11718 9114 11746
rect 9142 12361 9170 12367
rect 9142 12335 9143 12361
rect 9169 12335 9170 12361
rect 8862 11633 8890 11718
rect 9142 11690 9170 12335
rect 9198 11914 9226 11919
rect 9198 11867 9226 11886
rect 8862 11607 8863 11633
rect 8889 11607 8890 11633
rect 8862 11601 8890 11607
rect 9086 11662 9170 11690
rect 9254 11690 9282 15946
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9646 14042 9674 14047
rect 9310 13426 9338 13431
rect 9310 13379 9338 13398
rect 9646 13426 9674 14014
rect 10150 14042 10178 14047
rect 10178 14014 10290 14042
rect 10150 13995 10178 14014
rect 10262 13929 10290 14014
rect 10262 13903 10263 13929
rect 10289 13903 10290 13929
rect 10262 13897 10290 13903
rect 9646 13145 9674 13398
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9646 13119 9647 13145
rect 9673 13119 9674 13145
rect 9646 12810 9674 13119
rect 9982 13090 10010 13095
rect 9982 13043 10010 13062
rect 9674 12782 9786 12810
rect 9646 12777 9674 12782
rect 9254 11689 9562 11690
rect 9254 11663 9255 11689
rect 9281 11663 9562 11689
rect 9254 11662 9562 11663
rect 8022 11578 8050 11583
rect 8022 11521 8050 11550
rect 8022 11495 8023 11521
rect 8049 11495 8050 11521
rect 8022 11186 8050 11495
rect 8302 11578 8330 11583
rect 8078 11186 8106 11191
rect 8022 11185 8106 11186
rect 8022 11159 8079 11185
rect 8105 11159 8106 11185
rect 8022 11158 8106 11159
rect 8078 11153 8106 11158
rect 8302 11074 8330 11550
rect 8638 11578 8666 11583
rect 8638 11531 8666 11550
rect 8918 11578 8946 11583
rect 8918 11531 8946 11550
rect 8750 11521 8778 11527
rect 8750 11495 8751 11521
rect 8777 11495 8778 11521
rect 8750 11298 8778 11495
rect 8470 11270 8778 11298
rect 9086 11522 9114 11662
rect 9254 11657 9282 11662
rect 8470 11241 8498 11270
rect 8470 11215 8471 11241
rect 8497 11215 8498 11241
rect 8470 11209 8498 11215
rect 9086 11186 9114 11494
rect 9086 11153 9114 11158
rect 9142 11577 9170 11583
rect 9142 11551 9143 11577
rect 9169 11551 9170 11577
rect 7966 11046 8106 11074
rect 7910 10401 8050 10402
rect 7910 10375 7911 10401
rect 7937 10375 8050 10401
rect 7910 10374 8050 10375
rect 7910 10369 7938 10374
rect 7630 10345 7658 10351
rect 7630 10319 7631 10345
rect 7657 10319 7658 10345
rect 7630 9673 7658 10319
rect 7742 10346 7770 10351
rect 7742 10299 7770 10318
rect 7798 10290 7826 10295
rect 7798 10243 7826 10262
rect 7630 9647 7631 9673
rect 7657 9647 7658 9673
rect 7630 9641 7658 9647
rect 7574 9571 7602 9590
rect 7182 9225 7210 9534
rect 7742 9561 7770 9567
rect 7742 9535 7743 9561
rect 7769 9535 7770 9561
rect 7294 9338 7322 9343
rect 7294 9291 7322 9310
rect 7686 9338 7714 9343
rect 7686 9291 7714 9310
rect 7182 9199 7183 9225
rect 7209 9199 7210 9225
rect 7182 9193 7210 9199
rect 7406 9226 7434 9231
rect 7742 9226 7770 9535
rect 8022 9561 8050 10374
rect 8078 9673 8106 11046
rect 8078 9647 8079 9673
rect 8105 9647 8106 9673
rect 8078 9641 8106 9647
rect 8302 9617 8330 11046
rect 9142 10906 9170 11551
rect 9198 11578 9226 11583
rect 9198 11531 9226 11550
rect 9478 11578 9506 11583
rect 9478 11531 9506 11550
rect 9534 11241 9562 11662
rect 9534 11215 9535 11241
rect 9561 11215 9562 11241
rect 9534 11209 9562 11215
rect 9758 11241 9786 12782
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 10094 11858 10122 11863
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9870 11522 9898 11527
rect 9870 11475 9898 11494
rect 9758 11215 9759 11241
rect 9785 11215 9786 11241
rect 9170 10878 9226 10906
rect 9142 10873 9170 10878
rect 8414 10346 8442 10351
rect 8806 10346 8834 10351
rect 8414 10299 8442 10318
rect 8750 10345 8834 10346
rect 8750 10319 8807 10345
rect 8833 10319 8834 10345
rect 8750 10318 8834 10319
rect 8582 10289 8610 10295
rect 8582 10263 8583 10289
rect 8609 10263 8610 10289
rect 8358 9954 8386 9959
rect 8358 9907 8386 9926
rect 8582 9898 8610 10263
rect 8750 9954 8778 10318
rect 8806 10313 8834 10318
rect 8974 10290 9002 10295
rect 8974 10243 9002 10262
rect 9198 10178 9226 10878
rect 9758 10850 9786 11215
rect 10094 11129 10122 11830
rect 10598 11522 10626 18886
rect 10766 18746 10794 20600
rect 11102 19081 11130 20600
rect 11438 19138 11466 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 11438 19105 11466 19110
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 11102 19055 11103 19081
rect 11129 19055 11130 19081
rect 11102 19049 11130 19055
rect 11774 19025 11802 19031
rect 11774 18999 11775 19025
rect 11801 18999 11802 19025
rect 11774 18914 11802 18999
rect 11774 18881 11802 18886
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 10766 18713 10794 18718
rect 11382 18746 11410 18751
rect 11382 18699 11410 18718
rect 10990 18633 11018 18639
rect 10990 18607 10991 18633
rect 11017 18607 11018 18633
rect 10654 13874 10682 13879
rect 10654 13827 10682 13846
rect 10990 13454 11018 18607
rect 11046 13874 11074 13879
rect 11046 13649 11074 13846
rect 11046 13623 11047 13649
rect 11073 13623 11074 13649
rect 11046 13617 11074 13623
rect 11438 13874 11466 13879
rect 11102 13537 11130 13543
rect 11102 13511 11103 13537
rect 11129 13511 11130 13537
rect 11102 13454 11130 13511
rect 10990 13426 11074 13454
rect 11102 13426 11410 13454
rect 10654 13090 10682 13095
rect 10654 12865 10682 13062
rect 11046 13090 11074 13426
rect 11382 13257 11410 13426
rect 11382 13231 11383 13257
rect 11409 13231 11410 13257
rect 11382 13225 11410 13231
rect 11438 13257 11466 13846
rect 11718 13874 11746 13879
rect 11718 13827 11746 13846
rect 12278 13874 12306 18999
rect 20118 18689 20146 18695
rect 20118 18663 20119 18689
rect 20145 18663 20146 18689
rect 20118 18522 20146 18663
rect 20118 18489 20146 18494
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 12278 13841 12306 13846
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 13678 13594 13706 13599
rect 12278 13537 12306 13543
rect 12278 13511 12279 13537
rect 12305 13511 12306 13537
rect 12278 13482 12306 13511
rect 12278 13449 12306 13454
rect 12614 13482 12642 13487
rect 12614 13481 12810 13482
rect 12614 13455 12615 13481
rect 12641 13455 12810 13481
rect 12614 13454 12810 13455
rect 12614 13449 12642 13454
rect 11438 13231 11439 13257
rect 11465 13231 11466 13257
rect 11438 13225 11466 13231
rect 11494 13201 11522 13207
rect 11494 13175 11495 13201
rect 11521 13175 11522 13201
rect 11326 13145 11354 13151
rect 11326 13119 11327 13145
rect 11353 13119 11354 13145
rect 11046 13089 11130 13090
rect 11046 13063 11047 13089
rect 11073 13063 11130 13089
rect 11046 13062 11130 13063
rect 11046 13057 11074 13062
rect 10654 12839 10655 12865
rect 10681 12839 10682 12865
rect 10654 12833 10682 12839
rect 10710 12697 10738 12703
rect 10990 12698 11018 12703
rect 10710 12671 10711 12697
rect 10737 12671 10738 12697
rect 10710 12474 10738 12671
rect 10934 12670 10990 12698
rect 10766 12474 10794 12479
rect 10710 12473 10794 12474
rect 10710 12447 10767 12473
rect 10793 12447 10794 12473
rect 10710 12446 10794 12447
rect 10766 12441 10794 12446
rect 10710 12362 10738 12367
rect 10934 12362 10962 12670
rect 10990 12665 11018 12670
rect 10654 12361 10738 12362
rect 10654 12335 10711 12361
rect 10737 12335 10738 12361
rect 10654 12334 10738 12335
rect 10654 11858 10682 12334
rect 10710 12329 10738 12334
rect 10878 12334 10962 12362
rect 11046 12642 11074 12647
rect 11046 12417 11074 12614
rect 11046 12391 11047 12417
rect 11073 12391 11074 12417
rect 11046 12362 11074 12391
rect 11102 12418 11130 13062
rect 11158 12810 11186 12815
rect 11158 12763 11186 12782
rect 11158 12698 11186 12703
rect 11186 12670 11242 12698
rect 11158 12665 11186 12670
rect 11158 12418 11186 12423
rect 11102 12417 11186 12418
rect 11102 12391 11159 12417
rect 11185 12391 11186 12417
rect 11102 12390 11186 12391
rect 11158 12385 11186 12390
rect 11046 12334 11130 12362
rect 10822 12306 10850 12311
rect 10766 12305 10850 12306
rect 10766 12279 10823 12305
rect 10849 12279 10850 12305
rect 10766 12278 10850 12279
rect 10654 11825 10682 11830
rect 10710 11914 10738 11919
rect 10542 11354 10570 11359
rect 10094 11103 10095 11129
rect 10121 11103 10122 11129
rect 10094 11097 10122 11103
rect 10374 11298 10402 11303
rect 10206 11074 10234 11079
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 9702 10849 9786 10850
rect 9702 10823 9759 10849
rect 9785 10823 9786 10849
rect 9702 10822 9786 10823
rect 9198 10150 9338 10178
rect 9030 10066 9058 10071
rect 9030 10019 9058 10038
rect 9254 10066 9282 10071
rect 9310 10066 9338 10150
rect 9478 10066 9506 10071
rect 9310 10065 9506 10066
rect 9310 10039 9479 10065
rect 9505 10039 9506 10065
rect 9310 10038 9506 10039
rect 8750 9907 8778 9926
rect 9142 9954 9170 9959
rect 8582 9865 8610 9870
rect 8806 9898 8834 9903
rect 8302 9591 8303 9617
rect 8329 9591 8330 9617
rect 8302 9585 8330 9591
rect 8638 9730 8666 9735
rect 8638 9617 8666 9702
rect 8750 9674 8778 9679
rect 8806 9674 8834 9870
rect 8750 9673 8834 9674
rect 8750 9647 8751 9673
rect 8777 9647 8834 9673
rect 8750 9646 8834 9647
rect 8750 9641 8778 9646
rect 8638 9591 8639 9617
rect 8665 9591 8666 9617
rect 8022 9535 8023 9561
rect 8049 9535 8050 9561
rect 7910 9506 7938 9511
rect 7910 9505 7994 9506
rect 7910 9479 7911 9505
rect 7937 9479 7994 9505
rect 7910 9478 7994 9479
rect 7910 9473 7938 9478
rect 7854 9226 7882 9231
rect 7742 9225 7882 9226
rect 7742 9199 7855 9225
rect 7881 9199 7882 9225
rect 7742 9198 7882 9199
rect 7406 9179 7434 9198
rect 7350 9170 7378 9175
rect 7350 9123 7378 9142
rect 7854 9114 7882 9198
rect 7854 9081 7882 9086
rect 7966 8946 7994 9478
rect 8022 9338 8050 9535
rect 8078 9562 8106 9567
rect 8078 9515 8106 9534
rect 8470 9562 8498 9567
rect 8470 9505 8498 9534
rect 8470 9479 8471 9505
rect 8497 9479 8498 9505
rect 8470 9473 8498 9479
rect 8022 9305 8050 9310
rect 8190 9114 8218 9119
rect 8134 9086 8190 9114
rect 8022 8946 8050 8951
rect 7966 8918 8022 8946
rect 8022 8899 8050 8918
rect 8134 8777 8162 9086
rect 8190 9081 8218 9086
rect 8190 8890 8218 8895
rect 8358 8890 8386 8895
rect 8190 8889 8386 8890
rect 8190 8863 8191 8889
rect 8217 8863 8359 8889
rect 8385 8863 8386 8889
rect 8190 8862 8386 8863
rect 8190 8857 8218 8862
rect 8358 8857 8386 8862
rect 8526 8834 8554 8839
rect 8638 8834 8666 9591
rect 9142 9617 9170 9926
rect 9142 9591 9143 9617
rect 9169 9591 9170 9617
rect 9142 9585 9170 9591
rect 8526 8833 8666 8834
rect 8526 8807 8527 8833
rect 8553 8807 8666 8833
rect 8526 8806 8666 8807
rect 9030 9226 9058 9231
rect 8526 8801 8554 8806
rect 8134 8751 8135 8777
rect 8161 8751 8162 8777
rect 8134 8745 8162 8751
rect 7966 8722 7994 8727
rect 7350 8554 7378 8559
rect 7126 8553 7546 8554
rect 7126 8527 7351 8553
rect 7377 8527 7546 8553
rect 7126 8526 7546 8527
rect 7126 8441 7154 8526
rect 7350 8521 7378 8526
rect 7126 8415 7127 8441
rect 7153 8415 7154 8441
rect 7126 8409 7154 8415
rect 7518 8442 7546 8526
rect 7518 8414 7602 8442
rect 6790 8135 6791 8161
rect 6817 8135 6818 8161
rect 6790 8129 6818 8135
rect 5670 8073 5698 8078
rect 6734 8106 6762 8111
rect 6734 8059 6762 8078
rect 7574 8050 7602 8414
rect 7966 8105 7994 8694
rect 8414 8722 8442 8727
rect 8414 8675 8442 8694
rect 7966 8079 7967 8105
rect 7993 8079 7994 8105
rect 7966 8073 7994 8079
rect 8862 8442 8890 8447
rect 7630 8050 7658 8055
rect 7574 8049 7658 8050
rect 7574 8023 7631 8049
rect 7657 8023 7658 8049
rect 7574 8022 7658 8023
rect 7630 7658 7658 8022
rect 8694 7713 8722 7719
rect 8694 7687 8695 7713
rect 8721 7687 8722 7713
rect 7630 7625 7658 7630
rect 8022 7658 8050 7663
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 8022 7265 8050 7630
rect 8694 7574 8722 7687
rect 8862 7713 8890 8414
rect 9030 8105 9058 9198
rect 9030 8079 9031 8105
rect 9057 8079 9058 8105
rect 9030 8073 9058 8079
rect 9254 8105 9282 10038
rect 9478 9954 9506 10038
rect 9702 10066 9730 10822
rect 9758 10817 9786 10822
rect 10038 10794 10066 10799
rect 9758 10402 9786 10407
rect 9758 10355 9786 10374
rect 9870 10346 9898 10351
rect 9814 10345 9898 10346
rect 9814 10319 9871 10345
rect 9897 10319 9898 10345
rect 9814 10318 9898 10319
rect 9814 10122 9842 10318
rect 9870 10313 9898 10318
rect 10038 10345 10066 10766
rect 10038 10319 10039 10345
rect 10065 10319 10066 10345
rect 10038 10313 10066 10319
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9814 10094 9898 10122
rect 9702 10033 9730 10038
rect 9646 10010 9674 10015
rect 9646 9963 9674 9982
rect 9478 9921 9506 9926
rect 9478 9842 9506 9847
rect 9478 9618 9506 9814
rect 9814 9674 9842 9679
rect 9478 9561 9506 9590
rect 9646 9673 9842 9674
rect 9646 9647 9815 9673
rect 9841 9647 9842 9673
rect 9646 9646 9842 9647
rect 9646 9617 9674 9646
rect 9814 9641 9842 9646
rect 9646 9591 9647 9617
rect 9673 9591 9674 9617
rect 9590 9562 9618 9567
rect 9478 9535 9479 9561
rect 9505 9535 9506 9561
rect 9478 9529 9506 9535
rect 9534 9534 9590 9562
rect 9310 9506 9338 9511
rect 9310 9459 9338 9478
rect 9534 9170 9562 9534
rect 9590 9529 9618 9534
rect 9590 9282 9618 9287
rect 9646 9282 9674 9591
rect 9870 9618 9898 10094
rect 9870 9585 9898 9590
rect 9926 10066 9954 10071
rect 9926 9562 9954 10038
rect 10150 10066 10178 10071
rect 10150 10019 10178 10038
rect 10206 10065 10234 11046
rect 10262 11073 10290 11079
rect 10262 11047 10263 11073
rect 10289 11047 10290 11073
rect 10262 10402 10290 11047
rect 10262 10401 10346 10402
rect 10262 10375 10263 10401
rect 10289 10375 10346 10401
rect 10262 10374 10346 10375
rect 10262 10369 10290 10374
rect 10206 10039 10207 10065
rect 10233 10039 10234 10065
rect 10206 10033 10234 10039
rect 9982 10010 10010 10015
rect 9982 9730 10010 9982
rect 10094 10009 10122 10015
rect 10094 9983 10095 10009
rect 10121 9983 10122 10009
rect 10094 9842 10122 9983
rect 10094 9809 10122 9814
rect 10150 9730 10178 9735
rect 9982 9729 10178 9730
rect 9982 9703 9983 9729
rect 10009 9703 10151 9729
rect 10177 9703 10178 9729
rect 9982 9702 10178 9703
rect 9982 9697 10010 9702
rect 10150 9697 10178 9702
rect 9926 9529 9954 9534
rect 10206 9618 10234 9623
rect 10206 9561 10234 9590
rect 10206 9535 10207 9561
rect 10233 9535 10234 9561
rect 9870 9506 9898 9525
rect 9870 9473 9898 9478
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9702 9338 9730 9343
rect 9702 9291 9730 9310
rect 9590 9281 9674 9282
rect 9590 9255 9591 9281
rect 9617 9255 9674 9281
rect 9590 9254 9674 9255
rect 9590 9249 9618 9254
rect 10094 9226 10122 9231
rect 10206 9226 10234 9535
rect 10318 9338 10346 10374
rect 10374 10345 10402 11270
rect 10374 10319 10375 10345
rect 10401 10319 10402 10345
rect 10374 10313 10402 10319
rect 10318 9305 10346 9310
rect 10430 10009 10458 10015
rect 10430 9983 10431 10009
rect 10457 9983 10458 10009
rect 10122 9198 10234 9226
rect 10374 9282 10402 9287
rect 10374 9225 10402 9254
rect 10374 9199 10375 9225
rect 10401 9199 10402 9225
rect 10094 9179 10122 9198
rect 10374 9193 10402 9199
rect 10430 9226 10458 9983
rect 10542 9226 10570 11326
rect 10598 11074 10626 11494
rect 10598 11041 10626 11046
rect 10710 10906 10738 11886
rect 10766 11802 10794 12278
rect 10822 12273 10850 12278
rect 10878 12138 10906 12334
rect 11102 12306 11130 12334
rect 11102 12278 11186 12306
rect 10934 12250 10962 12255
rect 10934 12249 11130 12250
rect 10934 12223 10935 12249
rect 10961 12223 11130 12249
rect 10934 12222 11130 12223
rect 10934 12217 10962 12222
rect 10878 12110 10962 12138
rect 10934 12082 10962 12110
rect 10990 12082 11018 12087
rect 10934 12081 11018 12082
rect 10934 12055 10991 12081
rect 11017 12055 11018 12081
rect 10934 12054 11018 12055
rect 10990 12049 11018 12054
rect 10822 11970 10850 11975
rect 10934 11970 10962 11975
rect 10822 11969 10934 11970
rect 10822 11943 10823 11969
rect 10849 11943 10934 11969
rect 10822 11942 10934 11943
rect 10822 11937 10850 11942
rect 10822 11858 10850 11863
rect 10850 11830 10906 11858
rect 10822 11825 10850 11830
rect 10766 11130 10794 11774
rect 10766 11097 10794 11102
rect 10822 11410 10850 11415
rect 10710 10873 10738 10878
rect 10654 10402 10682 10407
rect 10654 10355 10682 10374
rect 10822 10121 10850 11382
rect 10878 11185 10906 11830
rect 10934 11746 10962 11942
rect 10934 11718 11018 11746
rect 10934 11521 10962 11527
rect 10934 11495 10935 11521
rect 10961 11495 10962 11521
rect 10934 11241 10962 11495
rect 10934 11215 10935 11241
rect 10961 11215 10962 11241
rect 10934 11209 10962 11215
rect 10878 11159 10879 11185
rect 10905 11159 10906 11185
rect 10878 11153 10906 11159
rect 10934 10794 10962 10799
rect 10990 10794 11018 11718
rect 11102 11242 11130 12222
rect 11158 11913 11186 12278
rect 11158 11887 11159 11913
rect 11185 11887 11186 11913
rect 11158 11881 11186 11887
rect 11102 11209 11130 11214
rect 11158 11466 11186 11471
rect 11158 11185 11186 11438
rect 11158 11159 11159 11185
rect 11185 11159 11186 11185
rect 11158 11153 11186 11159
rect 11214 11186 11242 12670
rect 11326 12586 11354 13119
rect 11326 12553 11354 12558
rect 11494 13146 11522 13175
rect 11326 12474 11354 12479
rect 11494 12474 11522 13118
rect 11326 12473 11522 12474
rect 11326 12447 11327 12473
rect 11353 12447 11522 12473
rect 11326 12446 11522 12447
rect 11718 13145 11746 13151
rect 11718 13119 11719 13145
rect 11745 13119 11746 13145
rect 11326 12441 11354 12446
rect 11438 12361 11466 12367
rect 11438 12335 11439 12361
rect 11465 12335 11466 12361
rect 11270 11969 11298 11975
rect 11270 11943 11271 11969
rect 11297 11943 11298 11969
rect 11270 11410 11298 11943
rect 11438 11970 11466 12335
rect 11718 12082 11746 13119
rect 12782 12809 12810 13454
rect 13230 13258 13258 13263
rect 13230 13211 13258 13230
rect 13678 13258 13706 13566
rect 20006 13593 20034 13599
rect 20006 13567 20007 13593
rect 20033 13567 20034 13593
rect 18830 13538 18858 13543
rect 18830 13491 18858 13510
rect 13678 13225 13706 13230
rect 13902 13482 13930 13487
rect 13902 13425 13930 13454
rect 13902 13399 13903 13425
rect 13929 13399 13930 13425
rect 12782 12783 12783 12809
rect 12809 12783 12810 12809
rect 12782 12777 12810 12783
rect 13118 13145 13146 13151
rect 13118 13119 13119 13145
rect 13145 13119 13146 13145
rect 13118 12753 13146 13119
rect 13118 12727 13119 12753
rect 13145 12727 13146 12753
rect 13118 12721 13146 12727
rect 13286 13145 13314 13151
rect 13286 13119 13287 13145
rect 13313 13119 13314 13145
rect 12838 12697 12866 12703
rect 12838 12671 12839 12697
rect 12865 12671 12866 12697
rect 12390 12586 12418 12591
rect 11718 12049 11746 12054
rect 12278 12082 12306 12087
rect 11438 11937 11466 11942
rect 11606 11969 11634 11975
rect 11606 11943 11607 11969
rect 11633 11943 11634 11969
rect 11606 11914 11634 11943
rect 12278 11969 12306 12054
rect 12278 11943 12279 11969
rect 12305 11943 12306 11969
rect 12278 11937 12306 11943
rect 11494 11857 11522 11863
rect 11494 11831 11495 11857
rect 11521 11831 11522 11857
rect 11494 11802 11522 11831
rect 11494 11769 11522 11774
rect 11326 11690 11354 11695
rect 11606 11690 11634 11886
rect 12390 11857 12418 12558
rect 12838 12474 12866 12671
rect 12950 12698 12978 12703
rect 12950 12651 12978 12670
rect 12838 12441 12866 12446
rect 13062 12641 13090 12647
rect 13062 12615 13063 12641
rect 13089 12615 13090 12641
rect 12670 12362 12698 12367
rect 12446 11914 12474 11919
rect 12446 11867 12474 11886
rect 12390 11831 12391 11857
rect 12417 11831 12418 11857
rect 11326 11577 11354 11662
rect 11326 11551 11327 11577
rect 11353 11551 11354 11577
rect 11326 11545 11354 11551
rect 11382 11662 11634 11690
rect 12054 11690 12082 11695
rect 11270 11377 11298 11382
rect 11214 11153 11242 11158
rect 11046 11130 11074 11135
rect 11046 11129 11130 11130
rect 11046 11103 11047 11129
rect 11073 11103 11130 11129
rect 11046 11102 11130 11103
rect 11046 11097 11074 11102
rect 11102 11018 11130 11102
rect 11102 10985 11130 10990
rect 10962 10766 11018 10794
rect 11158 10906 11186 10911
rect 10934 10761 10962 10766
rect 10822 10095 10823 10121
rect 10849 10095 10850 10121
rect 10822 10089 10850 10095
rect 11158 10290 11186 10878
rect 11158 10121 11186 10262
rect 11382 10234 11410 11662
rect 12054 11643 12082 11662
rect 11494 11577 11522 11583
rect 11494 11551 11495 11577
rect 11521 11551 11522 11577
rect 11494 11522 11522 11551
rect 11494 11489 11522 11494
rect 11606 11577 11634 11583
rect 11606 11551 11607 11577
rect 11633 11551 11634 11577
rect 11606 11410 11634 11551
rect 11718 11577 11746 11583
rect 11718 11551 11719 11577
rect 11745 11551 11746 11577
rect 11662 11521 11690 11527
rect 11662 11495 11663 11521
rect 11689 11495 11690 11521
rect 11662 11466 11690 11495
rect 11662 11433 11690 11438
rect 11606 11377 11634 11382
rect 11718 11298 11746 11551
rect 11774 11577 11802 11583
rect 11774 11551 11775 11577
rect 11801 11551 11802 11577
rect 11774 11354 11802 11551
rect 11774 11321 11802 11326
rect 11718 11265 11746 11270
rect 11550 11242 11578 11247
rect 11550 11186 11578 11214
rect 11718 11186 11746 11191
rect 11550 11185 11690 11186
rect 11550 11159 11551 11185
rect 11577 11159 11690 11185
rect 11550 11158 11690 11159
rect 11550 11153 11578 11158
rect 11438 11074 11466 11079
rect 11438 11027 11466 11046
rect 11606 11073 11634 11079
rect 11606 11047 11607 11073
rect 11633 11047 11634 11073
rect 11494 10793 11522 10799
rect 11494 10767 11495 10793
rect 11521 10767 11522 10793
rect 11494 10346 11522 10767
rect 11494 10313 11522 10318
rect 11382 10206 11578 10234
rect 11158 10095 11159 10121
rect 11185 10095 11186 10121
rect 11158 10089 11186 10095
rect 10654 10009 10682 10015
rect 10654 9983 10655 10009
rect 10681 9983 10682 10009
rect 10654 9898 10682 9983
rect 10766 10009 10794 10015
rect 10766 9983 10767 10009
rect 10793 9983 10794 10009
rect 10766 9954 10794 9983
rect 10766 9921 10794 9926
rect 10990 10009 11018 10015
rect 10990 9983 10991 10009
rect 11017 9983 11018 10009
rect 10654 9617 10682 9870
rect 10990 9674 11018 9983
rect 11102 10009 11130 10015
rect 11102 9983 11103 10009
rect 11129 9983 11130 10009
rect 11102 9954 11130 9983
rect 11102 9921 11130 9926
rect 11270 10009 11298 10015
rect 11270 9983 11271 10009
rect 11297 9983 11298 10009
rect 10990 9641 11018 9646
rect 11046 9730 11074 9735
rect 10766 9618 10794 9623
rect 10654 9591 10655 9617
rect 10681 9591 10682 9617
rect 10654 9585 10682 9591
rect 10710 9590 10766 9618
rect 10710 9506 10738 9590
rect 10766 9585 10794 9590
rect 11046 9617 11074 9702
rect 11046 9591 11047 9617
rect 11073 9591 11074 9617
rect 11046 9585 11074 9591
rect 10822 9562 10850 9567
rect 10542 9198 10626 9226
rect 10430 9193 10458 9198
rect 9646 9170 9674 9175
rect 9534 9142 9618 9170
rect 9590 8497 9618 9142
rect 9590 8471 9591 8497
rect 9617 8471 9618 8497
rect 9590 8465 9618 8471
rect 9646 8497 9674 9142
rect 10598 8666 10626 9198
rect 10710 9002 10738 9478
rect 10766 9505 10794 9511
rect 10766 9479 10767 9505
rect 10793 9479 10794 9505
rect 10766 9338 10794 9479
rect 10766 9305 10794 9310
rect 10822 9282 10850 9534
rect 11270 9561 11298 9983
rect 11494 9898 11522 9903
rect 11270 9535 11271 9561
rect 11297 9535 11298 9561
rect 11270 9529 11298 9535
rect 11326 9870 11494 9898
rect 11046 9506 11074 9511
rect 10822 9058 10850 9254
rect 10878 9281 10906 9287
rect 10878 9255 10879 9281
rect 10905 9255 10906 9281
rect 10878 9226 10906 9255
rect 10878 9193 10906 9198
rect 10990 9281 11018 9287
rect 10990 9255 10991 9281
rect 11017 9255 11018 9281
rect 10990 9226 11018 9255
rect 11046 9281 11074 9478
rect 11046 9255 11047 9281
rect 11073 9255 11074 9281
rect 11046 9249 11074 9255
rect 11102 9505 11130 9511
rect 11102 9479 11103 9505
rect 11129 9479 11130 9505
rect 10990 9193 11018 9198
rect 10822 9030 10906 9058
rect 10710 8974 10850 9002
rect 10822 8833 10850 8974
rect 10878 8889 10906 9030
rect 10878 8863 10879 8889
rect 10905 8863 10906 8889
rect 10878 8857 10906 8863
rect 11102 8834 11130 9479
rect 11158 9506 11186 9511
rect 11158 9459 11186 9478
rect 11270 8946 11298 8951
rect 11270 8834 11298 8918
rect 10822 8807 10823 8833
rect 10849 8807 10850 8833
rect 10822 8801 10850 8807
rect 10934 8806 11102 8834
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9646 8471 9647 8497
rect 9673 8471 9674 8497
rect 9646 8465 9674 8471
rect 9310 8442 9338 8447
rect 9310 8395 9338 8414
rect 9534 8441 9562 8447
rect 9534 8415 9535 8441
rect 9561 8415 9562 8441
rect 9534 8218 9562 8415
rect 10374 8442 10402 8447
rect 9534 8190 9954 8218
rect 9254 8079 9255 8105
rect 9281 8079 9282 8105
rect 8862 7687 8863 7713
rect 8889 7687 8890 7713
rect 8862 7681 8890 7687
rect 9198 7938 9226 7943
rect 8358 7546 8722 7574
rect 8358 7321 8386 7546
rect 8358 7295 8359 7321
rect 8385 7295 8386 7321
rect 8358 7289 8386 7295
rect 8022 7239 8023 7265
rect 8049 7239 8050 7265
rect 8022 7233 8050 7239
rect 9198 6985 9226 7910
rect 9254 7658 9282 8079
rect 9926 8049 9954 8190
rect 10318 8162 10346 8167
rect 9926 8023 9927 8049
rect 9953 8023 9954 8049
rect 9926 8017 9954 8023
rect 10094 8134 10318 8162
rect 10094 8049 10122 8134
rect 10318 8115 10346 8134
rect 10094 8023 10095 8049
rect 10121 8023 10122 8049
rect 10094 8017 10122 8023
rect 10374 8049 10402 8414
rect 10542 8442 10570 8447
rect 10542 8395 10570 8414
rect 10598 8441 10626 8638
rect 10598 8415 10599 8441
rect 10625 8415 10626 8441
rect 10598 8409 10626 8415
rect 10710 8441 10738 8447
rect 10710 8415 10711 8441
rect 10737 8415 10738 8441
rect 10654 8385 10682 8391
rect 10654 8359 10655 8385
rect 10681 8359 10682 8385
rect 10374 8023 10375 8049
rect 10401 8023 10402 8049
rect 10374 8017 10402 8023
rect 10486 8162 10514 8167
rect 10038 7938 10066 7957
rect 10038 7905 10066 7910
rect 10318 7938 10346 7943
rect 10318 7891 10346 7910
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9702 7714 9730 7719
rect 9702 7667 9730 7686
rect 9310 7658 9338 7663
rect 9282 7657 9338 7658
rect 9282 7631 9311 7657
rect 9337 7631 9338 7657
rect 9282 7630 9338 7631
rect 9254 7611 9282 7630
rect 9310 7574 9338 7630
rect 10206 7602 10234 7607
rect 9310 7546 9394 7574
rect 9366 7154 9394 7546
rect 9366 7121 9394 7126
rect 9422 7321 9450 7327
rect 9422 7295 9423 7321
rect 9449 7295 9450 7321
rect 9198 6959 9199 6985
rect 9225 6959 9226 6985
rect 9198 6953 9226 6959
rect 9142 6818 9170 6823
rect 9142 6771 9170 6790
rect 9422 6818 9450 7295
rect 9646 7154 9674 7159
rect 9646 7107 9674 7126
rect 9814 7154 9842 7159
rect 9814 6873 9842 7126
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 10206 6929 10234 7574
rect 10486 7266 10514 8134
rect 10654 8049 10682 8359
rect 10710 8162 10738 8415
rect 10710 8129 10738 8134
rect 10766 8441 10794 8447
rect 10766 8415 10767 8441
rect 10793 8415 10794 8441
rect 10654 8023 10655 8049
rect 10681 8023 10682 8049
rect 10654 8017 10682 8023
rect 10654 7937 10682 7943
rect 10654 7911 10655 7937
rect 10681 7911 10682 7937
rect 10654 7714 10682 7911
rect 10654 7681 10682 7686
rect 10766 7601 10794 8415
rect 10934 8386 10962 8806
rect 11102 8801 11130 8806
rect 11158 8833 11298 8834
rect 11158 8807 11271 8833
rect 11297 8807 11298 8833
rect 11158 8806 11298 8807
rect 10822 8358 10962 8386
rect 10990 8721 11018 8727
rect 10990 8695 10991 8721
rect 11017 8695 11018 8721
rect 10990 8442 11018 8695
rect 11158 8554 11186 8806
rect 11270 8801 11298 8806
rect 10822 8161 10850 8358
rect 10822 8135 10823 8161
rect 10849 8135 10850 8161
rect 10822 7658 10850 8135
rect 10934 8050 10962 8055
rect 10934 8003 10962 8022
rect 10990 7714 11018 8414
rect 11046 8553 11186 8554
rect 11046 8527 11159 8553
rect 11185 8527 11186 8553
rect 11046 8526 11186 8527
rect 11046 8049 11074 8526
rect 11158 8521 11186 8526
rect 11326 8777 11354 9870
rect 11494 9865 11522 9870
rect 11550 9226 11578 10206
rect 11326 8751 11327 8777
rect 11353 8751 11354 8777
rect 11046 8023 11047 8049
rect 11073 8023 11074 8049
rect 11046 8017 11074 8023
rect 11326 8050 11354 8751
rect 11438 8778 11466 8783
rect 11438 8731 11466 8750
rect 11550 8610 11578 9198
rect 11550 8577 11578 8582
rect 11326 8017 11354 8022
rect 11102 7770 11130 7775
rect 11046 7714 11074 7719
rect 10990 7686 11046 7714
rect 11046 7681 11074 7686
rect 11102 7713 11130 7742
rect 11550 7770 11578 7775
rect 11606 7770 11634 11047
rect 11662 10906 11690 11158
rect 11718 11139 11746 11158
rect 11718 11074 11746 11079
rect 11718 11018 11746 11046
rect 11998 11073 12026 11079
rect 11998 11047 11999 11073
rect 12025 11047 12026 11073
rect 11718 10990 11802 11018
rect 11718 10906 11746 10911
rect 11662 10905 11746 10906
rect 11662 10879 11719 10905
rect 11745 10879 11746 10905
rect 11662 10878 11746 10879
rect 11718 10873 11746 10878
rect 11662 10794 11690 10799
rect 11774 10794 11802 10990
rect 11662 10747 11690 10766
rect 11718 10766 11802 10794
rect 11830 10793 11858 10799
rect 11830 10767 11831 10793
rect 11857 10767 11858 10793
rect 11718 9898 11746 10766
rect 11830 10122 11858 10767
rect 11942 10793 11970 10799
rect 11942 10767 11943 10793
rect 11969 10767 11970 10793
rect 11942 10738 11970 10767
rect 11998 10794 12026 11047
rect 12166 11074 12194 11079
rect 12166 11027 12194 11046
rect 11998 10761 12026 10766
rect 11942 10705 11970 10710
rect 12334 10738 12362 10743
rect 12222 10122 12250 10127
rect 11830 10121 12250 10122
rect 11830 10095 12223 10121
rect 12249 10095 12250 10121
rect 11830 10094 12250 10095
rect 11830 9953 11858 10094
rect 12222 10089 12250 10094
rect 12278 10122 12306 10127
rect 12278 10065 12306 10094
rect 12278 10039 12279 10065
rect 12305 10039 12306 10065
rect 11942 10010 11970 10015
rect 11942 9963 11970 9982
rect 11830 9927 11831 9953
rect 11857 9927 11858 9953
rect 11830 9921 11858 9927
rect 11718 9851 11746 9870
rect 12278 9730 12306 10039
rect 11886 9702 12306 9730
rect 11830 9618 11858 9623
rect 11830 9571 11858 9590
rect 11830 9282 11858 9287
rect 11830 9235 11858 9254
rect 11886 9281 11914 9702
rect 11942 9506 11970 9511
rect 11942 9459 11970 9478
rect 11886 9255 11887 9281
rect 11913 9255 11914 9281
rect 11886 9249 11914 9255
rect 11830 9114 11858 9119
rect 11830 9067 11858 9086
rect 11942 8834 11970 8839
rect 11942 8787 11970 8806
rect 12054 8778 12082 8783
rect 12054 8731 12082 8750
rect 11942 8666 11970 8671
rect 11942 8105 11970 8638
rect 12110 8554 12138 9702
rect 12278 9618 12306 9623
rect 12278 9571 12306 9590
rect 12334 9506 12362 10710
rect 12390 10402 12418 11831
rect 12670 11690 12698 12334
rect 13006 12305 13034 12311
rect 13006 12279 13007 12305
rect 13033 12279 13034 12305
rect 13006 12025 13034 12279
rect 13006 11999 13007 12025
rect 13033 11999 13034 12025
rect 13006 11993 13034 11999
rect 13062 12082 13090 12615
rect 13286 12642 13314 13119
rect 13286 12609 13314 12614
rect 13902 13145 13930 13399
rect 13902 13119 13903 13145
rect 13929 13119 13930 13145
rect 12670 11657 12698 11662
rect 12838 11969 12866 11975
rect 12838 11943 12839 11969
rect 12865 11943 12866 11969
rect 12838 11689 12866 11943
rect 13062 11914 13090 12054
rect 13342 12474 13370 12479
rect 13342 12081 13370 12446
rect 13902 12362 13930 13119
rect 18830 13146 18858 13151
rect 18830 13099 18858 13118
rect 20006 13146 20034 13567
rect 20006 13113 20034 13118
rect 14294 13090 14322 13095
rect 14126 13089 14322 13090
rect 14126 13063 14295 13089
rect 14321 13063 14322 13089
rect 14126 13062 14322 13063
rect 14126 12865 14154 13062
rect 14294 13057 14322 13062
rect 15358 13090 15386 13095
rect 14126 12839 14127 12865
rect 14153 12839 14154 12865
rect 14126 12833 14154 12839
rect 14238 12754 14266 12759
rect 14238 12707 14266 12726
rect 14742 12754 14770 12759
rect 14742 12707 14770 12726
rect 14574 12697 14602 12703
rect 14574 12671 14575 12697
rect 14601 12671 14602 12697
rect 13342 12055 13343 12081
rect 13369 12055 13370 12081
rect 13342 12049 13370 12055
rect 13846 12334 13902 12362
rect 13846 12025 13874 12334
rect 13902 12329 13930 12334
rect 13958 12641 13986 12647
rect 13958 12615 13959 12641
rect 13985 12615 13986 12641
rect 13958 12474 13986 12615
rect 14070 12642 14098 12647
rect 14574 12642 14602 12671
rect 14630 12698 14658 12703
rect 14630 12651 14658 12670
rect 15358 12698 15386 13062
rect 15358 12665 15386 12670
rect 15582 13089 15610 13095
rect 15582 13063 15583 13089
rect 15609 13063 15610 13089
rect 14070 12641 14154 12642
rect 14070 12615 14071 12641
rect 14097 12615 14154 12641
rect 14070 12614 14154 12615
rect 14070 12609 14098 12614
rect 13846 11999 13847 12025
rect 13873 11999 13874 12025
rect 13846 11993 13874 11999
rect 13118 11914 13146 11919
rect 13062 11913 13146 11914
rect 13062 11887 13119 11913
rect 13145 11887 13146 11913
rect 13062 11886 13146 11887
rect 13118 11881 13146 11886
rect 13286 11914 13314 11919
rect 13958 11914 13986 12446
rect 14070 12305 14098 12311
rect 14070 12279 14071 12305
rect 14097 12279 14098 12305
rect 14070 12250 14098 12279
rect 14014 11914 14042 11919
rect 13958 11913 14042 11914
rect 13958 11887 14015 11913
rect 14041 11887 14042 11913
rect 13958 11886 14042 11887
rect 13286 11867 13314 11886
rect 14014 11881 14042 11886
rect 13006 11858 13034 11863
rect 13006 11857 13090 11858
rect 13006 11831 13007 11857
rect 13033 11831 13090 11857
rect 13006 11830 13090 11831
rect 13006 11825 13034 11830
rect 12838 11663 12839 11689
rect 12865 11663 12866 11689
rect 12838 11657 12866 11663
rect 12894 11633 12922 11639
rect 12894 11607 12895 11633
rect 12921 11607 12922 11633
rect 12782 11577 12810 11583
rect 12782 11551 12783 11577
rect 12809 11551 12810 11577
rect 12726 11298 12754 11303
rect 12390 10369 12418 10374
rect 12670 11073 12698 11079
rect 12670 11047 12671 11073
rect 12697 11047 12698 11073
rect 12558 10346 12586 10351
rect 12586 10318 12642 10346
rect 12558 10299 12586 10318
rect 12614 10009 12642 10318
rect 12670 10122 12698 11047
rect 12670 10089 12698 10094
rect 12614 9983 12615 10009
rect 12641 9983 12642 10009
rect 12614 9977 12642 9983
rect 12726 9786 12754 11270
rect 12782 11074 12810 11551
rect 12894 11130 12922 11607
rect 13006 11578 13034 11583
rect 13006 11531 13034 11550
rect 12950 11298 12978 11303
rect 13062 11298 13090 11830
rect 13342 11857 13370 11863
rect 13342 11831 13343 11857
rect 13369 11831 13370 11857
rect 13174 11578 13202 11583
rect 13174 11531 13202 11550
rect 13118 11298 13146 11303
rect 12978 11270 13034 11298
rect 13062 11270 13118 11298
rect 12950 11265 12978 11270
rect 13006 11186 13034 11270
rect 13118 11251 13146 11270
rect 13062 11186 13090 11191
rect 13342 11186 13370 11831
rect 14070 11634 14098 12222
rect 14126 11970 14154 12614
rect 14294 12362 14322 12367
rect 14294 12315 14322 12334
rect 14182 12306 14210 12311
rect 14182 12081 14210 12278
rect 14182 12055 14183 12081
rect 14209 12055 14210 12081
rect 14182 12049 14210 12055
rect 14294 11970 14322 11975
rect 14126 11942 14210 11970
rect 14070 11601 14098 11606
rect 14126 11857 14154 11863
rect 14126 11831 14127 11857
rect 14153 11831 14154 11857
rect 13006 11185 13370 11186
rect 13006 11159 13063 11185
rect 13089 11159 13370 11185
rect 13006 11158 13370 11159
rect 13566 11298 13594 11303
rect 13062 11153 13090 11158
rect 12894 11097 12922 11102
rect 13566 11129 13594 11270
rect 13566 11103 13567 11129
rect 13593 11103 13594 11129
rect 13566 11097 13594 11103
rect 13622 11241 13650 11247
rect 13622 11215 13623 11241
rect 13649 11215 13650 11241
rect 12782 10794 12810 11046
rect 12838 11073 12866 11079
rect 12838 11047 12839 11073
rect 12865 11047 12866 11073
rect 12838 11018 12866 11047
rect 13118 11073 13146 11079
rect 13118 11047 13119 11073
rect 13145 11047 13146 11073
rect 13118 11018 13146 11047
rect 12838 10990 13146 11018
rect 12782 10747 12810 10766
rect 12894 10849 12922 10855
rect 12894 10823 12895 10849
rect 12921 10823 12922 10849
rect 12894 10010 12922 10823
rect 12950 10849 12978 10855
rect 12950 10823 12951 10849
rect 12977 10823 12978 10849
rect 12950 10402 12978 10823
rect 12950 10369 12978 10374
rect 13118 10793 13146 10990
rect 13342 11018 13370 11023
rect 13118 10767 13119 10793
rect 13145 10767 13146 10793
rect 12726 9758 12866 9786
rect 12670 9730 12698 9735
rect 12334 9473 12362 9478
rect 12558 9617 12586 9623
rect 12558 9591 12559 9617
rect 12585 9591 12586 9617
rect 12558 9562 12586 9591
rect 12502 9282 12530 9287
rect 12558 9282 12586 9534
rect 12614 9561 12642 9567
rect 12614 9535 12615 9561
rect 12641 9535 12642 9561
rect 12614 9394 12642 9535
rect 12614 9361 12642 9366
rect 12670 9338 12698 9702
rect 12670 9291 12698 9310
rect 12726 9674 12754 9679
rect 12726 9618 12754 9646
rect 12782 9618 12810 9623
rect 12726 9617 12810 9618
rect 12726 9591 12783 9617
rect 12809 9591 12810 9617
rect 12726 9590 12810 9591
rect 12558 9254 12642 9282
rect 12502 8889 12530 9254
rect 12614 9225 12642 9254
rect 12614 9199 12615 9225
rect 12641 9199 12642 9225
rect 12614 9193 12642 9199
rect 12502 8863 12503 8889
rect 12529 8863 12530 8889
rect 12502 8857 12530 8863
rect 12222 8834 12250 8839
rect 12222 8787 12250 8806
rect 12166 8722 12194 8727
rect 12166 8675 12194 8694
rect 12166 8554 12194 8559
rect 12110 8553 12194 8554
rect 12110 8527 12167 8553
rect 12193 8527 12194 8553
rect 12110 8526 12194 8527
rect 11942 8079 11943 8105
rect 11969 8079 11970 8105
rect 11942 8073 11970 8079
rect 12166 8105 12194 8526
rect 12334 8498 12362 8503
rect 12334 8451 12362 8470
rect 12670 8442 12698 8447
rect 12670 8395 12698 8414
rect 12726 8162 12754 9590
rect 12782 9585 12810 9590
rect 12838 9562 12866 9758
rect 12894 9674 12922 9982
rect 13118 10346 13146 10767
rect 13174 10962 13202 10967
rect 13174 10737 13202 10934
rect 13342 10906 13370 10990
rect 13454 10906 13482 10911
rect 13174 10711 13175 10737
rect 13201 10711 13202 10737
rect 13174 10705 13202 10711
rect 13230 10905 13482 10906
rect 13230 10879 13455 10905
rect 13481 10879 13482 10905
rect 13230 10878 13482 10879
rect 12894 9646 13090 9674
rect 12894 9562 12922 9567
rect 12838 9561 12922 9562
rect 12838 9535 12895 9561
rect 12921 9535 12922 9561
rect 12838 9534 12922 9535
rect 12894 9529 12922 9534
rect 12950 9506 12978 9511
rect 12950 9459 12978 9478
rect 13006 9505 13034 9511
rect 13006 9479 13007 9505
rect 13033 9479 13034 9505
rect 12894 9450 12922 9455
rect 12894 8834 12922 9422
rect 13006 9394 13034 9479
rect 13006 9361 13034 9366
rect 13062 9282 13090 9646
rect 13118 9617 13146 10318
rect 13118 9591 13119 9617
rect 13145 9591 13146 9617
rect 13118 9585 13146 9591
rect 13062 9235 13090 9254
rect 13174 9226 13202 9231
rect 13174 9179 13202 9198
rect 13230 9058 13258 10878
rect 13454 10873 13482 10878
rect 13510 10849 13538 10855
rect 13510 10823 13511 10849
rect 13537 10823 13538 10849
rect 13342 10794 13370 10799
rect 13342 10402 13370 10766
rect 13510 10738 13538 10823
rect 13622 10850 13650 11215
rect 13846 11186 13874 11191
rect 13846 11139 13874 11158
rect 13678 11074 13706 11079
rect 13678 11073 13762 11074
rect 13678 11047 13679 11073
rect 13705 11047 13762 11073
rect 13678 11046 13762 11047
rect 13678 11041 13706 11046
rect 13622 10817 13650 10822
rect 13678 10794 13706 10799
rect 13678 10747 13706 10766
rect 13538 10710 13650 10738
rect 13510 10705 13538 10710
rect 13454 10402 13482 10407
rect 13342 10401 13482 10402
rect 13342 10375 13455 10401
rect 13481 10375 13482 10401
rect 13342 10374 13482 10375
rect 13454 10369 13482 10374
rect 13566 10346 13594 10351
rect 13566 10299 13594 10318
rect 13622 10345 13650 10710
rect 13734 10737 13762 11046
rect 14126 10962 14154 11831
rect 14182 11186 14210 11942
rect 14294 11923 14322 11942
rect 14574 11969 14602 12614
rect 15582 12362 15610 13063
rect 19950 13089 19978 13095
rect 19950 13063 19951 13089
rect 19977 13063 19978 13089
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 19950 12810 19978 13063
rect 19950 12777 19978 12782
rect 20006 12809 20034 12815
rect 20006 12783 20007 12809
rect 20033 12783 20034 12809
rect 18830 12753 18858 12759
rect 18830 12727 18831 12753
rect 18857 12727 18858 12753
rect 18830 12418 18858 12727
rect 20006 12474 20034 12783
rect 20006 12441 20034 12446
rect 18830 12385 18858 12390
rect 15582 12329 15610 12334
rect 15918 12362 15946 12367
rect 14630 12306 14658 12311
rect 14630 12259 14658 12278
rect 15694 12306 15722 12311
rect 14574 11943 14575 11969
rect 14601 11943 14602 11969
rect 14574 11937 14602 11943
rect 14742 11970 14770 11975
rect 14742 11923 14770 11942
rect 14630 11914 14658 11919
rect 14630 11867 14658 11886
rect 15694 11914 15722 12278
rect 15694 11881 15722 11886
rect 15918 12305 15946 12334
rect 15918 12279 15919 12305
rect 15945 12279 15946 12305
rect 14182 11153 14210 11158
rect 14126 10929 14154 10934
rect 14406 10850 14434 10855
rect 14406 10803 14434 10822
rect 13734 10711 13735 10737
rect 13761 10711 13762 10737
rect 13734 10705 13762 10711
rect 14014 10793 14042 10799
rect 14014 10767 14015 10793
rect 14041 10767 14042 10793
rect 13622 10319 13623 10345
rect 13649 10319 13650 10345
rect 13622 10313 13650 10319
rect 13846 10401 13874 10407
rect 13846 10375 13847 10401
rect 13873 10375 13874 10401
rect 13510 10289 13538 10295
rect 13510 10263 13511 10289
rect 13537 10263 13538 10289
rect 13510 10094 13538 10263
rect 13286 10066 13314 10071
rect 13286 9617 13314 10038
rect 13286 9591 13287 9617
rect 13313 9591 13314 9617
rect 13286 9585 13314 9591
rect 13398 10066 13538 10094
rect 13846 10066 13874 10375
rect 13398 9617 13426 10066
rect 13846 10033 13874 10038
rect 13398 9591 13399 9617
rect 13425 9591 13426 9617
rect 13398 9585 13426 9591
rect 13454 9561 13482 9567
rect 13454 9535 13455 9561
rect 13481 9535 13482 9561
rect 13454 9506 13482 9535
rect 13678 9562 13706 9567
rect 13958 9562 13986 9567
rect 13678 9561 13986 9562
rect 13678 9535 13679 9561
rect 13705 9535 13959 9561
rect 13985 9535 13986 9561
rect 13678 9534 13986 9535
rect 13678 9529 13706 9534
rect 13958 9529 13986 9534
rect 13454 9473 13482 9478
rect 13790 9450 13818 9455
rect 13566 9394 13594 9399
rect 13342 9338 13370 9343
rect 13370 9310 13482 9338
rect 13342 9305 13370 9310
rect 13454 9225 13482 9310
rect 13454 9199 13455 9225
rect 13481 9199 13482 9225
rect 13454 9193 13482 9199
rect 13510 9226 13538 9231
rect 13062 9030 13426 9058
rect 12950 8834 12978 8839
rect 12894 8833 12978 8834
rect 12894 8807 12951 8833
rect 12977 8807 12978 8833
rect 12894 8806 12978 8807
rect 12950 8801 12978 8806
rect 13006 8834 13034 8839
rect 13006 8787 13034 8806
rect 13062 8833 13090 9030
rect 13062 8807 13063 8833
rect 13089 8807 13090 8833
rect 13062 8801 13090 8807
rect 13286 8834 13314 8839
rect 13286 8787 13314 8806
rect 13398 8777 13426 9030
rect 13398 8751 13399 8777
rect 13425 8751 13426 8777
rect 13398 8745 13426 8751
rect 13510 8833 13538 9198
rect 13566 9225 13594 9366
rect 13734 9281 13762 9287
rect 13734 9255 13735 9281
rect 13761 9255 13762 9281
rect 13566 9199 13567 9225
rect 13593 9199 13594 9225
rect 13566 9193 13594 9199
rect 13678 9225 13706 9231
rect 13678 9199 13679 9225
rect 13705 9199 13706 9225
rect 13678 8946 13706 9199
rect 13734 9226 13762 9255
rect 13790 9281 13818 9422
rect 13790 9255 13791 9281
rect 13817 9255 13818 9281
rect 13790 9249 13818 9255
rect 13734 9193 13762 9198
rect 14014 9225 14042 10767
rect 15470 10794 15498 10799
rect 15470 10737 15498 10766
rect 15694 10738 15722 10743
rect 15918 10738 15946 12279
rect 18830 12250 18858 12255
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 18830 11969 18858 12222
rect 18830 11943 18831 11969
rect 18857 11943 18858 11969
rect 18830 11937 18858 11943
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 20006 11802 20034 11999
rect 20006 11769 20034 11774
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 18830 11185 18858 11191
rect 18830 11159 18831 11185
rect 18857 11159 18858 11185
rect 18830 10794 18858 11159
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 18830 10761 18858 10766
rect 15470 10711 15471 10737
rect 15497 10711 15498 10737
rect 15470 10705 15498 10711
rect 15638 10737 15946 10738
rect 15638 10711 15695 10737
rect 15721 10711 15946 10737
rect 15638 10710 15946 10711
rect 15414 10066 15442 10071
rect 15414 10019 15442 10038
rect 14630 9953 14658 9959
rect 14630 9927 14631 9953
rect 14657 9927 14658 9953
rect 14630 9617 14658 9927
rect 15470 9953 15498 9959
rect 15470 9927 15471 9953
rect 15497 9927 15498 9953
rect 15470 9674 15498 9927
rect 15470 9641 15498 9646
rect 14630 9591 14631 9617
rect 14657 9591 14658 9617
rect 14126 9562 14154 9567
rect 14126 9515 14154 9534
rect 14014 9199 14015 9225
rect 14041 9199 14042 9225
rect 13678 8913 13706 8918
rect 13510 8807 13511 8833
rect 13537 8807 13538 8833
rect 12782 8722 12810 8727
rect 13006 8722 13034 8727
rect 12782 8721 12922 8722
rect 12782 8695 12783 8721
rect 12809 8695 12922 8721
rect 12782 8694 12922 8695
rect 12782 8689 12810 8694
rect 12726 8129 12754 8134
rect 12166 8079 12167 8105
rect 12193 8079 12194 8105
rect 12166 8073 12194 8079
rect 11578 7742 11634 7770
rect 12222 8049 12250 8055
rect 12894 8050 12922 8694
rect 12222 8023 12223 8049
rect 12249 8023 12250 8049
rect 12222 7770 12250 8023
rect 11550 7723 11578 7742
rect 12222 7737 12250 7742
rect 12614 8049 12922 8050
rect 12614 8023 12895 8049
rect 12921 8023 12922 8049
rect 12614 8022 12922 8023
rect 11102 7687 11103 7713
rect 11129 7687 11130 7713
rect 11102 7681 11130 7687
rect 11382 7714 11410 7719
rect 11382 7667 11410 7686
rect 11438 7713 11466 7719
rect 11438 7687 11439 7713
rect 11465 7687 11466 7713
rect 10822 7625 10850 7630
rect 10878 7657 10906 7663
rect 10878 7631 10879 7657
rect 10905 7631 10906 7657
rect 10766 7575 10767 7601
rect 10793 7575 10794 7601
rect 10654 7266 10682 7271
rect 10486 7265 10682 7266
rect 10486 7239 10655 7265
rect 10681 7239 10682 7265
rect 10486 7238 10682 7239
rect 10654 7233 10682 7238
rect 10206 6903 10207 6929
rect 10233 6903 10234 6929
rect 10206 6897 10234 6903
rect 10710 7153 10738 7159
rect 10710 7127 10711 7153
rect 10737 7127 10738 7153
rect 9814 6847 9815 6873
rect 9841 6847 9842 6873
rect 9814 6841 9842 6847
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 854 2450 882 2455
rect 854 2403 882 2422
rect 9422 2169 9450 6790
rect 10710 6818 10738 7127
rect 10710 6785 10738 6790
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 10766 4214 10794 7575
rect 10822 7266 10850 7271
rect 10878 7266 10906 7631
rect 11158 7658 11186 7663
rect 10990 7602 11018 7621
rect 11158 7611 11186 7630
rect 10990 7569 11018 7574
rect 11438 7574 11466 7687
rect 12614 7713 12642 8022
rect 12894 8017 12922 8022
rect 12950 8610 12978 8615
rect 12838 7938 12866 7943
rect 12838 7891 12866 7910
rect 12670 7770 12698 7775
rect 12670 7723 12698 7742
rect 12894 7770 12922 7775
rect 12950 7770 12978 8582
rect 13006 8497 13034 8694
rect 13006 8471 13007 8497
rect 13033 8471 13034 8497
rect 13006 8465 13034 8471
rect 13510 8498 13538 8807
rect 13118 8050 13146 8055
rect 13118 8003 13146 8022
rect 13510 7994 13538 8470
rect 14014 8442 14042 9199
rect 14350 9226 14378 9231
rect 14350 9179 14378 9198
rect 14630 9170 14658 9591
rect 14966 9562 14994 9567
rect 14966 9515 14994 9534
rect 14014 8409 14042 8414
rect 14070 8834 14098 8839
rect 14070 8385 14098 8806
rect 14630 8721 14658 9142
rect 15414 9169 15442 9175
rect 15414 9143 15415 9169
rect 15441 9143 15442 9169
rect 14910 9114 14938 9119
rect 14854 8946 14882 8951
rect 14854 8899 14882 8918
rect 14910 8889 14938 9086
rect 15414 9114 15442 9143
rect 15638 9170 15666 10710
rect 15694 10705 15722 10710
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 20006 10457 20034 10463
rect 20006 10431 20007 10457
rect 20033 10431 20034 10457
rect 18830 10401 18858 10407
rect 18830 10375 18831 10401
rect 18857 10375 18858 10401
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 16030 9674 16058 9679
rect 16030 9627 16058 9646
rect 18830 9674 18858 10375
rect 20006 10122 20034 10431
rect 20006 10089 20034 10094
rect 18830 9641 18858 9646
rect 18830 9226 18858 9231
rect 18830 9179 18858 9198
rect 15638 9123 15666 9142
rect 15414 9081 15442 9086
rect 20006 9114 20034 9119
rect 20006 9067 20034 9086
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 14910 8863 14911 8889
rect 14937 8863 14938 8889
rect 14910 8857 14938 8863
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 14630 8695 14631 8721
rect 14657 8695 14658 8721
rect 14070 8359 14071 8385
rect 14097 8359 14098 8385
rect 14070 8353 14098 8359
rect 14294 8442 14322 8447
rect 13510 7947 13538 7966
rect 13342 7937 13370 7943
rect 13342 7911 13343 7937
rect 13369 7911 13370 7937
rect 12894 7769 12978 7770
rect 12894 7743 12895 7769
rect 12921 7743 12978 7769
rect 12894 7742 12978 7743
rect 13006 7770 13034 7775
rect 12894 7737 12922 7742
rect 12614 7687 12615 7713
rect 12641 7687 12642 7713
rect 11438 7546 11522 7574
rect 10822 7265 10906 7266
rect 10822 7239 10823 7265
rect 10849 7239 10906 7265
rect 10822 7238 10906 7239
rect 10822 7233 10850 7238
rect 11494 7210 11522 7546
rect 12614 7546 12642 7687
rect 12614 7513 12642 7518
rect 11494 7177 11522 7182
rect 12390 7210 12418 7215
rect 10990 7154 11018 7159
rect 10990 7107 11018 7126
rect 11830 7154 11858 7159
rect 11830 6985 11858 7126
rect 11830 6959 11831 6985
rect 11857 6959 11858 6985
rect 11830 6953 11858 6959
rect 11606 6930 11634 6935
rect 11606 6929 11802 6930
rect 11606 6903 11607 6929
rect 11633 6903 11802 6929
rect 11606 6902 11802 6903
rect 11606 6897 11634 6902
rect 11438 6873 11466 6879
rect 11438 6847 11439 6873
rect 11465 6847 11466 6873
rect 11270 6818 11298 6823
rect 11438 6818 11466 6847
rect 11298 6790 11466 6818
rect 11270 4214 11298 6790
rect 10654 4186 10794 4214
rect 11102 4186 11298 4214
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 10430 2618 10458 2623
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9422 2143 9423 2169
rect 9449 2143 9450 2169
rect 9422 2137 9450 2143
rect 9422 2058 9450 2063
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 9422 400 9450 2030
rect 9926 2058 9954 2063
rect 9926 2011 9954 2030
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10430 400 10458 2590
rect 10654 2561 10682 4186
rect 10654 2535 10655 2561
rect 10681 2535 10682 2561
rect 10654 2529 10682 2535
rect 11102 2169 11130 4186
rect 11158 2618 11186 2623
rect 11158 2571 11186 2590
rect 11102 2143 11103 2169
rect 11129 2143 11130 2169
rect 11102 2137 11130 2143
rect 10766 2058 10794 2063
rect 10766 400 10794 2030
rect 11382 2058 11410 2063
rect 11382 2011 11410 2030
rect 11774 1777 11802 6902
rect 12054 6818 12082 6823
rect 12054 6481 12082 6790
rect 12390 6537 12418 7182
rect 12558 7210 12586 7215
rect 12558 7163 12586 7182
rect 12726 7210 12754 7215
rect 12894 7210 12922 7215
rect 12726 7209 12922 7210
rect 12726 7183 12727 7209
rect 12753 7183 12895 7209
rect 12921 7183 12922 7209
rect 12726 7182 12922 7183
rect 12726 7177 12754 7182
rect 12894 7177 12922 7182
rect 13006 6929 13034 7742
rect 13174 7601 13202 7607
rect 13174 7575 13175 7601
rect 13201 7575 13202 7601
rect 13062 7545 13090 7551
rect 13062 7519 13063 7545
rect 13089 7519 13090 7545
rect 13062 7378 13090 7519
rect 13174 7546 13202 7575
rect 13174 7513 13202 7518
rect 13062 7350 13314 7378
rect 13230 7265 13258 7271
rect 13230 7239 13231 7265
rect 13257 7239 13258 7265
rect 13230 7154 13258 7239
rect 13286 7266 13314 7350
rect 13342 7266 13370 7911
rect 13286 7265 13370 7266
rect 13286 7239 13343 7265
rect 13369 7239 13370 7265
rect 13286 7238 13370 7239
rect 13230 7121 13258 7126
rect 13006 6903 13007 6929
rect 13033 6903 13034 6929
rect 13006 6897 13034 6903
rect 12614 6873 12642 6879
rect 12614 6847 12615 6873
rect 12641 6847 12642 6873
rect 12614 6818 12642 6847
rect 12614 6785 12642 6790
rect 12390 6511 12391 6537
rect 12417 6511 12418 6537
rect 12390 6505 12418 6511
rect 13342 6538 13370 7238
rect 13566 7546 13594 7551
rect 13566 7209 13594 7518
rect 13566 7183 13567 7209
rect 13593 7183 13594 7209
rect 13566 7177 13594 7183
rect 13734 7154 13762 7159
rect 13734 7107 13762 7126
rect 14070 7154 14098 7159
rect 13734 6818 13762 6823
rect 13454 6538 13482 6543
rect 13342 6537 13482 6538
rect 13342 6511 13455 6537
rect 13481 6511 13482 6537
rect 13342 6510 13482 6511
rect 13454 6505 13482 6510
rect 13734 6537 13762 6790
rect 14070 6817 14098 7126
rect 14070 6791 14071 6817
rect 14097 6791 14098 6817
rect 14070 6785 14098 6791
rect 14294 6818 14322 8414
rect 14630 8442 14658 8695
rect 14630 8409 14658 8414
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 14294 6771 14322 6790
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 13734 6511 13735 6537
rect 13761 6511 13762 6537
rect 13734 6505 13762 6511
rect 12054 6455 12055 6481
rect 12081 6455 12082 6481
rect 12054 6449 12082 6455
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 20118 2449 20146 2455
rect 20118 2423 20119 2449
rect 20145 2423 20146 2449
rect 20118 2394 20146 2423
rect 20118 2361 20146 2366
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 11774 1751 11775 1777
rect 11801 1751 11802 1777
rect 11774 1745 11802 1751
rect 11102 1721 11130 1727
rect 11102 1695 11103 1721
rect 11129 1695 11130 1721
rect 11102 400 11130 1695
rect 9408 0 9464 400
rect 10416 0 10472 400
rect 10752 0 10808 400
rect 11088 0 11144 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 8414 18326 8442 18354
rect 9030 18353 9058 18354
rect 9030 18327 9031 18353
rect 9031 18327 9057 18353
rect 9057 18327 9058 18353
rect 9030 18326 9058 18327
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 7350 13790 7378 13818
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 2086 13454 2114 13482
rect 966 12782 994 12810
rect 966 11465 994 11466
rect 966 11439 967 11465
rect 967 11439 993 11465
rect 993 11439 994 11465
rect 966 11438 994 11439
rect 966 11241 994 11242
rect 966 11215 967 11241
rect 967 11215 993 11241
rect 993 11215 994 11241
rect 966 11214 994 11215
rect 7910 13817 7938 13818
rect 7910 13791 7911 13817
rect 7911 13791 7937 13817
rect 7937 13791 7938 13817
rect 7910 13790 7938 13791
rect 2142 13145 2170 13146
rect 2142 13119 2143 13145
rect 2143 13119 2169 13145
rect 2169 13119 2170 13145
rect 2142 13118 2170 13119
rect 6118 13118 6146 13146
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 6118 12670 6146 12698
rect 7798 13118 7826 13146
rect 7014 12614 7042 12642
rect 7406 12670 7434 12698
rect 7574 12558 7602 12586
rect 7630 12446 7658 12474
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 6734 11969 6762 11970
rect 6734 11943 6735 11969
rect 6735 11943 6761 11969
rect 6761 11943 6762 11969
rect 6734 11942 6762 11943
rect 2142 11577 2170 11578
rect 2142 11551 2143 11577
rect 2143 11551 2169 11577
rect 2169 11551 2170 11577
rect 2142 11550 2170 11551
rect 5838 11550 5866 11578
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 2142 11185 2170 11186
rect 2142 11159 2143 11185
rect 2143 11159 2169 11185
rect 2169 11159 2170 11185
rect 2142 11158 2170 11159
rect 5782 11158 5810 11186
rect 5782 11046 5810 11074
rect 6902 11913 6930 11914
rect 6902 11887 6903 11913
rect 6903 11887 6929 11913
rect 6929 11887 6930 11913
rect 6902 11886 6930 11887
rect 7294 11942 7322 11970
rect 7798 12614 7826 12642
rect 7406 11886 7434 11914
rect 7238 11718 7266 11746
rect 7462 11662 7490 11690
rect 6902 11382 6930 11410
rect 7294 11577 7322 11578
rect 7294 11551 7295 11577
rect 7295 11551 7321 11577
rect 7321 11551 7322 11577
rect 7294 11550 7322 11551
rect 7574 11494 7602 11522
rect 7630 11382 7658 11410
rect 7910 11718 7938 11746
rect 7742 11550 7770 11578
rect 7798 11494 7826 11522
rect 7742 11326 7770 11354
rect 7462 11073 7490 11074
rect 7462 11047 7463 11073
rect 7463 11047 7489 11073
rect 7489 11047 7490 11073
rect 7462 11046 7490 11047
rect 6790 10766 6818 10794
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 2086 10374 2114 10402
rect 966 10094 994 10122
rect 6342 10262 6370 10290
rect 6790 10289 6818 10290
rect 6790 10263 6791 10289
rect 6791 10263 6817 10289
rect 6817 10263 6818 10289
rect 6790 10262 6818 10263
rect 6846 10150 6874 10178
rect 2142 9926 2170 9954
rect 5278 9953 5306 9954
rect 5278 9927 5279 9953
rect 5279 9927 5305 9953
rect 5305 9927 5306 9953
rect 5278 9926 5306 9927
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 6790 9870 6818 9898
rect 6902 9729 6930 9730
rect 6902 9703 6903 9729
rect 6903 9703 6929 9729
rect 6929 9703 6930 9729
rect 6902 9702 6930 9703
rect 7294 10150 7322 10178
rect 6734 9142 6762 9170
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 966 8889 994 8890
rect 966 8863 967 8889
rect 967 8863 993 8889
rect 993 8863 994 8889
rect 966 8862 994 8863
rect 2142 8833 2170 8834
rect 2142 8807 2143 8833
rect 2143 8807 2169 8833
rect 2169 8807 2170 8833
rect 2142 8806 2170 8807
rect 5670 8806 5698 8834
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 7182 10038 7210 10066
rect 7798 10905 7826 10906
rect 7798 10879 7799 10905
rect 7799 10879 7825 10905
rect 7825 10879 7826 10905
rect 7798 10878 7826 10879
rect 7630 10766 7658 10794
rect 8134 13118 8162 13146
rect 8022 12838 8050 12866
rect 10598 18913 10626 18914
rect 10598 18887 10599 18913
rect 10599 18887 10625 18913
rect 10625 18887 10626 18913
rect 10598 18886 10626 18887
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 9422 18718 9450 18746
rect 9926 18745 9954 18746
rect 9926 18719 9927 18745
rect 9927 18719 9953 18745
rect 9953 18719 9954 18745
rect 9926 18718 9954 18719
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 9142 13398 9170 13426
rect 8694 13145 8722 13146
rect 8694 13119 8695 13145
rect 8695 13119 8721 13145
rect 8721 13119 8722 13145
rect 8694 13118 8722 13119
rect 8414 12838 8442 12866
rect 8246 12446 8274 12474
rect 8694 12473 8722 12474
rect 8694 12447 8695 12473
rect 8695 12447 8721 12473
rect 8721 12447 8722 12473
rect 8694 12446 8722 12447
rect 8862 11886 8890 11914
rect 9086 11830 9114 11858
rect 8806 11606 8834 11634
rect 9198 11913 9226 11914
rect 9198 11887 9199 11913
rect 9199 11887 9225 11913
rect 9225 11887 9226 11913
rect 9198 11886 9226 11887
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 9646 14014 9674 14042
rect 9310 13425 9338 13426
rect 9310 13399 9311 13425
rect 9311 13399 9337 13425
rect 9337 13399 9338 13425
rect 9310 13398 9338 13399
rect 10150 14041 10178 14042
rect 10150 14015 10151 14041
rect 10151 14015 10177 14041
rect 10177 14015 10178 14041
rect 10150 14014 10178 14015
rect 9646 13398 9674 13426
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9982 13089 10010 13090
rect 9982 13063 9983 13089
rect 9983 13063 10009 13089
rect 10009 13063 10010 13089
rect 9982 13062 10010 13063
rect 9646 12782 9674 12810
rect 8022 11550 8050 11578
rect 8302 11550 8330 11578
rect 8638 11577 8666 11578
rect 8638 11551 8639 11577
rect 8639 11551 8665 11577
rect 8665 11551 8666 11577
rect 8638 11550 8666 11551
rect 8918 11577 8946 11578
rect 8918 11551 8919 11577
rect 8919 11551 8945 11577
rect 8945 11551 8946 11577
rect 8918 11550 8946 11551
rect 9086 11494 9114 11522
rect 9086 11158 9114 11186
rect 7742 10345 7770 10346
rect 7742 10319 7743 10345
rect 7743 10319 7769 10345
rect 7769 10319 7770 10345
rect 7742 10318 7770 10319
rect 7798 10289 7826 10290
rect 7798 10263 7799 10289
rect 7799 10263 7825 10289
rect 7825 10263 7826 10289
rect 7798 10262 7826 10263
rect 7574 9617 7602 9618
rect 7574 9591 7575 9617
rect 7575 9591 7601 9617
rect 7601 9591 7602 9617
rect 7574 9590 7602 9591
rect 7182 9534 7210 9562
rect 7294 9337 7322 9338
rect 7294 9311 7295 9337
rect 7295 9311 7321 9337
rect 7321 9311 7322 9337
rect 7294 9310 7322 9311
rect 7686 9337 7714 9338
rect 7686 9311 7687 9337
rect 7687 9311 7713 9337
rect 7713 9311 7714 9337
rect 7686 9310 7714 9311
rect 7406 9225 7434 9226
rect 7406 9199 7407 9225
rect 7407 9199 7433 9225
rect 7433 9199 7434 9225
rect 7406 9198 7434 9199
rect 8302 11046 8330 11074
rect 9198 11577 9226 11578
rect 9198 11551 9199 11577
rect 9199 11551 9225 11577
rect 9225 11551 9226 11577
rect 9198 11550 9226 11551
rect 9478 11577 9506 11578
rect 9478 11551 9479 11577
rect 9479 11551 9505 11577
rect 9505 11551 9506 11577
rect 9478 11550 9506 11551
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 10094 11830 10122 11858
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 9870 11521 9898 11522
rect 9870 11495 9871 11521
rect 9871 11495 9897 11521
rect 9897 11495 9898 11521
rect 9870 11494 9898 11495
rect 9142 10878 9170 10906
rect 8414 10345 8442 10346
rect 8414 10319 8415 10345
rect 8415 10319 8441 10345
rect 8441 10319 8442 10345
rect 8414 10318 8442 10319
rect 8358 9953 8386 9954
rect 8358 9927 8359 9953
rect 8359 9927 8385 9953
rect 8385 9927 8386 9953
rect 8358 9926 8386 9927
rect 8974 10289 9002 10290
rect 8974 10263 8975 10289
rect 8975 10263 9001 10289
rect 9001 10263 9002 10289
rect 8974 10262 9002 10263
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 11438 19110 11466 19138
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 11774 18886 11802 18914
rect 10766 18718 10794 18746
rect 11382 18745 11410 18746
rect 11382 18719 11383 18745
rect 11383 18719 11409 18745
rect 11409 18719 11410 18745
rect 11382 18718 11410 18719
rect 10654 13873 10682 13874
rect 10654 13847 10655 13873
rect 10655 13847 10681 13873
rect 10681 13847 10682 13873
rect 10654 13846 10682 13847
rect 11046 13846 11074 13874
rect 11438 13846 11466 13874
rect 10654 13062 10682 13090
rect 11718 13873 11746 13874
rect 11718 13847 11719 13873
rect 11719 13847 11745 13873
rect 11745 13847 11746 13873
rect 11718 13846 11746 13847
rect 20118 18494 20146 18522
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 12278 13846 12306 13874
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 13678 13593 13706 13594
rect 13678 13567 13679 13593
rect 13679 13567 13705 13593
rect 13705 13567 13706 13593
rect 13678 13566 13706 13567
rect 12278 13454 12306 13482
rect 10990 12670 11018 12698
rect 11046 12614 11074 12642
rect 11158 12809 11186 12810
rect 11158 12783 11159 12809
rect 11159 12783 11185 12809
rect 11185 12783 11186 12809
rect 11158 12782 11186 12783
rect 11158 12670 11186 12698
rect 10654 11830 10682 11858
rect 10710 11913 10738 11914
rect 10710 11887 10711 11913
rect 10711 11887 10737 11913
rect 10737 11887 10738 11913
rect 10710 11886 10738 11887
rect 10598 11494 10626 11522
rect 10542 11326 10570 11354
rect 10374 11270 10402 11298
rect 10206 11046 10234 11074
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 9030 10065 9058 10066
rect 9030 10039 9031 10065
rect 9031 10039 9057 10065
rect 9057 10039 9058 10065
rect 9030 10038 9058 10039
rect 9254 10038 9282 10066
rect 8750 9953 8778 9954
rect 8750 9927 8751 9953
rect 8751 9927 8777 9953
rect 8777 9927 8778 9953
rect 8750 9926 8778 9927
rect 9142 9926 9170 9954
rect 8582 9870 8610 9898
rect 8806 9897 8834 9898
rect 8806 9871 8807 9897
rect 8807 9871 8833 9897
rect 8833 9871 8834 9897
rect 8806 9870 8834 9871
rect 8638 9702 8666 9730
rect 7350 9169 7378 9170
rect 7350 9143 7351 9169
rect 7351 9143 7377 9169
rect 7377 9143 7378 9169
rect 7350 9142 7378 9143
rect 7854 9086 7882 9114
rect 8078 9561 8106 9562
rect 8078 9535 8079 9561
rect 8079 9535 8105 9561
rect 8105 9535 8106 9561
rect 8078 9534 8106 9535
rect 8470 9534 8498 9562
rect 8022 9310 8050 9338
rect 8190 9086 8218 9114
rect 8022 8945 8050 8946
rect 8022 8919 8023 8945
rect 8023 8919 8049 8945
rect 8049 8919 8050 8945
rect 8022 8918 8050 8919
rect 9030 9198 9058 9226
rect 7966 8694 7994 8722
rect 5670 8078 5698 8106
rect 6734 8105 6762 8106
rect 6734 8079 6735 8105
rect 6735 8079 6761 8105
rect 6761 8079 6762 8105
rect 6734 8078 6762 8079
rect 8414 8721 8442 8722
rect 8414 8695 8415 8721
rect 8415 8695 8441 8721
rect 8441 8695 8442 8721
rect 8414 8694 8442 8695
rect 8862 8414 8890 8442
rect 7630 7630 7658 7658
rect 8022 7630 8050 7658
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 10038 10766 10066 10794
rect 9758 10401 9786 10402
rect 9758 10375 9759 10401
rect 9759 10375 9785 10401
rect 9785 10375 9786 10401
rect 9758 10374 9786 10375
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9702 10038 9730 10066
rect 9646 10009 9674 10010
rect 9646 9983 9647 10009
rect 9647 9983 9673 10009
rect 9673 9983 9674 10009
rect 9646 9982 9674 9983
rect 9478 9926 9506 9954
rect 9478 9814 9506 9842
rect 9478 9590 9506 9618
rect 9590 9534 9618 9562
rect 9310 9505 9338 9506
rect 9310 9479 9311 9505
rect 9311 9479 9337 9505
rect 9337 9479 9338 9505
rect 9310 9478 9338 9479
rect 9870 9590 9898 9618
rect 9926 10038 9954 10066
rect 10150 10065 10178 10066
rect 10150 10039 10151 10065
rect 10151 10039 10177 10065
rect 10177 10039 10178 10065
rect 10150 10038 10178 10039
rect 9982 9982 10010 10010
rect 10094 9814 10122 9842
rect 9926 9534 9954 9562
rect 10206 9590 10234 9618
rect 9870 9505 9898 9506
rect 9870 9479 9871 9505
rect 9871 9479 9897 9505
rect 9897 9479 9898 9505
rect 9870 9478 9898 9479
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9702 9337 9730 9338
rect 9702 9311 9703 9337
rect 9703 9311 9729 9337
rect 9729 9311 9730 9337
rect 9702 9310 9730 9311
rect 10318 9310 10346 9338
rect 10094 9225 10122 9226
rect 10094 9199 10095 9225
rect 10095 9199 10121 9225
rect 10121 9199 10122 9225
rect 10094 9198 10122 9199
rect 10374 9254 10402 9282
rect 10430 9198 10458 9226
rect 10598 11046 10626 11074
rect 10934 11942 10962 11970
rect 10822 11830 10850 11858
rect 10766 11774 10794 11802
rect 10766 11102 10794 11130
rect 10822 11382 10850 11410
rect 10710 10878 10738 10906
rect 10654 10401 10682 10402
rect 10654 10375 10655 10401
rect 10655 10375 10681 10401
rect 10681 10375 10682 10401
rect 10654 10374 10682 10375
rect 11102 11214 11130 11242
rect 11158 11438 11186 11466
rect 11326 12558 11354 12586
rect 11494 13118 11522 13146
rect 13230 13257 13258 13258
rect 13230 13231 13231 13257
rect 13231 13231 13257 13257
rect 13257 13231 13258 13257
rect 13230 13230 13258 13231
rect 18830 13537 18858 13538
rect 18830 13511 18831 13537
rect 18831 13511 18857 13537
rect 18857 13511 18858 13537
rect 18830 13510 18858 13511
rect 13678 13230 13706 13258
rect 13902 13454 13930 13482
rect 12390 12558 12418 12586
rect 11718 12054 11746 12082
rect 12278 12054 12306 12082
rect 11438 11942 11466 11970
rect 11606 11886 11634 11914
rect 11494 11774 11522 11802
rect 12950 12697 12978 12698
rect 12950 12671 12951 12697
rect 12951 12671 12977 12697
rect 12977 12671 12978 12697
rect 12950 12670 12978 12671
rect 12838 12446 12866 12474
rect 12670 12361 12698 12362
rect 12670 12335 12671 12361
rect 12671 12335 12697 12361
rect 12697 12335 12698 12361
rect 12670 12334 12698 12335
rect 12446 11913 12474 11914
rect 12446 11887 12447 11913
rect 12447 11887 12473 11913
rect 12473 11887 12474 11913
rect 12446 11886 12474 11887
rect 11326 11662 11354 11690
rect 12054 11689 12082 11690
rect 12054 11663 12055 11689
rect 12055 11663 12081 11689
rect 12081 11663 12082 11689
rect 12054 11662 12082 11663
rect 11270 11382 11298 11410
rect 11214 11158 11242 11186
rect 11102 10990 11130 11018
rect 10934 10766 10962 10794
rect 11158 10878 11186 10906
rect 11158 10262 11186 10290
rect 11494 11494 11522 11522
rect 11662 11438 11690 11466
rect 11606 11382 11634 11410
rect 11774 11326 11802 11354
rect 11718 11270 11746 11298
rect 11550 11214 11578 11242
rect 11438 11073 11466 11074
rect 11438 11047 11439 11073
rect 11439 11047 11465 11073
rect 11465 11047 11466 11073
rect 11438 11046 11466 11047
rect 11494 10318 11522 10346
rect 10766 9926 10794 9954
rect 10654 9870 10682 9898
rect 11102 9926 11130 9954
rect 10990 9646 11018 9674
rect 11046 9702 11074 9730
rect 10766 9590 10794 9618
rect 10822 9561 10850 9562
rect 10822 9535 10823 9561
rect 10823 9535 10849 9561
rect 10849 9535 10850 9561
rect 10822 9534 10850 9535
rect 10710 9478 10738 9506
rect 9646 9169 9674 9170
rect 9646 9143 9647 9169
rect 9647 9143 9673 9169
rect 9673 9143 9674 9169
rect 9646 9142 9674 9143
rect 10766 9310 10794 9338
rect 11494 9870 11522 9898
rect 11046 9478 11074 9506
rect 10822 9254 10850 9282
rect 10878 9198 10906 9226
rect 10990 9198 11018 9226
rect 11158 9505 11186 9506
rect 11158 9479 11159 9505
rect 11159 9479 11185 9505
rect 11185 9479 11186 9505
rect 11158 9478 11186 9479
rect 11270 8918 11298 8946
rect 11102 8806 11130 8834
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 10598 8638 10626 8666
rect 9310 8441 9338 8442
rect 9310 8415 9311 8441
rect 9311 8415 9337 8441
rect 9337 8415 9338 8441
rect 9310 8414 9338 8415
rect 10374 8414 10402 8442
rect 9198 7910 9226 7938
rect 10318 8161 10346 8162
rect 10318 8135 10319 8161
rect 10319 8135 10345 8161
rect 10345 8135 10346 8161
rect 10318 8134 10346 8135
rect 10542 8441 10570 8442
rect 10542 8415 10543 8441
rect 10543 8415 10569 8441
rect 10569 8415 10570 8441
rect 10542 8414 10570 8415
rect 10486 8134 10514 8162
rect 10038 7937 10066 7938
rect 10038 7911 10039 7937
rect 10039 7911 10065 7937
rect 10065 7911 10066 7937
rect 10038 7910 10066 7911
rect 10318 7937 10346 7938
rect 10318 7911 10319 7937
rect 10319 7911 10345 7937
rect 10345 7911 10346 7937
rect 10318 7910 10346 7911
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 9702 7713 9730 7714
rect 9702 7687 9703 7713
rect 9703 7687 9729 7713
rect 9729 7687 9730 7713
rect 9702 7686 9730 7687
rect 9254 7630 9282 7658
rect 10206 7574 10234 7602
rect 9366 7126 9394 7154
rect 9142 6817 9170 6818
rect 9142 6791 9143 6817
rect 9143 6791 9169 6817
rect 9169 6791 9170 6817
rect 9142 6790 9170 6791
rect 9646 7153 9674 7154
rect 9646 7127 9647 7153
rect 9647 7127 9673 7153
rect 9673 7127 9674 7153
rect 9646 7126 9674 7127
rect 9814 7126 9842 7154
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 10710 8134 10738 8162
rect 10654 7686 10682 7714
rect 10990 8441 11018 8442
rect 10990 8415 10991 8441
rect 10991 8415 11017 8441
rect 11017 8415 11018 8441
rect 10990 8414 11018 8415
rect 10934 8049 10962 8050
rect 10934 8023 10935 8049
rect 10935 8023 10961 8049
rect 10961 8023 10962 8049
rect 10934 8022 10962 8023
rect 11550 9198 11578 9226
rect 11438 8777 11466 8778
rect 11438 8751 11439 8777
rect 11439 8751 11465 8777
rect 11465 8751 11466 8777
rect 11438 8750 11466 8751
rect 11550 8582 11578 8610
rect 11326 8022 11354 8050
rect 11102 7742 11130 7770
rect 11046 7686 11074 7714
rect 11718 11185 11746 11186
rect 11718 11159 11719 11185
rect 11719 11159 11745 11185
rect 11745 11159 11746 11185
rect 11718 11158 11746 11159
rect 11718 11046 11746 11074
rect 11662 10793 11690 10794
rect 11662 10767 11663 10793
rect 11663 10767 11689 10793
rect 11689 10767 11690 10793
rect 11662 10766 11690 10767
rect 12166 11073 12194 11074
rect 12166 11047 12167 11073
rect 12167 11047 12193 11073
rect 12193 11047 12194 11073
rect 12166 11046 12194 11047
rect 11998 10766 12026 10794
rect 11942 10710 11970 10738
rect 12334 10710 12362 10738
rect 12278 10094 12306 10122
rect 11942 10009 11970 10010
rect 11942 9983 11943 10009
rect 11943 9983 11969 10009
rect 11969 9983 11970 10009
rect 11942 9982 11970 9983
rect 11718 9897 11746 9898
rect 11718 9871 11719 9897
rect 11719 9871 11745 9897
rect 11745 9871 11746 9897
rect 11718 9870 11746 9871
rect 11830 9617 11858 9618
rect 11830 9591 11831 9617
rect 11831 9591 11857 9617
rect 11857 9591 11858 9617
rect 11830 9590 11858 9591
rect 11830 9281 11858 9282
rect 11830 9255 11831 9281
rect 11831 9255 11857 9281
rect 11857 9255 11858 9281
rect 11830 9254 11858 9255
rect 11942 9505 11970 9506
rect 11942 9479 11943 9505
rect 11943 9479 11969 9505
rect 11969 9479 11970 9505
rect 11942 9478 11970 9479
rect 11830 9113 11858 9114
rect 11830 9087 11831 9113
rect 11831 9087 11857 9113
rect 11857 9087 11858 9113
rect 11830 9086 11858 9087
rect 11942 8833 11970 8834
rect 11942 8807 11943 8833
rect 11943 8807 11969 8833
rect 11969 8807 11970 8833
rect 11942 8806 11970 8807
rect 12054 8777 12082 8778
rect 12054 8751 12055 8777
rect 12055 8751 12081 8777
rect 12081 8751 12082 8777
rect 12054 8750 12082 8751
rect 11942 8638 11970 8666
rect 12278 9617 12306 9618
rect 12278 9591 12279 9617
rect 12279 9591 12305 9617
rect 12305 9591 12306 9617
rect 12278 9590 12306 9591
rect 13286 12614 13314 12642
rect 13062 12054 13090 12082
rect 12670 11662 12698 11690
rect 13342 12446 13370 12474
rect 18830 13145 18858 13146
rect 18830 13119 18831 13145
rect 18831 13119 18857 13145
rect 18857 13119 18858 13145
rect 18830 13118 18858 13119
rect 20006 13118 20034 13146
rect 15358 13089 15386 13090
rect 15358 13063 15359 13089
rect 15359 13063 15385 13089
rect 15385 13063 15386 13089
rect 15358 13062 15386 13063
rect 14238 12753 14266 12754
rect 14238 12727 14239 12753
rect 14239 12727 14265 12753
rect 14265 12727 14266 12753
rect 14238 12726 14266 12727
rect 14742 12753 14770 12754
rect 14742 12727 14743 12753
rect 14743 12727 14769 12753
rect 14769 12727 14770 12753
rect 14742 12726 14770 12727
rect 13902 12334 13930 12362
rect 14630 12697 14658 12698
rect 14630 12671 14631 12697
rect 14631 12671 14657 12697
rect 14657 12671 14658 12697
rect 14630 12670 14658 12671
rect 15358 12670 15386 12698
rect 13958 12446 13986 12474
rect 13286 11913 13314 11914
rect 13286 11887 13287 11913
rect 13287 11887 13313 11913
rect 13313 11887 13314 11913
rect 13286 11886 13314 11887
rect 14070 12222 14098 12250
rect 12726 11270 12754 11298
rect 12390 10374 12418 10402
rect 12558 10345 12586 10346
rect 12558 10319 12559 10345
rect 12559 10319 12585 10345
rect 12585 10319 12586 10345
rect 12558 10318 12586 10319
rect 12670 10094 12698 10122
rect 13006 11577 13034 11578
rect 13006 11551 13007 11577
rect 13007 11551 13033 11577
rect 13033 11551 13034 11577
rect 13006 11550 13034 11551
rect 13174 11577 13202 11578
rect 13174 11551 13175 11577
rect 13175 11551 13201 11577
rect 13201 11551 13202 11577
rect 13174 11550 13202 11551
rect 12950 11270 12978 11298
rect 13118 11297 13146 11298
rect 13118 11271 13119 11297
rect 13119 11271 13145 11297
rect 13145 11271 13146 11297
rect 13118 11270 13146 11271
rect 14574 12614 14602 12642
rect 14294 12361 14322 12362
rect 14294 12335 14295 12361
rect 14295 12335 14321 12361
rect 14321 12335 14322 12361
rect 14294 12334 14322 12335
rect 14182 12278 14210 12306
rect 14070 11606 14098 11634
rect 13566 11270 13594 11298
rect 12894 11102 12922 11130
rect 12782 11046 12810 11074
rect 12782 10793 12810 10794
rect 12782 10767 12783 10793
rect 12783 10767 12809 10793
rect 12809 10767 12810 10793
rect 12782 10766 12810 10767
rect 12950 10374 12978 10402
rect 13342 10990 13370 11018
rect 12894 9982 12922 10010
rect 12670 9702 12698 9730
rect 12334 9478 12362 9506
rect 12558 9534 12586 9562
rect 12502 9254 12530 9282
rect 12614 9366 12642 9394
rect 12670 9337 12698 9338
rect 12670 9311 12671 9337
rect 12671 9311 12697 9337
rect 12697 9311 12698 9337
rect 12670 9310 12698 9311
rect 12726 9646 12754 9674
rect 12222 8833 12250 8834
rect 12222 8807 12223 8833
rect 12223 8807 12249 8833
rect 12249 8807 12250 8833
rect 12222 8806 12250 8807
rect 12166 8721 12194 8722
rect 12166 8695 12167 8721
rect 12167 8695 12193 8721
rect 12193 8695 12194 8721
rect 12166 8694 12194 8695
rect 12334 8497 12362 8498
rect 12334 8471 12335 8497
rect 12335 8471 12361 8497
rect 12361 8471 12362 8497
rect 12334 8470 12362 8471
rect 12670 8441 12698 8442
rect 12670 8415 12671 8441
rect 12671 8415 12697 8441
rect 12697 8415 12698 8441
rect 12670 8414 12698 8415
rect 13174 10934 13202 10962
rect 13118 10318 13146 10346
rect 12950 9505 12978 9506
rect 12950 9479 12951 9505
rect 12951 9479 12977 9505
rect 12977 9479 12978 9505
rect 12950 9478 12978 9479
rect 12894 9422 12922 9450
rect 13006 9366 13034 9394
rect 13062 9281 13090 9282
rect 13062 9255 13063 9281
rect 13063 9255 13089 9281
rect 13089 9255 13090 9281
rect 13062 9254 13090 9255
rect 13174 9225 13202 9226
rect 13174 9199 13175 9225
rect 13175 9199 13201 9225
rect 13201 9199 13202 9225
rect 13174 9198 13202 9199
rect 13342 10793 13370 10794
rect 13342 10767 13343 10793
rect 13343 10767 13369 10793
rect 13369 10767 13370 10793
rect 13342 10766 13370 10767
rect 13846 11185 13874 11186
rect 13846 11159 13847 11185
rect 13847 11159 13873 11185
rect 13873 11159 13874 11185
rect 13846 11158 13874 11159
rect 13622 10822 13650 10850
rect 13678 10793 13706 10794
rect 13678 10767 13679 10793
rect 13679 10767 13705 10793
rect 13705 10767 13706 10793
rect 13678 10766 13706 10767
rect 13510 10710 13538 10738
rect 13566 10345 13594 10346
rect 13566 10319 13567 10345
rect 13567 10319 13593 10345
rect 13593 10319 13594 10345
rect 13566 10318 13594 10319
rect 14294 11969 14322 11970
rect 14294 11943 14295 11969
rect 14295 11943 14321 11969
rect 14321 11943 14322 11969
rect 14294 11942 14322 11943
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 19950 12782 19978 12810
rect 20006 12446 20034 12474
rect 18830 12390 18858 12418
rect 15582 12334 15610 12362
rect 15918 12334 15946 12362
rect 14630 12305 14658 12306
rect 14630 12279 14631 12305
rect 14631 12279 14657 12305
rect 14657 12279 14658 12305
rect 14630 12278 14658 12279
rect 15694 12305 15722 12306
rect 15694 12279 15695 12305
rect 15695 12279 15721 12305
rect 15721 12279 15722 12305
rect 15694 12278 15722 12279
rect 14742 11969 14770 11970
rect 14742 11943 14743 11969
rect 14743 11943 14769 11969
rect 14769 11943 14770 11969
rect 14742 11942 14770 11943
rect 14630 11913 14658 11914
rect 14630 11887 14631 11913
rect 14631 11887 14657 11913
rect 14657 11887 14658 11913
rect 14630 11886 14658 11887
rect 15694 11886 15722 11914
rect 14182 11158 14210 11186
rect 14126 10934 14154 10962
rect 14406 10849 14434 10850
rect 14406 10823 14407 10849
rect 14407 10823 14433 10849
rect 14433 10823 14434 10849
rect 14406 10822 14434 10823
rect 13286 10038 13314 10066
rect 13846 10038 13874 10066
rect 13454 9478 13482 9506
rect 13790 9422 13818 9450
rect 13566 9366 13594 9394
rect 13342 9310 13370 9338
rect 13510 9198 13538 9226
rect 13006 8833 13034 8834
rect 13006 8807 13007 8833
rect 13007 8807 13033 8833
rect 13033 8807 13034 8833
rect 13006 8806 13034 8807
rect 13286 8833 13314 8834
rect 13286 8807 13287 8833
rect 13287 8807 13313 8833
rect 13313 8807 13314 8833
rect 13286 8806 13314 8807
rect 13734 9198 13762 9226
rect 15470 10766 15498 10794
rect 18830 12222 18858 12250
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 20006 11774 20034 11802
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 20006 11102 20034 11130
rect 18830 10766 18858 10794
rect 15414 10065 15442 10066
rect 15414 10039 15415 10065
rect 15415 10039 15441 10065
rect 15441 10039 15442 10065
rect 15414 10038 15442 10039
rect 15470 9646 15498 9674
rect 14126 9561 14154 9562
rect 14126 9535 14127 9561
rect 14127 9535 14153 9561
rect 14153 9535 14154 9561
rect 14126 9534 14154 9535
rect 13678 8918 13706 8946
rect 12726 8134 12754 8162
rect 11550 7769 11578 7770
rect 11550 7743 11551 7769
rect 11551 7743 11577 7769
rect 11577 7743 11578 7769
rect 11550 7742 11578 7743
rect 13006 8694 13034 8722
rect 12222 7742 12250 7770
rect 11382 7713 11410 7714
rect 11382 7687 11383 7713
rect 11383 7687 11409 7713
rect 11409 7687 11410 7713
rect 11382 7686 11410 7687
rect 10822 7630 10850 7658
rect 9422 6790 9450 6818
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 854 2449 882 2450
rect 854 2423 855 2449
rect 855 2423 881 2449
rect 881 2423 882 2449
rect 854 2422 882 2423
rect 10710 6790 10738 6818
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 11158 7657 11186 7658
rect 11158 7631 11159 7657
rect 11159 7631 11185 7657
rect 11185 7631 11186 7657
rect 11158 7630 11186 7631
rect 10990 7601 11018 7602
rect 10990 7575 10991 7601
rect 10991 7575 11017 7601
rect 11017 7575 11018 7601
rect 10990 7574 11018 7575
rect 12950 8582 12978 8610
rect 12838 7937 12866 7938
rect 12838 7911 12839 7937
rect 12839 7911 12865 7937
rect 12865 7911 12866 7937
rect 12838 7910 12866 7911
rect 12670 7769 12698 7770
rect 12670 7743 12671 7769
rect 12671 7743 12697 7769
rect 12697 7743 12698 7769
rect 12670 7742 12698 7743
rect 13510 8470 13538 8498
rect 13118 8049 13146 8050
rect 13118 8023 13119 8049
rect 13119 8023 13145 8049
rect 13145 8023 13146 8049
rect 13118 8022 13146 8023
rect 14350 9225 14378 9226
rect 14350 9199 14351 9225
rect 14351 9199 14377 9225
rect 14377 9199 14378 9225
rect 14350 9198 14378 9199
rect 14966 9561 14994 9562
rect 14966 9535 14967 9561
rect 14967 9535 14993 9561
rect 14993 9535 14994 9561
rect 14966 9534 14994 9535
rect 14630 9142 14658 9170
rect 14014 8414 14042 8442
rect 14070 8806 14098 8834
rect 14910 9086 14938 9114
rect 14854 8945 14882 8946
rect 14854 8919 14855 8945
rect 14855 8919 14881 8945
rect 14881 8919 14882 8945
rect 14854 8918 14882 8919
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 16030 9673 16058 9674
rect 16030 9647 16031 9673
rect 16031 9647 16057 9673
rect 16057 9647 16058 9673
rect 16030 9646 16058 9647
rect 20006 10094 20034 10122
rect 18830 9646 18858 9674
rect 18830 9225 18858 9226
rect 18830 9199 18831 9225
rect 18831 9199 18857 9225
rect 18857 9199 18858 9225
rect 18830 9198 18858 9199
rect 15638 9169 15666 9170
rect 15638 9143 15639 9169
rect 15639 9143 15665 9169
rect 15665 9143 15666 9169
rect 15638 9142 15666 9143
rect 15414 9086 15442 9114
rect 20006 9113 20034 9114
rect 20006 9087 20007 9113
rect 20007 9087 20033 9113
rect 20033 9087 20034 9113
rect 20006 9086 20034 9087
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 20006 8750 20034 8778
rect 14294 8441 14322 8442
rect 14294 8415 14295 8441
rect 14295 8415 14321 8441
rect 14321 8415 14322 8441
rect 14294 8414 14322 8415
rect 13510 7993 13538 7994
rect 13510 7967 13511 7993
rect 13511 7967 13537 7993
rect 13537 7967 13538 7993
rect 13510 7966 13538 7967
rect 13006 7742 13034 7770
rect 12614 7518 12642 7546
rect 11494 7182 11522 7210
rect 12390 7182 12418 7210
rect 10990 7153 11018 7154
rect 10990 7127 10991 7153
rect 10991 7127 11017 7153
rect 11017 7127 11018 7153
rect 10990 7126 11018 7127
rect 11830 7126 11858 7154
rect 11270 6817 11298 6818
rect 11270 6791 11271 6817
rect 11271 6791 11297 6817
rect 11297 6791 11298 6817
rect 11270 6790 11298 6791
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 10430 2590 10458 2618
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9422 2030 9450 2058
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9926 2057 9954 2058
rect 9926 2031 9927 2057
rect 9927 2031 9953 2057
rect 9953 2031 9954 2057
rect 9926 2030 9954 2031
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 11158 2617 11186 2618
rect 11158 2591 11159 2617
rect 11159 2591 11185 2617
rect 11185 2591 11186 2617
rect 11158 2590 11186 2591
rect 10766 2030 10794 2058
rect 11382 2057 11410 2058
rect 11382 2031 11383 2057
rect 11383 2031 11409 2057
rect 11409 2031 11410 2057
rect 11382 2030 11410 2031
rect 12054 6790 12082 6818
rect 12558 7209 12586 7210
rect 12558 7183 12559 7209
rect 12559 7183 12585 7209
rect 12585 7183 12586 7209
rect 12558 7182 12586 7183
rect 13174 7518 13202 7546
rect 13230 7126 13258 7154
rect 12614 6790 12642 6818
rect 13566 7518 13594 7546
rect 13734 7153 13762 7154
rect 13734 7127 13735 7153
rect 13735 7127 13761 7153
rect 13761 7127 13762 7153
rect 13734 7126 13762 7127
rect 14070 7126 14098 7154
rect 13734 6790 13762 6818
rect 14630 8414 14658 8442
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 14294 6817 14322 6818
rect 14294 6791 14295 6817
rect 14295 6791 14321 6817
rect 14321 6791 14322 6817
rect 14294 6790 14322 6791
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 20118 2366 20146 2394
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 11433 19110 11438 19138
rect 11466 19110 12782 19138
rect 12810 19110 12815 19138
rect 10593 18886 10598 18914
rect 10626 18886 11774 18914
rect 11802 18886 11807 18914
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 9417 18718 9422 18746
rect 9450 18718 9926 18746
rect 9954 18718 9959 18746
rect 10761 18718 10766 18746
rect 10794 18718 11382 18746
rect 11410 18718 11415 18746
rect 20600 18522 21000 18536
rect 20113 18494 20118 18522
rect 20146 18494 21000 18522
rect 20600 18480 21000 18494
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 8409 18326 8414 18354
rect 8442 18326 9030 18354
rect 9058 18326 9063 18354
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 9641 14014 9646 14042
rect 9674 14014 10150 14042
rect 10178 14014 10183 14042
rect 10649 13846 10654 13874
rect 10682 13846 11046 13874
rect 11074 13846 11079 13874
rect 11433 13846 11438 13874
rect 11466 13846 11718 13874
rect 11746 13846 12278 13874
rect 12306 13846 12311 13874
rect 7345 13790 7350 13818
rect 7378 13790 7910 13818
rect 7938 13790 7943 13818
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 13673 13566 13678 13594
rect 13706 13566 15974 13594
rect 15946 13538 15974 13566
rect 15946 13510 18830 13538
rect 18858 13510 18863 13538
rect 0 13482 400 13496
rect 0 13454 2086 13482
rect 2114 13454 2119 13482
rect 12273 13454 12278 13482
rect 12306 13454 13902 13482
rect 13930 13454 13935 13482
rect 0 13440 400 13454
rect 9137 13398 9142 13426
rect 9170 13398 9310 13426
rect 9338 13398 9646 13426
rect 9674 13398 9679 13426
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 13225 13230 13230 13258
rect 13258 13230 13678 13258
rect 13706 13230 13711 13258
rect 20600 13146 21000 13160
rect 2137 13118 2142 13146
rect 2170 13118 6118 13146
rect 6146 13118 6151 13146
rect 7793 13118 7798 13146
rect 7826 13118 8134 13146
rect 8162 13118 8694 13146
rect 8722 13118 11494 13146
rect 11522 13118 11527 13146
rect 15946 13118 18830 13146
rect 18858 13118 18863 13146
rect 20001 13118 20006 13146
rect 20034 13118 21000 13146
rect 15946 13090 15974 13118
rect 20600 13104 21000 13118
rect 9977 13062 9982 13090
rect 10010 13062 10654 13090
rect 10682 13062 10687 13090
rect 15353 13062 15358 13090
rect 15386 13062 15974 13090
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 8017 12838 8022 12866
rect 8050 12838 8414 12866
rect 8442 12838 8447 12866
rect 0 12810 400 12824
rect 20600 12810 21000 12824
rect 0 12782 966 12810
rect 994 12782 999 12810
rect 9641 12782 9646 12810
rect 9674 12782 11158 12810
rect 11186 12782 11191 12810
rect 19945 12782 19950 12810
rect 19978 12782 21000 12810
rect 0 12768 400 12782
rect 20600 12768 21000 12782
rect 14233 12726 14238 12754
rect 14266 12726 14742 12754
rect 14770 12726 14775 12754
rect 6113 12670 6118 12698
rect 6146 12670 7406 12698
rect 7434 12670 7439 12698
rect 10985 12670 10990 12698
rect 11018 12670 11158 12698
rect 11186 12670 12950 12698
rect 12978 12670 12983 12698
rect 14625 12670 14630 12698
rect 14658 12670 15358 12698
rect 15386 12670 15391 12698
rect 7009 12614 7014 12642
rect 7042 12614 7798 12642
rect 7826 12614 7831 12642
rect 11041 12614 11046 12642
rect 11074 12614 13286 12642
rect 13314 12614 14574 12642
rect 14602 12614 14607 12642
rect 7574 12586 7602 12614
rect 7569 12558 7574 12586
rect 7602 12558 7607 12586
rect 11321 12558 11326 12586
rect 11354 12558 12390 12586
rect 12418 12558 12423 12586
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 20600 12474 21000 12488
rect 7625 12446 7630 12474
rect 7658 12446 8246 12474
rect 8274 12446 8694 12474
rect 8722 12446 8727 12474
rect 12833 12446 12838 12474
rect 12866 12446 13342 12474
rect 13370 12446 13958 12474
rect 13986 12446 13991 12474
rect 20001 12446 20006 12474
rect 20034 12446 21000 12474
rect 20600 12432 21000 12446
rect 18825 12390 18830 12418
rect 18858 12390 18863 12418
rect 12665 12334 12670 12362
rect 12698 12334 13902 12362
rect 13930 12334 14294 12362
rect 14322 12334 15582 12362
rect 15610 12334 15918 12362
rect 15946 12334 15951 12362
rect 18830 12306 18858 12390
rect 14177 12278 14182 12306
rect 14210 12278 14630 12306
rect 14658 12278 14663 12306
rect 15689 12278 15694 12306
rect 15722 12278 18858 12306
rect 14065 12222 14070 12250
rect 14098 12222 18830 12250
rect 18858 12222 18863 12250
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 11713 12054 11718 12082
rect 11746 12054 12278 12082
rect 12306 12054 13062 12082
rect 13090 12054 13095 12082
rect 6729 11942 6734 11970
rect 6762 11942 7294 11970
rect 7322 11942 7327 11970
rect 10929 11942 10934 11970
rect 10962 11942 11438 11970
rect 11466 11942 11471 11970
rect 14289 11942 14294 11970
rect 14322 11942 14742 11970
rect 14770 11942 14775 11970
rect 6897 11886 6902 11914
rect 6930 11886 7406 11914
rect 7434 11886 7439 11914
rect 8857 11886 8862 11914
rect 8890 11886 9198 11914
rect 9226 11886 10710 11914
rect 10738 11886 10743 11914
rect 11601 11886 11606 11914
rect 11634 11886 12446 11914
rect 12474 11886 13286 11914
rect 13314 11886 13319 11914
rect 14625 11886 14630 11914
rect 14658 11886 15694 11914
rect 15722 11886 15727 11914
rect 9081 11830 9086 11858
rect 9114 11830 10094 11858
rect 10122 11830 10654 11858
rect 10682 11830 10822 11858
rect 10850 11830 10855 11858
rect 20600 11802 21000 11816
rect 10761 11774 10766 11802
rect 10794 11774 11494 11802
rect 11522 11774 11527 11802
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 20600 11760 21000 11774
rect 7233 11718 7238 11746
rect 7266 11718 7910 11746
rect 7938 11718 7943 11746
rect 7457 11662 7462 11690
rect 7490 11662 8834 11690
rect 11321 11662 11326 11690
rect 11354 11662 12054 11690
rect 12082 11662 12670 11690
rect 12698 11662 12703 11690
rect 8806 11634 8834 11662
rect 8801 11606 8806 11634
rect 8834 11606 9506 11634
rect 9478 11578 9506 11606
rect 13426 11606 14070 11634
rect 14098 11606 14103 11634
rect 13426 11578 13454 11606
rect 2137 11550 2142 11578
rect 2170 11550 5838 11578
rect 5866 11550 5871 11578
rect 7289 11550 7294 11578
rect 7322 11550 7742 11578
rect 7770 11550 8022 11578
rect 8050 11550 8055 11578
rect 8297 11550 8302 11578
rect 8330 11550 8638 11578
rect 8666 11550 8671 11578
rect 8913 11550 8918 11578
rect 8946 11550 9198 11578
rect 9226 11550 9231 11578
rect 9473 11550 9478 11578
rect 9506 11550 13006 11578
rect 13034 11550 13039 11578
rect 13169 11550 13174 11578
rect 13202 11550 13454 11578
rect 5838 11522 5866 11550
rect 5838 11494 7574 11522
rect 7602 11494 7607 11522
rect 7793 11494 7798 11522
rect 7826 11494 9086 11522
rect 9114 11494 9119 11522
rect 9865 11494 9870 11522
rect 9898 11494 10598 11522
rect 10626 11494 11494 11522
rect 11522 11494 11527 11522
rect 0 11466 400 11480
rect 0 11438 966 11466
rect 994 11438 999 11466
rect 11153 11438 11158 11466
rect 11186 11438 11662 11466
rect 11690 11438 11695 11466
rect 0 11424 400 11438
rect 6897 11382 6902 11410
rect 6930 11382 7630 11410
rect 7658 11382 7663 11410
rect 10817 11382 10822 11410
rect 10850 11382 11270 11410
rect 11298 11382 11606 11410
rect 11634 11382 11639 11410
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 7737 11326 7742 11354
rect 7770 11326 10542 11354
rect 10570 11326 11774 11354
rect 11802 11326 11807 11354
rect 10369 11270 10374 11298
rect 10402 11270 11718 11298
rect 11746 11270 12726 11298
rect 12754 11270 12950 11298
rect 12978 11270 12983 11298
rect 13113 11270 13118 11298
rect 13146 11270 13566 11298
rect 13594 11270 13599 11298
rect 961 11214 966 11242
rect 994 11214 999 11242
rect 11097 11214 11102 11242
rect 11130 11214 11550 11242
rect 11578 11214 11583 11242
rect 13426 11214 13874 11242
rect 0 11130 400 11144
rect 966 11130 994 11214
rect 13426 11186 13454 11214
rect 13846 11186 13874 11214
rect 2137 11158 2142 11186
rect 2170 11158 5782 11186
rect 5810 11158 5815 11186
rect 9081 11158 9086 11186
rect 9114 11158 10962 11186
rect 11041 11158 11046 11186
rect 11074 11158 11214 11186
rect 11242 11158 11247 11186
rect 11713 11158 11718 11186
rect 11746 11158 13454 11186
rect 13841 11158 13846 11186
rect 13874 11158 14182 11186
rect 14210 11158 14215 11186
rect 10934 11130 10962 11158
rect 20600 11130 21000 11144
rect 0 11102 994 11130
rect 10206 11102 10766 11130
rect 10794 11102 10799 11130
rect 10934 11102 11746 11130
rect 12889 11102 12894 11130
rect 12922 11102 12927 11130
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 0 11088 400 11102
rect 10206 11074 10234 11102
rect 11718 11074 11746 11102
rect 5777 11046 5782 11074
rect 5810 11046 7462 11074
rect 7490 11046 7495 11074
rect 8297 11046 8302 11074
rect 8330 11046 10206 11074
rect 10234 11046 10239 11074
rect 10593 11046 10598 11074
rect 10626 11046 11438 11074
rect 11466 11046 11471 11074
rect 11713 11046 11718 11074
rect 11746 11046 11751 11074
rect 12161 11046 12166 11074
rect 12194 11046 12782 11074
rect 12810 11046 12815 11074
rect 12894 11018 12922 11102
rect 20600 11088 21000 11102
rect 11097 10990 11102 11018
rect 11130 10990 13342 11018
rect 13370 10990 13375 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 13169 10934 13174 10962
rect 13202 10934 14126 10962
rect 14154 10934 14159 10962
rect 7793 10878 7798 10906
rect 7826 10878 9142 10906
rect 9170 10878 9175 10906
rect 10705 10878 10710 10906
rect 10738 10878 11158 10906
rect 11186 10878 11191 10906
rect 13617 10822 13622 10850
rect 13650 10822 14406 10850
rect 14434 10822 14439 10850
rect 6785 10766 6790 10794
rect 6818 10766 6902 10794
rect 6930 10766 7630 10794
rect 7658 10766 7663 10794
rect 10033 10766 10038 10794
rect 10066 10766 10934 10794
rect 10962 10766 11662 10794
rect 11690 10766 11998 10794
rect 12026 10766 12031 10794
rect 12777 10766 12782 10794
rect 12810 10766 13342 10794
rect 13370 10766 13375 10794
rect 13673 10766 13678 10794
rect 13706 10766 15470 10794
rect 15498 10766 18830 10794
rect 18858 10766 18863 10794
rect 11937 10710 11942 10738
rect 11970 10710 12334 10738
rect 12362 10710 13510 10738
rect 13538 10710 13543 10738
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 2081 10374 2086 10402
rect 2114 10374 9758 10402
rect 9786 10374 10654 10402
rect 10682 10374 10687 10402
rect 11382 10374 12390 10402
rect 12418 10374 12950 10402
rect 12978 10374 12983 10402
rect 11382 10346 11410 10374
rect 7737 10318 7742 10346
rect 7770 10318 8414 10346
rect 8442 10318 11410 10346
rect 11489 10318 11494 10346
rect 11522 10318 12558 10346
rect 12586 10318 12591 10346
rect 13113 10318 13118 10346
rect 13146 10318 13566 10346
rect 13594 10318 13599 10346
rect 6337 10262 6342 10290
rect 6370 10262 6790 10290
rect 6818 10262 6823 10290
rect 7793 10262 7798 10290
rect 7826 10262 7831 10290
rect 8969 10262 8974 10290
rect 9002 10262 11158 10290
rect 11186 10262 11191 10290
rect 7798 10178 7826 10262
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 6841 10150 6846 10178
rect 6874 10150 6879 10178
rect 7289 10150 7294 10178
rect 7322 10150 7826 10178
rect 0 10122 400 10136
rect 0 10094 966 10122
rect 994 10094 999 10122
rect 0 10080 400 10094
rect 6846 10066 6874 10150
rect 20600 10122 21000 10136
rect 12273 10094 12278 10122
rect 12306 10094 12670 10122
rect 12698 10094 12703 10122
rect 20001 10094 20006 10122
rect 20034 10094 21000 10122
rect 20600 10080 21000 10094
rect 6846 10038 7182 10066
rect 7210 10038 7215 10066
rect 9025 10038 9030 10066
rect 9058 10038 9254 10066
rect 9282 10038 9702 10066
rect 9730 10038 9735 10066
rect 9921 10038 9926 10066
rect 9954 10038 10150 10066
rect 10178 10038 13286 10066
rect 13314 10038 13319 10066
rect 13841 10038 13846 10066
rect 13874 10038 15414 10066
rect 15442 10038 15447 10066
rect 9641 9982 9646 10010
rect 9674 9982 9982 10010
rect 10010 9982 10015 10010
rect 11937 9982 11942 10010
rect 11970 9982 12894 10010
rect 12922 9982 12927 10010
rect 2137 9926 2142 9954
rect 2170 9926 5278 9954
rect 5306 9926 6818 9954
rect 8353 9926 8358 9954
rect 8386 9926 8750 9954
rect 8778 9926 9142 9954
rect 9170 9926 9175 9954
rect 9473 9926 9478 9954
rect 9506 9926 10766 9954
rect 10794 9926 11102 9954
rect 11130 9926 11135 9954
rect 6790 9898 6818 9926
rect 6785 9870 6790 9898
rect 6818 9870 6823 9898
rect 8577 9870 8582 9898
rect 8610 9870 8806 9898
rect 8834 9870 10654 9898
rect 10682 9870 10687 9898
rect 11489 9870 11494 9898
rect 11522 9870 11718 9898
rect 11746 9870 11751 9898
rect 9473 9814 9478 9842
rect 9506 9814 10094 9842
rect 10122 9814 10127 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 6883 9702 6902 9730
rect 6930 9702 6935 9730
rect 8633 9702 8638 9730
rect 8666 9702 11046 9730
rect 11074 9702 12670 9730
rect 12698 9702 12703 9730
rect 10985 9646 10990 9674
rect 11018 9646 12726 9674
rect 12754 9646 12759 9674
rect 15465 9646 15470 9674
rect 15498 9646 16030 9674
rect 16058 9646 18830 9674
rect 18858 9646 18863 9674
rect 7569 9590 7574 9618
rect 7602 9590 9478 9618
rect 9506 9590 9511 9618
rect 9865 9590 9870 9618
rect 9898 9590 10206 9618
rect 10234 9590 10239 9618
rect 10761 9590 10766 9618
rect 10794 9590 11830 9618
rect 11858 9590 12278 9618
rect 12306 9590 12311 9618
rect 7177 9534 7182 9562
rect 7210 9534 8078 9562
rect 8106 9534 8470 9562
rect 8498 9534 8503 9562
rect 9585 9534 9590 9562
rect 9618 9534 9926 9562
rect 9954 9534 9959 9562
rect 10817 9534 10822 9562
rect 10850 9534 12558 9562
rect 12586 9534 12591 9562
rect 14121 9534 14126 9562
rect 14154 9534 14966 9562
rect 14994 9534 14999 9562
rect 9305 9478 9310 9506
rect 9338 9478 9870 9506
rect 9898 9478 10710 9506
rect 10738 9478 10743 9506
rect 11027 9478 11046 9506
rect 11074 9478 11079 9506
rect 11153 9478 11158 9506
rect 11186 9478 11942 9506
rect 11970 9478 12334 9506
rect 12362 9478 12367 9506
rect 12945 9478 12950 9506
rect 12978 9478 13454 9506
rect 13482 9478 13487 9506
rect 11046 9450 11074 9478
rect 11046 9422 12894 9450
rect 12922 9422 13790 9450
rect 13818 9422 13823 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 12609 9366 12614 9394
rect 12642 9366 13006 9394
rect 13034 9366 13566 9394
rect 13594 9366 13599 9394
rect 7289 9310 7294 9338
rect 7322 9310 7686 9338
rect 7714 9310 8022 9338
rect 8050 9310 8055 9338
rect 9697 9310 9702 9338
rect 9730 9310 10318 9338
rect 10346 9310 10766 9338
rect 10794 9310 10799 9338
rect 12665 9310 12670 9338
rect 12698 9310 13342 9338
rect 13370 9310 13375 9338
rect 10369 9254 10374 9282
rect 10402 9254 10822 9282
rect 10850 9254 10855 9282
rect 11825 9254 11830 9282
rect 11858 9254 12502 9282
rect 12530 9254 13062 9282
rect 13090 9254 13095 9282
rect 7401 9198 7406 9226
rect 7434 9198 7574 9226
rect 9025 9198 9030 9226
rect 9058 9198 10094 9226
rect 10122 9198 10127 9226
rect 10425 9198 10430 9226
rect 10458 9198 10878 9226
rect 10906 9198 10911 9226
rect 10985 9198 10990 9226
rect 11018 9198 11550 9226
rect 11578 9198 11583 9226
rect 13169 9198 13174 9226
rect 13202 9198 13510 9226
rect 13538 9198 13543 9226
rect 13729 9198 13734 9226
rect 13762 9198 14350 9226
rect 14378 9198 14383 9226
rect 15946 9198 18830 9226
rect 18858 9198 18863 9226
rect 7546 9170 7574 9198
rect 6729 9142 6734 9170
rect 6762 9142 7350 9170
rect 7378 9142 7383 9170
rect 7546 9142 9646 9170
rect 9674 9142 9679 9170
rect 14625 9142 14630 9170
rect 14658 9142 15638 9170
rect 15666 9142 15671 9170
rect 15946 9114 15974 9198
rect 20600 9114 21000 9128
rect 7849 9086 7854 9114
rect 7882 9086 8190 9114
rect 8218 9086 11830 9114
rect 11858 9086 11863 9114
rect 14905 9086 14910 9114
rect 14938 9086 15414 9114
rect 15442 9086 15974 9114
rect 20001 9086 20006 9114
rect 20034 9086 21000 9114
rect 20600 9072 21000 9086
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 8017 8918 8022 8946
rect 8050 8918 11270 8946
rect 11298 8918 11303 8946
rect 13673 8918 13678 8946
rect 13706 8918 14854 8946
rect 14882 8918 14887 8946
rect 961 8862 966 8890
rect 994 8862 999 8890
rect 0 8778 400 8792
rect 966 8778 994 8862
rect 2137 8806 2142 8834
rect 2170 8806 5670 8834
rect 5698 8806 5703 8834
rect 11097 8806 11102 8834
rect 11130 8806 11942 8834
rect 11970 8806 11975 8834
rect 12217 8806 12222 8834
rect 12250 8806 13006 8834
rect 13034 8806 13039 8834
rect 13281 8806 13286 8834
rect 13314 8806 14070 8834
rect 14098 8806 18830 8834
rect 18858 8806 18863 8834
rect 20600 8778 21000 8792
rect 0 8750 994 8778
rect 11433 8750 11438 8778
rect 11466 8750 12054 8778
rect 12082 8750 12087 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 0 8736 400 8750
rect 20600 8736 21000 8750
rect 7961 8694 7966 8722
rect 7994 8694 8414 8722
rect 8442 8694 8447 8722
rect 12161 8694 12166 8722
rect 12194 8694 13006 8722
rect 13034 8694 13039 8722
rect 10593 8638 10598 8666
rect 10626 8638 11942 8666
rect 11970 8638 11975 8666
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 11545 8582 11550 8610
rect 11578 8582 12950 8610
rect 12978 8582 12983 8610
rect 12329 8470 12334 8498
rect 12362 8470 13510 8498
rect 13538 8470 13543 8498
rect 8857 8414 8862 8442
rect 8890 8414 9310 8442
rect 9338 8414 9343 8442
rect 10369 8414 10374 8442
rect 10402 8414 10542 8442
rect 10570 8414 10990 8442
rect 11018 8414 11023 8442
rect 12665 8414 12670 8442
rect 12698 8414 14014 8442
rect 14042 8414 14294 8442
rect 14322 8414 14630 8442
rect 14658 8414 14663 8442
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 10313 8134 10318 8162
rect 10346 8134 10486 8162
rect 10514 8134 10710 8162
rect 10738 8134 10743 8162
rect 12721 8134 12726 8162
rect 12754 8134 12759 8162
rect 5665 8078 5670 8106
rect 5698 8078 6734 8106
rect 6762 8078 6767 8106
rect 10929 8022 10934 8050
rect 10962 8022 11326 8050
rect 11354 8022 11359 8050
rect 12726 7938 12754 8134
rect 13113 8022 13118 8050
rect 13146 8022 13454 8050
rect 13426 7994 13454 8022
rect 13426 7966 13510 7994
rect 13538 7966 13543 7994
rect 9193 7910 9198 7938
rect 9226 7910 10038 7938
rect 10066 7910 10071 7938
rect 10313 7910 10318 7938
rect 10346 7910 12838 7938
rect 12866 7910 12871 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 11097 7742 11102 7770
rect 11130 7742 11550 7770
rect 11578 7742 11583 7770
rect 12217 7742 12222 7770
rect 12250 7742 12670 7770
rect 12698 7742 13006 7770
rect 13034 7742 13039 7770
rect 9697 7686 9702 7714
rect 9730 7686 10654 7714
rect 10682 7686 10687 7714
rect 11041 7686 11046 7714
rect 11074 7686 11382 7714
rect 11410 7686 11415 7714
rect 7625 7630 7630 7658
rect 7658 7630 8022 7658
rect 8050 7630 9254 7658
rect 9282 7630 9287 7658
rect 10817 7630 10822 7658
rect 10850 7630 11158 7658
rect 11186 7630 11191 7658
rect 10201 7574 10206 7602
rect 10234 7574 10990 7602
rect 11018 7574 11023 7602
rect 12609 7518 12614 7546
rect 12642 7518 13174 7546
rect 13202 7518 13566 7546
rect 13594 7518 13599 7546
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 11489 7182 11494 7210
rect 11522 7182 12390 7210
rect 12418 7182 12558 7210
rect 12586 7182 12591 7210
rect 9361 7126 9366 7154
rect 9394 7126 9646 7154
rect 9674 7126 9814 7154
rect 9842 7126 10990 7154
rect 11018 7126 11830 7154
rect 11858 7126 11863 7154
rect 13225 7126 13230 7154
rect 13258 7126 13734 7154
rect 13762 7126 14070 7154
rect 14098 7126 14103 7154
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 9137 6790 9142 6818
rect 9170 6790 9422 6818
rect 9450 6790 9455 6818
rect 10705 6790 10710 6818
rect 10738 6790 11270 6818
rect 11298 6790 11303 6818
rect 12049 6790 12054 6818
rect 12082 6790 12614 6818
rect 12642 6790 13734 6818
rect 13762 6790 14294 6818
rect 14322 6790 14327 6818
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 10425 2590 10430 2618
rect 10458 2590 11158 2618
rect 11186 2590 11191 2618
rect 849 2422 854 2450
rect 882 2422 887 2450
rect 0 2394 400 2408
rect 854 2394 882 2422
rect 20600 2394 21000 2408
rect 0 2366 882 2394
rect 20113 2366 20118 2394
rect 20146 2366 21000 2394
rect 0 2352 400 2366
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 20600 2352 21000 2366
rect 9417 2030 9422 2058
rect 9450 2030 9926 2058
rect 9954 2030 9959 2058
rect 10761 2030 10766 2058
rect 10794 2030 11382 2058
rect 11410 2030 11415 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 11046 11158 11074 11186
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 6902 10766 6930 10794
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 6902 9702 6930 9730
rect 11046 9478 11074 9506
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 6902 10794 6930 10799
rect 6902 9730 6930 10766
rect 6902 9697 6930 9702
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 9422 10064 10178
rect 11046 11186 11074 11191
rect 11046 9506 11074 11158
rect 11046 9473 11074 9478
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8680 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10024 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10920 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10360 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform -1 0 13832 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13272 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform -1 0 11760 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _120_
timestamp 1698175906
transform -1 0 10304 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform -1 0 9744 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8736 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698175906
transform -1 0 9296 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9072 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform -1 0 7896 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _127_
timestamp 1698175906
transform 1 0 9072 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _128_
timestamp 1698175906
transform -1 0 10080 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_
timestamp 1698175906
transform -1 0 9744 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _130_
timestamp 1698175906
transform -1 0 12880 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform 1 0 13272 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform -1 0 12432 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _133_
timestamp 1698175906
transform -1 0 12376 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _134_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12152 0 -1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7896 0 -1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _136_
timestamp 1698175906
transform -1 0 7000 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _137_
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13496 0 1 7056
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _139_
timestamp 1698175906
transform -1 0 12824 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _140_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _141_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11984 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _142_
timestamp 1698175906
transform -1 0 11144 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _143_
timestamp 1698175906
transform 1 0 10920 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _144_
timestamp 1698175906
transform 1 0 7952 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _145_
timestamp 1698175906
transform 1 0 8288 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _146_
timestamp 1698175906
transform -1 0 8680 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _147_
timestamp 1698175906
transform -1 0 7952 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _148_
timestamp 1698175906
transform -1 0 7840 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _149_
timestamp 1698175906
transform -1 0 8008 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _150_
timestamp 1698175906
transform 1 0 9800 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _151_
timestamp 1698175906
transform -1 0 11592 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _152_
timestamp 1698175906
transform -1 0 12544 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _153_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11256 0 -1 13328
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _154_
timestamp 1698175906
transform -1 0 11200 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _155_
timestamp 1698175906
transform -1 0 13664 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _156_
timestamp 1698175906
transform 1 0 10136 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _157_
timestamp 1698175906
transform -1 0 12432 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _158_
timestamp 1698175906
transform 1 0 12712 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _159_
timestamp 1698175906
transform -1 0 11032 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _160_
timestamp 1698175906
transform 1 0 11424 0 -1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _161_
timestamp 1698175906
transform 1 0 10808 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _162_
timestamp 1698175906
transform -1 0 15008 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _163_
timestamp 1698175906
transform 1 0 10640 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _164_
timestamp 1698175906
transform 1 0 12040 0 1 9408
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _165_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13888 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _166_
timestamp 1698175906
transform 1 0 11200 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _167_
timestamp 1698175906
transform 1 0 12880 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _168_
timestamp 1698175906
transform 1 0 11704 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _169_
timestamp 1698175906
transform 1 0 11032 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _170_
timestamp 1698175906
transform 1 0 10976 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _171_
timestamp 1698175906
transform -1 0 12320 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _172_
timestamp 1698175906
transform -1 0 10472 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _173_
timestamp 1698175906
transform -1 0 10920 0 -1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _174_
timestamp 1698175906
transform -1 0 11144 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _175_
timestamp 1698175906
transform 1 0 9520 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _176_
timestamp 1698175906
transform -1 0 11144 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _177_
timestamp 1698175906
transform 1 0 10024 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _178_
timestamp 1698175906
transform 1 0 9072 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _179_
timestamp 1698175906
transform -1 0 10192 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _180_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9800 0 -1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _181_
timestamp 1698175906
transform -1 0 8960 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _182_
timestamp 1698175906
transform 1 0 12600 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _183_
timestamp 1698175906
transform 1 0 12992 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _184_
timestamp 1698175906
transform 1 0 11928 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _185_
timestamp 1698175906
transform 1 0 13272 0 -1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _186_
timestamp 1698175906
transform 1 0 11312 0 -1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _187_
timestamp 1698175906
transform 1 0 11592 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _188_
timestamp 1698175906
transform 1 0 11480 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _189_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13888 0 1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _190_
timestamp 1698175906
transform -1 0 15568 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _191_
timestamp 1698175906
transform 1 0 13384 0 1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _192_
timestamp 1698175906
transform -1 0 13216 0 1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _193_
timestamp 1698175906
transform 1 0 13216 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _194_
timestamp 1698175906
transform 1 0 13888 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _195_
timestamp 1698175906
transform 1 0 12712 0 -1 11760
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _196_
timestamp 1698175906
transform 1 0 12824 0 1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _197_
timestamp 1698175906
transform 1 0 13216 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _198_
timestamp 1698175906
transform 1 0 12712 0 -1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _199_
timestamp 1698175906
transform -1 0 11424 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _200_
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _201_
timestamp 1698175906
transform -1 0 14336 0 1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _202_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11256 0 -1 12544
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _203_
timestamp 1698175906
transform -1 0 10808 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _204_
timestamp 1698175906
transform -1 0 13384 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _205_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13272 0 1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _206_
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _207_
timestamp 1698175906
transform -1 0 14280 0 1 12544
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _208_
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _209_
timestamp 1698175906
transform 1 0 10864 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _210_
timestamp 1698175906
transform -1 0 7784 0 1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _211_
timestamp 1698175906
transform -1 0 7000 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _212_
timestamp 1698175906
transform -1 0 9240 0 -1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _213_
timestamp 1698175906
transform -1 0 8960 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _214_
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _215_
timestamp 1698175906
transform -1 0 8680 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _216_
timestamp 1698175906
transform -1 0 8848 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _217_
timestamp 1698175906
transform -1 0 7000 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _218_
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _219_
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _220_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7000 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _221_
timestamp 1698175906
transform 1 0 8064 0 -1 14112
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _222_
timestamp 1698175906
transform 1 0 7840 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _223_
timestamp 1698175906
transform -1 0 8064 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _224_
timestamp 1698175906
transform -1 0 7840 0 1 12544
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _225_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7728 0 1 11760
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8008 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform -1 0 7392 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 11928 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 7504 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 6832 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 10192 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform -1 0 11424 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 13888 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform 1 0 9240 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 7896 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698175906
transform 1 0 13944 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _240_
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _241_
timestamp 1698175906
transform 1 0 14168 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _242_
timestamp 1698175906
transform 1 0 9520 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _243_
timestamp 1698175906
transform 1 0 12152 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _244_
timestamp 1698175906
transform 1 0 13832 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _245_
timestamp 1698175906
transform 1 0 9744 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _246_
timestamp 1698175906
transform -1 0 7336 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _247_
timestamp 1698175906
transform 1 0 7560 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _248_
timestamp 1698175906
transform -1 0 6832 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _249_
timestamp 1698175906
transform -1 0 7224 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _250_
timestamp 1698175906
transform 1 0 6888 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _251_
timestamp 1698175906
transform -1 0 7672 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _255_
timestamp 1698175906
transform 1 0 11368 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__160__B2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11480 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 9744 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 8008 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 14280 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform -1 0 13776 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 9240 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 9016 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform -1 0 10192 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 12040 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 15624 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 14280 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform 1 0 10976 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 9632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform 1 0 15680 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform 1 0 14616 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__CLK
timestamp 1698175906
transform 1 0 13832 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__CLK
timestamp 1698175906
transform 1 0 15904 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__CLK
timestamp 1698175906
transform 1 0 11144 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__CLK
timestamp 1698175906
transform 1 0 13888 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__CLK
timestamp 1698175906
transform 1 0 15568 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__CLK
timestamp 1698175906
transform 1 0 11816 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__CLK
timestamp 1698175906
transform 1 0 7448 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__CLK
timestamp 1698175906
transform 1 0 9296 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__CLK
timestamp 1698175906
transform 1 0 7112 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__CLK
timestamp 1698175906
transform 1 0 7336 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__CLK
timestamp 1698175906
transform 1 0 9128 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__CLK
timestamp 1698175906
transform 1 0 7784 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 9800 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output23_I
timestamp 1698175906
transform -1 0 10640 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 11592 0 -1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698175906
transform 1 0 9072 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_154
timestamp 1698175906
transform 1 0 9296 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 12264 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 16128 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_6 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1008 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_22
timestamp 1698175906
transform 1 0 1904 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_30
timestamp 1698175906
transform 1 0 2352 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_203
timestamp 1698175906
transform 1 0 12040 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_235
timestamp 1698175906
transform 1 0 13832 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_243
timestamp 1698175906
transform 1 0 14280 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_333
timestamp 1698175906
transform 1 0 19320 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_341
timestamp 1698175906
transform 1 0 19768 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 10248 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_193
timestamp 1698175906
transform 1 0 11480 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_230
timestamp 1698175906
transform 1 0 13552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_234
timestamp 1698175906
transform 1 0 13776 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_242
timestamp 1698175906
transform 1 0 14224 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698175906
transform 1 0 14336 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_154
timestamp 1698175906
transform 1 0 9296 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_197
timestamp 1698175906
transform 1 0 11704 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_201
timestamp 1698175906
transform 1 0 11928 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 12376 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_241
timestamp 1698175906
transform 1 0 14168 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_245
timestamp 1698175906
transform 1 0 14392 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_277
timestamp 1698175906
transform 1 0 16184 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698175906
transform 1 0 16296 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_123
timestamp 1698175906
transform 1 0 7560 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_127
timestamp 1698175906
transform 1 0 7784 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_158
timestamp 1698175906
transform 1 0 9520 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_162
timestamp 1698175906
transform 1 0 9744 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_170
timestamp 1698175906
transform 1 0 10192 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 10416 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_182
timestamp 1698175906
transform 1 0 10864 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_186
timestamp 1698175906
transform 1 0 11088 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_202
timestamp 1698175906
transform 1 0 11984 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_210
timestamp 1698175906
transform 1 0 12432 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_235
timestamp 1698175906
transform 1 0 13832 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698175906
transform 1 0 14280 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 8288 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_148
timestamp 1698175906
transform 1 0 8960 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_152
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_195
timestamp 1698175906
transform 1 0 11592 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_203
timestamp 1698175906
transform 1 0 12040 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698175906
transform 1 0 12264 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 12376 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_216
timestamp 1698175906
transform 1 0 12768 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_225
timestamp 1698175906
transform 1 0 13272 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_257
timestamp 1698175906
transform 1 0 15064 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_273
timestamp 1698175906
transform 1 0 15960 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698175906
transform 1 0 16184 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 16296 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_111
timestamp 1698175906
transform 1 0 6888 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_119
timestamp 1698175906
transform 1 0 7336 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_121
timestamp 1698175906
transform 1 0 7448 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_151
timestamp 1698175906
transform 1 0 9128 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_155
timestamp 1698175906
transform 1 0 9352 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_163
timestamp 1698175906
transform 1 0 9800 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_187
timestamp 1698175906
transform 1 0 11144 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_195
timestamp 1698175906
transform 1 0 11592 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_199
timestamp 1698175906
transform 1 0 11816 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_210
timestamp 1698175906
transform 1 0 12432 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_214
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_231
timestamp 1698175906
transform 1 0 13608 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_239
timestamp 1698175906
transform 1 0 14056 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 14280 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_117
timestamp 1698175906
transform 1 0 7224 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_121
timestamp 1698175906
transform 1 0 7448 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698175906
transform 1 0 8344 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 8456 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_150
timestamp 1698175906
transform 1 0 9072 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_152
timestamp 1698175906
transform 1 0 9184 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_163
timestamp 1698175906
transform 1 0 9800 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_171
timestamp 1698175906
transform 1 0 10248 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_173
timestamp 1698175906
transform 1 0 10360 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_189
timestamp 1698175906
transform 1 0 11256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_197
timestamp 1698175906
transform 1 0 11704 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_201
timestamp 1698175906
transform 1 0 11928 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_203
timestamp 1698175906
transform 1 0 12040 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_241
timestamp 1698175906
transform 1 0 14168 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_245
timestamp 1698175906
transform 1 0 14392 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698175906
transform 1 0 16184 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 16296 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 20048 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 20160 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_123
timestamp 1698175906
transform 1 0 7560 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_127
timestamp 1698175906
transform 1 0 7784 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_129
timestamp 1698175906
transform 1 0 7896 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_142
timestamp 1698175906
transform 1 0 8624 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 10416 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_187
timestamp 1698175906
transform 1 0 11144 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_193
timestamp 1698175906
transform 1 0 11480 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_197
timestamp 1698175906
transform 1 0 11704 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_199
timestamp 1698175906
transform 1 0 11816 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_208
timestamp 1698175906
transform 1 0 12320 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_232
timestamp 1698175906
transform 1 0 13664 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_240
timestamp 1698175906
transform 1 0 14112 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 14336 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_251
timestamp 1698175906
transform 1 0 14728 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_256
timestamp 1698175906
transform 1 0 15008 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_288
timestamp 1698175906
transform 1 0 16800 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_304
timestamp 1698175906
transform 1 0 17696 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_312
timestamp 1698175906
transform 1 0 18144 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698175906
transform 1 0 18256 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_104
timestamp 1698175906
transform 1 0 6496 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_112
timestamp 1698175906
transform 1 0 6944 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_123
timestamp 1698175906
transform 1 0 7560 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_130
timestamp 1698175906
transform 1 0 7952 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698175906
transform 1 0 8400 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_164
timestamp 1698175906
transform 1 0 9856 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_166
timestamp 1698175906
transform 1 0 9968 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_175
timestamp 1698175906
transform 1 0 10472 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_179
timestamp 1698175906
transform 1 0 10696 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_181
timestamp 1698175906
transform 1 0 10808 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_187
timestamp 1698175906
transform 1 0 11144 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_195
timestamp 1698175906
transform 1 0 11592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_202
timestamp 1698175906
transform 1 0 11984 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_225
timestamp 1698175906
transform 1 0 13272 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_265
timestamp 1698175906
transform 1 0 15512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_269
timestamp 1698175906
transform 1 0 15736 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698175906
transform 1 0 16184 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 16296 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 18256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 18704 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_113
timestamp 1698175906
transform 1 0 7000 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_117
timestamp 1698175906
transform 1 0 7224 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_121
timestamp 1698175906
transform 1 0 7448 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_146
timestamp 1698175906
transform 1 0 8848 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_172
timestamp 1698175906
transform 1 0 10304 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698175906
transform 1 0 10416 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_183
timestamp 1698175906
transform 1 0 10920 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_192
timestamp 1698175906
transform 1 0 11424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_196
timestamp 1698175906
transform 1 0 11648 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_234
timestamp 1698175906
transform 1 0 13776 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_242
timestamp 1698175906
transform 1 0 14224 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 14336 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_276
timestamp 1698175906
transform 1 0 16128 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_308
timestamp 1698175906
transform 1 0 17920 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698175906
transform 1 0 18144 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698175906
transform 1 0 18256 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_80
timestamp 1698175906
transform 1 0 5152 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 8456 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_142
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_147
timestamp 1698175906
transform 1 0 8904 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_151
timestamp 1698175906
transform 1 0 9128 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_155
timestamp 1698175906
transform 1 0 9352 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_162
timestamp 1698175906
transform 1 0 9744 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_166
timestamp 1698175906
transform 1 0 9968 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_175
timestamp 1698175906
transform 1 0 10472 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_190
timestamp 1698175906
transform 1 0 11312 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_194
timestamp 1698175906
transform 1 0 11536 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 12376 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_266
timestamp 1698175906
transform 1 0 15568 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_274
timestamp 1698175906
transform 1 0 16016 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 16240 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 20048 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 20160 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698175906
transform 1 0 2240 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698175906
transform 1 0 2464 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_113
timestamp 1698175906
transform 1 0 7000 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_121
timestamp 1698175906
transform 1 0 7448 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_131
timestamp 1698175906
transform 1 0 8008 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_135
timestamp 1698175906
transform 1 0 8232 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_143
timestamp 1698175906
transform 1 0 8680 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_150
timestamp 1698175906
transform 1 0 9072 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_158
timestamp 1698175906
transform 1 0 9520 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_160
timestamp 1698175906
transform 1 0 9632 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_237
timestamp 1698175906
transform 1 0 13944 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 18648 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_88
timestamp 1698175906
transform 1 0 5600 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_119
timestamp 1698175906
transform 1 0 7336 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_129
timestamp 1698175906
transform 1 0 7896 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_137
timestamp 1698175906
transform 1 0 8344 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698175906
transform 1 0 8456 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_144
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_203
timestamp 1698175906
transform 1 0 12040 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_207
timestamp 1698175906
transform 1 0 12264 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 12376 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_214
timestamp 1698175906
transform 1 0 12656 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_235
timestamp 1698175906
transform 1 0 13832 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_266
timestamp 1698175906
transform 1 0 15568 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_270
timestamp 1698175906
transform 1 0 15792 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 16240 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 20048 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 20160 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 2240 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 2464 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_113
timestamp 1698175906
transform 1 0 7000 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_117
timestamp 1698175906
transform 1 0 7224 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_127
timestamp 1698175906
transform 1 0 7784 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_160
timestamp 1698175906
transform 1 0 9632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_164
timestamp 1698175906
transform 1 0 9856 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_166
timestamp 1698175906
transform 1 0 9968 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_173
timestamp 1698175906
transform 1 0 10360 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_177
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_189
timestamp 1698175906
transform 1 0 11256 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_198
timestamp 1698175906
transform 1 0 11760 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_200
timestamp 1698175906
transform 1 0 11872 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_207
timestamp 1698175906
transform 1 0 12264 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_211
timestamp 1698175906
transform 1 0 12488 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_219
timestamp 1698175906
transform 1 0 12936 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_225
timestamp 1698175906
transform 1 0 13272 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_236
timestamp 1698175906
transform 1 0 13888 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 14336 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 2240 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 4032 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 4480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_88
timestamp 1698175906
transform 1 0 5600 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_90
timestamp 1698175906
transform 1 0 5712 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_129
timestamp 1698175906
transform 1 0 7896 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_133
timestamp 1698175906
transform 1 0 8120 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698175906
transform 1 0 8344 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 8456 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_158
timestamp 1698175906
transform 1 0 9520 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_162
timestamp 1698175906
transform 1 0 9744 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_201
timestamp 1698175906
transform 1 0 11928 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_205
timestamp 1698175906
transform 1 0 12152 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_214
timestamp 1698175906
transform 1 0 12656 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_225
timestamp 1698175906
transform 1 0 13272 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_257
timestamp 1698175906
transform 1 0 15064 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698175906
transform 1 0 15960 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 16184 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 16296 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 20048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 20160 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_113
timestamp 1698175906
transform 1 0 7000 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_126
timestamp 1698175906
transform 1 0 7728 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_142
timestamp 1698175906
transform 1 0 8624 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_146
timestamp 1698175906
transform 1 0 8848 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_154
timestamp 1698175906
transform 1 0 9296 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_170
timestamp 1698175906
transform 1 0 10192 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 10416 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_198
timestamp 1698175906
transform 1 0 11760 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_206
timestamp 1698175906
transform 1 0 12208 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_212
timestamp 1698175906
transform 1 0 12544 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_216
timestamp 1698175906
transform 1 0 12768 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_229
timestamp 1698175906
transform 1 0 13496 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_233
timestamp 1698175906
transform 1 0 13720 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 14336 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_252
timestamp 1698175906
transform 1 0 14784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_284
timestamp 1698175906
transform 1 0 16576 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_300
timestamp 1698175906
transform 1 0 17472 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_308
timestamp 1698175906
transform 1 0 17920 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_312
timestamp 1698175906
transform 1 0 18144 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698175906
transform 1 0 18256 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_88
timestamp 1698175906
transform 1 0 5600 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_125
timestamp 1698175906
transform 1 0 7672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_129
timestamp 1698175906
transform 1 0 7896 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_137
timestamp 1698175906
transform 1 0 8344 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 8456 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_153
timestamp 1698175906
transform 1 0 9240 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_169
timestamp 1698175906
transform 1 0 10136 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_177
timestamp 1698175906
transform 1 0 10584 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_195
timestamp 1698175906
transform 1 0 11592 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_203
timestamp 1698175906
transform 1 0 12040 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_207
timestamp 1698175906
transform 1 0 12264 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698175906
transform 1 0 12376 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_270
timestamp 1698175906
transform 1 0 15792 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_274
timestamp 1698175906
transform 1 0 16016 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698175906
transform 1 0 16240 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_115
timestamp 1698175906
transform 1 0 7112 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_119
timestamp 1698175906
transform 1 0 7336 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_128
timestamp 1698175906
transform 1 0 7840 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_136
timestamp 1698175906
transform 1 0 8288 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_143
timestamp 1698175906
transform 1 0 8680 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_181
timestamp 1698175906
transform 1 0 10808 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_185
timestamp 1698175906
transform 1 0 11032 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_189
timestamp 1698175906
transform 1 0 11256 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_205
timestamp 1698175906
transform 1 0 12152 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_213
timestamp 1698175906
transform 1 0 12600 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_215
timestamp 1698175906
transform 1 0 12712 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_225
timestamp 1698175906
transform 1 0 13272 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_233
timestamp 1698175906
transform 1 0 13720 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_235
timestamp 1698175906
transform 1 0 13832 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698175906
transform 1 0 14280 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_252
timestamp 1698175906
transform 1 0 14784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_284
timestamp 1698175906
transform 1 0 16576 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_300
timestamp 1698175906
transform 1 0 17472 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_308
timestamp 1698175906
transform 1 0 17920 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_312
timestamp 1698175906
transform 1 0 18144 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698175906
transform 1 0 18256 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 18648 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 2240 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 4032 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 4480 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_104
timestamp 1698175906
transform 1 0 6496 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_108
timestamp 1698175906
transform 1 0 6720 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_110
timestamp 1698175906
transform 1 0 6832 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_149
timestamp 1698175906
transform 1 0 9016 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_153
timestamp 1698175906
transform 1 0 9240 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_157
timestamp 1698175906
transform 1 0 9464 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_187
timestamp 1698175906
transform 1 0 11144 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_199
timestamp 1698175906
transform 1 0 11816 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698175906
transform 1 0 12264 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 12376 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_212
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_220
timestamp 1698175906
transform 1 0 12992 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_227
timestamp 1698175906
transform 1 0 13384 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_264
timestamp 1698175906
transform 1 0 15456 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_268
timestamp 1698175906
transform 1 0 15680 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 16128 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_152
timestamp 1698175906
transform 1 0 9184 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_156
timestamp 1698175906
transform 1 0 9408 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_172
timestamp 1698175906
transform 1 0 10304 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698175906
transform 1 0 10416 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_181
timestamp 1698175906
transform 1 0 10808 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_183
timestamp 1698175906
transform 1 0 10920 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_188
timestamp 1698175906
transform 1 0 11200 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_204
timestamp 1698175906
transform 1 0 12096 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_234
timestamp 1698175906
transform 1 0 13776 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698175906
transform 1 0 14000 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 14224 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 18648 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_104
timestamp 1698175906
transform 1 0 6496 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_120
timestamp 1698175906
transform 1 0 7392 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_124
timestamp 1698175906
transform 1 0 7616 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_126
timestamp 1698175906
transform 1 0 7728 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698175906
transform 1 0 8456 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_158
timestamp 1698175906
transform 1 0 9520 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_166
timestamp 1698175906
transform 1 0 9968 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_199
timestamp 1698175906
transform 1 0 11816 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698175906
transform 1 0 12264 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 12376 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_165
timestamp 1698175906
transform 1 0 9912 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_173
timestamp 1698175906
transform 1 0 10360 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_150
timestamp 1698175906
transform 1 0 9072 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_154
timestamp 1698175906
transform 1 0 9296 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 16128 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_314
timestamp 1698175906
transform 1 0 18256 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_330
timestamp 1698175906
transform 1 0 19152 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_338
timestamp 1698175906
transform 1 0 19600 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_342
timestamp 1698175906
transform 1 0 19824 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_344
timestamp 1698175906
transform 1 0 19936 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita50_24 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19992 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita50_25
timestamp 1698175906
transform 1 0 19992 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita50_26
timestamp 1698175906
transform -1 0 1008 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18760 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 8456 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 12096 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 10808 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18760 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 10808 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 18760 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 9352 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 8736 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 2240 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 18760 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 2240 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform -1 0 2240 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 2240 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 9352 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 12096 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13440 400 13496 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 20600 18480 21000 18536 0 FreeSans 224 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 20600 10080 21000 10136 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 8400 20600 8456 21000 0 FreeSans 224 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 20600 2352 21000 2408 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 0 8736 400 8792 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 11088 0 11144 400 0 FreeSans 224 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 0 2352 400 2408 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 10752 0 10808 400 0 FreeSans 224 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 20600 12432 21000 12488 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 10752 20600 10808 21000 0 FreeSans 224 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 9408 0 9464 400 0 FreeSans 224 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 9072 20600 9128 21000 0 FreeSans 224 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 10080 400 10136 0 FreeSans 224 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 10416 0 10472 400 0 FreeSans 224 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 20600 9072 21000 9128 0 FreeSans 224 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 11424 20600 11480 21000 0 FreeSans 224 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 11088 400 11144 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 0 11424 400 11480 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 12768 400 12824 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 9408 20600 9464 21000 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 8372 7434 8372 7434 0 _000_
rlabel metal3 14028 10836 14028 10836 0 _001_
rlabel metal3 14560 9548 14560 9548 0 _002_
rlabel metal2 13020 12152 13020 12152 0 _003_
rlabel metal2 14196 12180 14196 12180 0 _004_
rlabel metal2 10668 12964 10668 12964 0 _005_
rlabel metal2 12712 13468 12712 13468 0 _006_
rlabel metal2 14140 12964 14140 12964 0 _007_
rlabel metal3 10612 7588 10612 7588 0 _008_
rlabel metal2 6916 10836 6916 10836 0 _009_
rlabel metal2 8428 12796 8428 12796 0 _010_
rlabel metal2 6356 10164 6356 10164 0 _011_
rlabel metal2 6748 8820 6748 8820 0 _012_
rlabel metal3 7644 13804 7644 13804 0 _013_
rlabel metal2 7196 12068 7196 12068 0 _014_
rlabel metal2 8484 11256 8484 11256 0 _015_
rlabel metal2 6804 11368 6804 11368 0 _016_
rlabel metal3 12460 7756 12460 7756 0 _017_
rlabel metal3 12040 7196 12040 7196 0 _018_
rlabel metal2 7980 8400 7980 8400 0 _019_
rlabel metal3 7812 10220 7812 10220 0 _020_
rlabel metal2 11060 13748 11060 13748 0 _021_
rlabel metal2 10948 11368 10948 11368 0 _022_
rlabel metal2 13748 9240 13748 9240 0 _023_
rlabel metal2 13020 8596 13020 8596 0 _024_
rlabel metal3 10192 7700 10192 7700 0 _025_
rlabel metal2 11172 11312 11172 11312 0 _026_
rlabel metal3 14280 8932 14280 8932 0 _027_
rlabel metal2 13804 9352 13804 9352 0 _028_
rlabel metal2 13580 9296 13580 9296 0 _029_
rlabel metal3 11760 8764 11760 8764 0 _030_
rlabel metal3 12628 8820 12628 8820 0 _031_
rlabel metal2 13524 10780 13524 10780 0 _032_
rlabel metal2 11284 9772 11284 9772 0 _033_
rlabel metal3 11536 8820 11536 8820 0 _034_
rlabel metal2 10584 7252 10584 7252 0 _035_
rlabel metal2 10668 8204 10668 8204 0 _036_
rlabel metal2 9660 8820 9660 8820 0 _037_
rlabel metal2 10892 9240 10892 9240 0 _038_
rlabel metal3 11732 10052 11732 10052 0 _039_
rlabel metal3 9632 7924 9632 7924 0 _040_
rlabel metal2 9940 8120 9940 8120 0 _041_
rlabel metal2 8876 8064 8876 8064 0 _042_
rlabel metal2 13132 10192 13132 10192 0 _043_
rlabel metal2 13580 11200 13580 11200 0 _044_
rlabel metal2 13356 10584 13356 10584 0 _045_
rlabel metal2 13748 10892 13748 10892 0 _046_
rlabel metal2 11592 7756 11592 7756 0 _047_
rlabel metal2 11032 12236 11032 12236 0 _048_
rlabel metal3 14028 11172 14028 11172 0 _049_
rlabel metal3 14644 10052 14644 10052 0 _050_
rlabel metal2 13524 10178 13524 10178 0 _051_
rlabel metal2 13468 9520 13468 9520 0 _052_
rlabel metal2 13832 9548 13832 9548 0 _053_
rlabel metal2 12852 11816 12852 11816 0 _054_
rlabel metal2 13972 12544 13972 12544 0 _055_
rlabel metal2 14140 11396 14140 11396 0 _056_
rlabel metal2 14588 12292 14588 12292 0 _057_
rlabel metal3 14532 11956 14532 11956 0 _058_
rlabel metal2 10752 12460 10752 12460 0 _059_
rlabel metal2 13132 12936 13132 12936 0 _060_
rlabel metal3 14504 12740 14504 12740 0 _061_
rlabel metal2 10864 7252 10864 7252 0 _062_
rlabel metal2 7532 11564 7532 11564 0 _063_
rlabel metal2 8904 12460 8904 12460 0 _064_
rlabel metal2 7644 12432 7644 12432 0 _065_
rlabel metal2 8596 12880 8596 12880 0 _066_
rlabel metal2 8484 9520 8484 9520 0 _067_
rlabel metal2 6748 9800 6748 9800 0 _068_
rlabel metal2 6804 8624 6804 8624 0 _069_
rlabel metal2 8064 14028 8064 14028 0 _070_
rlabel metal2 8036 11060 8036 11060 0 _071_
rlabel metal2 7672 12068 7672 12068 0 _072_
rlabel metal2 10668 9800 10668 9800 0 _073_
rlabel metal2 12628 9240 12628 9240 0 _074_
rlabel metal2 10780 9408 10780 9408 0 _075_
rlabel metal2 8876 11676 8876 11676 0 _076_
rlabel metal3 12908 7532 12908 7532 0 _077_
rlabel metal2 11004 9240 11004 9240 0 _078_
rlabel metal3 8484 11564 8484 11564 0 _079_
rlabel metal2 9996 9856 9996 9856 0 _080_
rlabel metal2 9156 11228 9156 11228 0 _081_
rlabel metal2 10724 11396 10724 11396 0 _082_
rlabel metal3 11256 11564 11256 11564 0 _083_
rlabel metal3 9072 11564 9072 11564 0 _084_
rlabel metal2 7336 12012 7336 12012 0 _085_
rlabel metal3 12068 9604 12068 9604 0 _086_
rlabel metal2 9660 9632 9660 9632 0 _087_
rlabel metal2 7588 11228 7588 11228 0 _088_
rlabel metal2 13076 9464 13076 9464 0 _089_
rlabel metal2 13524 8400 13524 8400 0 _090_
rlabel metal2 12292 10080 12292 10080 0 _091_
rlabel metal2 11844 10360 11844 10360 0 _092_
rlabel metal2 9156 12012 9156 12012 0 _093_
rlabel metal2 7644 11452 7644 11452 0 _094_
rlabel metal2 12824 7196 12824 7196 0 _095_
rlabel metal2 13468 9268 13468 9268 0 _096_
rlabel metal2 8148 8932 8148 8932 0 _097_
rlabel metal2 11004 8064 11004 8064 0 _098_
rlabel metal2 8008 8932 8008 8932 0 _099_
rlabel metal2 8288 8876 8288 8876 0 _100_
rlabel metal3 8092 10332 8092 10332 0 _101_
rlabel metal2 7924 11060 7924 11060 0 _102_
rlabel metal2 7644 9996 7644 9996 0 _103_
rlabel metal3 10864 10780 10864 10780 0 _104_
rlabel metal2 11508 12824 11508 12824 0 _105_
rlabel metal2 12292 12012 12292 12012 0 _106_
rlabel metal2 11116 13482 11116 13482 0 _107_
rlabel metal2 12908 11368 12908 11368 0 _108_
rlabel metal2 11732 11424 11732 11424 0 _109_
rlabel metal2 11788 11452 11788 11452 0 _110_
rlabel metal3 11592 7924 11592 7924 0 _111_
rlabel metal2 11284 11676 11284 11676 0 _112_
rlabel metal3 1239 13468 1239 13468 0 clk
rlabel metal2 12600 10332 12600 10332 0 clknet_0_clk
rlabel metal2 10276 13972 10276 13972 0 clknet_1_0__leaf_clk
rlabel metal2 15680 10724 15680 10724 0 clknet_1_1__leaf_clk
rlabel metal3 13916 7140 13916 7140 0 dut50.count\[0\]
rlabel metal2 13356 6888 13356 6888 0 dut50.count\[1\]
rlabel metal3 9576 9212 9576 9212 0 dut50.count\[2\]
rlabel metal3 8960 9940 8960 9940 0 dut50.count\[3\]
rlabel metal2 15484 9800 15484 9800 0 net1
rlabel metal2 11004 16030 11004 16030 0 net10
rlabel metal2 13692 13412 13692 13412 0 net11
rlabel metal3 9296 6804 9296 6804 0 net12
rlabel metal2 9016 13580 9016 13580 0 net13
rlabel metal3 3724 9940 3724 9940 0 net14
rlabel metal2 10668 3374 10668 3374 0 net15
rlabel metal2 14084 8596 14084 8596 0 net16
rlabel metal2 15428 9128 15428 9128 0 net17
rlabel metal3 12012 13860 12012 13860 0 net18
rlabel metal2 5796 10948 5796 10948 0 net19
rlabel metal2 8400 14028 8400 14028 0 net2
rlabel metal2 7588 11536 7588 11536 0 net20
rlabel metal2 6132 12712 6132 12712 0 net21
rlabel metal2 9352 15960 9352 15960 0 net22
rlabel metal2 11788 18956 11788 18956 0 net23
rlabel metal2 20132 18592 20132 18592 0 net24
rlabel metal2 20132 2408 20132 2408 0 net25
rlabel metal3 623 2380 623 2380 0 net26
rlabel metal2 14084 12264 14084 12264 0 net3
rlabel metal2 15372 12880 15372 12880 0 net4
rlabel metal2 5684 8596 5684 8596 0 net5
rlabel metal2 11704 6916 11704 6916 0 net6
rlabel metal2 11116 3178 11116 3178 0 net7
rlabel metal2 15708 12096 15708 12096 0 net8
rlabel metal2 15484 10752 15484 10752 0 net9
rlabel metal2 20020 10276 20020 10276 0 segm[10]
rlabel metal2 8428 19481 8428 19481 0 segm[11]
rlabel metal2 20020 11900 20020 11900 0 segm[12]
rlabel metal2 19964 12936 19964 12936 0 segm[13]
rlabel metal3 679 8764 679 8764 0 segm[2]
rlabel metal2 11116 1043 11116 1043 0 segm[3]
rlabel metal2 10780 1211 10780 1211 0 segm[5]
rlabel metal2 20020 12628 20020 12628 0 segm[6]
rlabel metal2 20020 11172 20020 11172 0 segm[7]
rlabel metal2 10780 19677 10780 19677 0 segm[8]
rlabel metal2 20020 13356 20020 13356 0 segm[9]
rlabel metal2 9436 1211 9436 1211 0 sel[0]
rlabel metal2 9100 19873 9100 19873 0 sel[10]
rlabel metal3 679 10108 679 10108 0 sel[11]
rlabel metal2 10444 1491 10444 1491 0 sel[1]
rlabel metal2 20020 8820 20020 8820 0 sel[2]
rlabel metal3 20321 9100 20321 9100 0 sel[3]
rlabel metal2 11452 19873 11452 19873 0 sel[4]
rlabel metal3 679 11116 679 11116 0 sel[5]
rlabel metal3 679 11452 679 11452 0 sel[6]
rlabel metal3 679 12796 679 12796 0 sel[7]
rlabel metal3 9688 18732 9688 18732 0 sel[8]
rlabel metal2 11116 19845 11116 19845 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
