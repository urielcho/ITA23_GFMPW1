magic
tech gf180mcuD
magscale 1 10
timestamp 1699641651
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 18834 38110 18846 38162
rect 18898 38110 18910 38162
rect 22194 38110 22206 38162
rect 22258 38110 22270 38162
rect 17826 37998 17838 38050
rect 17890 37998 17902 38050
rect 23650 37998 23662 38050
rect 23714 37998 23726 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 18734 37490 18786 37502
rect 18734 37426 18786 37438
rect 22094 37490 22146 37502
rect 22094 37426 22146 37438
rect 27470 37490 27522 37502
rect 27470 37426 27522 37438
rect 17714 37214 17726 37266
rect 17778 37214 17790 37266
rect 21522 37214 21534 37266
rect 21586 37214 21598 37266
rect 26450 37214 26462 37266
rect 26514 37214 26526 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 40238 36370 40290 36382
rect 40238 36306 40290 36318
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 21522 28590 21534 28642
rect 21586 28590 21598 28642
rect 21310 28418 21362 28430
rect 21310 28354 21362 28366
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 17502 28082 17554 28094
rect 17502 28018 17554 28030
rect 25230 27970 25282 27982
rect 20738 27918 20750 27970
rect 20802 27918 20814 27970
rect 25230 27906 25282 27918
rect 17278 27858 17330 27870
rect 17278 27794 17330 27806
rect 17614 27858 17666 27870
rect 23438 27858 23490 27870
rect 19954 27806 19966 27858
rect 20018 27806 20030 27858
rect 25442 27806 25454 27858
rect 25506 27806 25518 27858
rect 17614 27794 17666 27806
rect 23438 27794 23490 27806
rect 22866 27694 22878 27746
rect 22930 27694 22942 27746
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 20738 27246 20750 27298
rect 20802 27246 20814 27298
rect 40014 27186 40066 27198
rect 15922 27134 15934 27186
rect 15986 27134 15998 27186
rect 24322 27134 24334 27186
rect 24386 27134 24398 27186
rect 26450 27134 26462 27186
rect 26514 27134 26526 27186
rect 40014 27122 40066 27134
rect 19294 27074 19346 27086
rect 18834 27022 18846 27074
rect 18898 27022 18910 27074
rect 19294 27010 19346 27022
rect 20190 27074 20242 27086
rect 20190 27010 20242 27022
rect 20414 27074 20466 27086
rect 20414 27010 20466 27022
rect 21422 27074 21474 27086
rect 21422 27010 21474 27022
rect 21758 27074 21810 27086
rect 23538 27022 23550 27074
rect 23602 27022 23614 27074
rect 28242 27022 28254 27074
rect 28306 27022 28318 27074
rect 37650 27022 37662 27074
rect 37714 27022 37726 27074
rect 21758 27010 21810 27022
rect 26910 26962 26962 26974
rect 18050 26910 18062 26962
rect 18114 26910 18126 26962
rect 21970 26910 21982 26962
rect 22034 26910 22046 26962
rect 22418 26910 22430 26962
rect 22482 26910 22494 26962
rect 28466 26910 28478 26962
rect 28530 26910 28542 26962
rect 26910 26898 26962 26910
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 24658 26462 24670 26514
rect 24722 26462 24734 26514
rect 17950 26402 18002 26414
rect 17950 26338 18002 26350
rect 17838 26290 17890 26302
rect 24110 26290 24162 26302
rect 4050 26238 4062 26290
rect 4114 26238 4126 26290
rect 14018 26238 14030 26290
rect 14082 26238 14094 26290
rect 23874 26238 23886 26290
rect 23938 26238 23950 26290
rect 17838 26226 17890 26238
rect 24110 26226 24162 26238
rect 24222 26290 24274 26302
rect 24222 26226 24274 26238
rect 25342 26290 25394 26302
rect 25778 26238 25790 26290
rect 25842 26238 25854 26290
rect 37874 26238 37886 26290
rect 37938 26238 37950 26290
rect 25342 26226 25394 26238
rect 17614 26178 17666 26190
rect 14690 26126 14702 26178
rect 14754 26126 14766 26178
rect 16818 26126 16830 26178
rect 16882 26126 16894 26178
rect 26450 26126 26462 26178
rect 26514 26126 26526 26178
rect 28578 26126 28590 26178
rect 28642 26126 28654 26178
rect 39890 26126 39902 26178
rect 39954 26126 39966 26178
rect 17614 26114 17666 26126
rect 1934 26066 1986 26078
rect 17950 26066 18002 26078
rect 17266 26014 17278 26066
rect 17330 26063 17342 26066
rect 17490 26063 17502 26066
rect 17330 26017 17502 26063
rect 17330 26014 17342 26017
rect 17490 26014 17502 26017
rect 17554 26014 17566 26066
rect 1934 26002 1986 26014
rect 17950 26002 18002 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 24334 25730 24386 25742
rect 24334 25666 24386 25678
rect 21982 25618 22034 25630
rect 2034 25566 2046 25618
rect 2098 25566 2110 25618
rect 13458 25566 13470 25618
rect 13522 25566 13534 25618
rect 20738 25566 20750 25618
rect 20802 25566 20814 25618
rect 21982 25554 22034 25566
rect 24894 25618 24946 25630
rect 24894 25554 24946 25566
rect 26686 25618 26738 25630
rect 26686 25554 26738 25566
rect 27582 25618 27634 25630
rect 27582 25554 27634 25566
rect 16606 25506 16658 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 16370 25454 16382 25506
rect 16434 25454 16446 25506
rect 16606 25442 16658 25454
rect 16942 25506 16994 25518
rect 16942 25442 16994 25454
rect 17278 25506 17330 25518
rect 17278 25442 17330 25454
rect 17614 25506 17666 25518
rect 24670 25506 24722 25518
rect 17938 25454 17950 25506
rect 18002 25454 18014 25506
rect 17614 25442 17666 25454
rect 24670 25442 24722 25454
rect 26126 25506 26178 25518
rect 26126 25442 26178 25454
rect 12910 25394 12962 25406
rect 16830 25394 16882 25406
rect 15586 25342 15598 25394
rect 15650 25342 15662 25394
rect 12910 25330 12962 25342
rect 16830 25330 16882 25342
rect 17390 25394 17442 25406
rect 21422 25394 21474 25406
rect 18610 25342 18622 25394
rect 18674 25342 18686 25394
rect 17390 25330 17442 25342
rect 21422 25330 21474 25342
rect 21534 25394 21586 25406
rect 21534 25330 21586 25342
rect 26798 25394 26850 25406
rect 26798 25330 26850 25342
rect 12798 25282 12850 25294
rect 12798 25218 12850 25230
rect 21198 25282 21250 25294
rect 23774 25282 23826 25294
rect 23426 25230 23438 25282
rect 23490 25230 23502 25282
rect 21198 25218 21250 25230
rect 23774 25218 23826 25230
rect 26574 25282 26626 25294
rect 26574 25218 26626 25230
rect 27470 25282 27522 25294
rect 27470 25218 27522 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 15486 24946 15538 24958
rect 15486 24882 15538 24894
rect 15598 24946 15650 24958
rect 15598 24882 15650 24894
rect 16606 24946 16658 24958
rect 19966 24946 20018 24958
rect 17602 24894 17614 24946
rect 17666 24894 17678 24946
rect 16606 24882 16658 24894
rect 19966 24882 20018 24894
rect 12786 24782 12798 24834
rect 12850 24782 12862 24834
rect 15710 24722 15762 24734
rect 19854 24722 19906 24734
rect 12114 24670 12126 24722
rect 12178 24670 12190 24722
rect 15250 24670 15262 24722
rect 15314 24670 15326 24722
rect 15922 24670 15934 24722
rect 15986 24670 15998 24722
rect 17826 24670 17838 24722
rect 17890 24670 17902 24722
rect 15710 24658 15762 24670
rect 19854 24658 19906 24670
rect 20078 24722 20130 24734
rect 20078 24658 20130 24670
rect 20526 24722 20578 24734
rect 20526 24658 20578 24670
rect 14914 24558 14926 24610
rect 14978 24558 14990 24610
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 13918 24162 13970 24174
rect 13918 24098 13970 24110
rect 15150 24050 15202 24062
rect 15150 23986 15202 23998
rect 25342 24050 25394 24062
rect 40014 24050 40066 24062
rect 28578 23998 28590 24050
rect 28642 23998 28654 24050
rect 25342 23986 25394 23998
rect 40014 23986 40066 23998
rect 14590 23938 14642 23950
rect 22306 23886 22318 23938
rect 22370 23886 22382 23938
rect 25666 23886 25678 23938
rect 25730 23886 25742 23938
rect 37874 23886 37886 23938
rect 37938 23886 37950 23938
rect 14590 23874 14642 23886
rect 14030 23826 14082 23838
rect 14030 23762 14082 23774
rect 14254 23826 14306 23838
rect 14254 23762 14306 23774
rect 14478 23826 14530 23838
rect 14478 23762 14530 23774
rect 21982 23826 22034 23838
rect 26450 23774 26462 23826
rect 26514 23774 26526 23826
rect 21982 23762 22034 23774
rect 13918 23714 13970 23726
rect 13918 23650 13970 23662
rect 22094 23714 22146 23726
rect 22094 23650 22146 23662
rect 22654 23714 22706 23726
rect 22978 23662 22990 23714
rect 23042 23662 23054 23714
rect 22654 23650 22706 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 15598 23378 15650 23390
rect 19742 23378 19794 23390
rect 17378 23326 17390 23378
rect 17442 23326 17454 23378
rect 15598 23314 15650 23326
rect 19742 23314 19794 23326
rect 23550 23378 23602 23390
rect 23550 23314 23602 23326
rect 26014 23378 26066 23390
rect 26014 23314 26066 23326
rect 17950 23266 18002 23278
rect 17950 23202 18002 23214
rect 18734 23266 18786 23278
rect 18734 23202 18786 23214
rect 19518 23266 19570 23278
rect 19518 23202 19570 23214
rect 24110 23266 24162 23278
rect 24110 23202 24162 23214
rect 24222 23266 24274 23278
rect 24222 23202 24274 23214
rect 17838 23154 17890 23166
rect 12338 23102 12350 23154
rect 12402 23102 12414 23154
rect 17838 23090 17890 23102
rect 18062 23154 18114 23166
rect 18062 23090 18114 23102
rect 18510 23154 18562 23166
rect 24446 23154 24498 23166
rect 20290 23102 20302 23154
rect 20354 23102 20366 23154
rect 26338 23102 26350 23154
rect 26402 23102 26414 23154
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 18510 23090 18562 23102
rect 24446 23090 24498 23102
rect 13010 22990 13022 23042
rect 13074 22990 13086 23042
rect 15138 22990 15150 23042
rect 15202 22990 15214 23042
rect 18834 22990 18846 23042
rect 18898 22990 18910 23042
rect 20962 22990 20974 23042
rect 21026 22990 21038 23042
rect 23090 22990 23102 23042
rect 23154 22990 23166 23042
rect 27122 22990 27134 23042
rect 27186 22990 27198 23042
rect 29250 22990 29262 23042
rect 29314 22990 29326 23042
rect 19854 22930 19906 22942
rect 19854 22866 19906 22878
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 27134 22594 27186 22606
rect 20178 22542 20190 22594
rect 20242 22542 20254 22594
rect 27134 22530 27186 22542
rect 14142 22482 14194 22494
rect 14142 22418 14194 22430
rect 16270 22482 16322 22494
rect 16270 22418 16322 22430
rect 20638 22482 20690 22494
rect 27470 22482 27522 22494
rect 26338 22430 26350 22482
rect 26402 22430 26414 22482
rect 20638 22418 20690 22430
rect 27470 22418 27522 22430
rect 27918 22482 27970 22494
rect 27918 22418 27970 22430
rect 40014 22482 40066 22494
rect 40014 22418 40066 22430
rect 18846 22370 18898 22382
rect 17378 22318 17390 22370
rect 17442 22318 17454 22370
rect 19058 22318 19070 22370
rect 19122 22318 19134 22370
rect 19954 22318 19966 22370
rect 20018 22318 20030 22370
rect 21858 22318 21870 22370
rect 21922 22318 21934 22370
rect 28130 22318 28142 22370
rect 28194 22318 28206 22370
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 18846 22306 18898 22318
rect 16382 22258 16434 22270
rect 20750 22258 20802 22270
rect 17714 22206 17726 22258
rect 17778 22206 17790 22258
rect 18050 22206 18062 22258
rect 18114 22206 18126 22258
rect 20514 22206 20526 22258
rect 20578 22206 20590 22258
rect 16382 22194 16434 22206
rect 20750 22194 20802 22206
rect 27806 22258 27858 22270
rect 27806 22194 27858 22206
rect 13806 22146 13858 22158
rect 13806 22082 13858 22094
rect 14030 22146 14082 22158
rect 14030 22082 14082 22094
rect 14254 22146 14306 22158
rect 14254 22082 14306 22094
rect 14702 22146 14754 22158
rect 14702 22082 14754 22094
rect 17054 22146 17106 22158
rect 18958 22146 19010 22158
rect 18386 22094 18398 22146
rect 18450 22094 18462 22146
rect 17054 22082 17106 22094
rect 18958 22082 19010 22094
rect 27246 22146 27298 22158
rect 27246 22082 27298 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 15038 21810 15090 21822
rect 15038 21746 15090 21758
rect 24446 21810 24498 21822
rect 24446 21746 24498 21758
rect 27134 21810 27186 21822
rect 27134 21746 27186 21758
rect 27246 21810 27298 21822
rect 27246 21746 27298 21758
rect 14478 21698 14530 21710
rect 14478 21634 14530 21646
rect 15150 21698 15202 21710
rect 16146 21646 16158 21698
rect 16210 21646 16222 21698
rect 16818 21646 16830 21698
rect 16882 21646 16894 21698
rect 21858 21646 21870 21698
rect 21922 21646 21934 21698
rect 15150 21634 15202 21646
rect 14814 21586 14866 21598
rect 23998 21586 24050 21598
rect 10994 21534 11006 21586
rect 11058 21534 11070 21586
rect 15922 21534 15934 21586
rect 15986 21534 15998 21586
rect 16594 21534 16606 21586
rect 16658 21534 16670 21586
rect 17490 21534 17502 21586
rect 17554 21534 17566 21586
rect 18498 21534 18510 21586
rect 18562 21534 18574 21586
rect 14814 21522 14866 21534
rect 23998 21522 24050 21534
rect 24222 21586 24274 21598
rect 24222 21522 24274 21534
rect 26014 21586 26066 21598
rect 26014 21522 26066 21534
rect 26238 21586 26290 21598
rect 26238 21522 26290 21534
rect 26686 21586 26738 21598
rect 37874 21534 37886 21586
rect 37938 21534 37950 21586
rect 26686 21522 26738 21534
rect 14366 21474 14418 21486
rect 24110 21474 24162 21486
rect 11778 21422 11790 21474
rect 11842 21422 11854 21474
rect 13906 21422 13918 21474
rect 13970 21422 13982 21474
rect 17826 21422 17838 21474
rect 17890 21422 17902 21474
rect 14366 21410 14418 21422
rect 24110 21410 24162 21422
rect 26126 21474 26178 21486
rect 26126 21410 26178 21422
rect 26462 21474 26514 21486
rect 26462 21410 26514 21422
rect 27022 21474 27074 21486
rect 39890 21422 39902 21474
rect 39954 21422 39966 21474
rect 27022 21410 27074 21422
rect 14254 21362 14306 21374
rect 14254 21298 14306 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 20638 21026 20690 21038
rect 20638 20962 20690 20974
rect 21422 21026 21474 21038
rect 21422 20962 21474 20974
rect 22206 20914 22258 20926
rect 26686 20914 26738 20926
rect 15250 20862 15262 20914
rect 15314 20862 15326 20914
rect 23426 20862 23438 20914
rect 23490 20862 23502 20914
rect 25554 20862 25566 20914
rect 25618 20862 25630 20914
rect 26226 20862 26238 20914
rect 26290 20862 26302 20914
rect 22206 20850 22258 20862
rect 26686 20850 26738 20862
rect 40014 20914 40066 20926
rect 40014 20850 40066 20862
rect 22430 20802 22482 20814
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 22082 20750 22094 20802
rect 22146 20750 22158 20802
rect 22754 20750 22766 20802
rect 22818 20750 22830 20802
rect 37650 20750 37662 20802
rect 37714 20750 37726 20802
rect 22430 20738 22482 20750
rect 20526 20690 20578 20702
rect 14466 20638 14478 20690
rect 14530 20638 14542 20690
rect 20526 20626 20578 20638
rect 21310 20690 21362 20702
rect 21310 20626 21362 20638
rect 21870 20690 21922 20702
rect 21870 20626 21922 20638
rect 25902 20690 25954 20702
rect 25902 20626 25954 20638
rect 14142 20578 14194 20590
rect 14142 20514 14194 20526
rect 20638 20578 20690 20590
rect 20638 20514 20690 20526
rect 21422 20578 21474 20590
rect 21422 20514 21474 20526
rect 26126 20578 26178 20590
rect 26126 20514 26178 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 19170 20190 19182 20242
rect 19234 20190 19246 20242
rect 15262 20130 15314 20142
rect 15262 20066 15314 20078
rect 15374 20130 15426 20142
rect 15374 20066 15426 20078
rect 15934 20130 15986 20142
rect 15934 20066 15986 20078
rect 16158 20130 16210 20142
rect 16158 20066 16210 20078
rect 16494 20130 16546 20142
rect 23886 20130 23938 20142
rect 16818 20078 16830 20130
rect 16882 20078 16894 20130
rect 18162 20078 18174 20130
rect 18226 20078 18238 20130
rect 19282 20078 19294 20130
rect 19346 20078 19358 20130
rect 19842 20078 19854 20130
rect 19906 20078 19918 20130
rect 20850 20078 20862 20130
rect 20914 20078 20926 20130
rect 23202 20078 23214 20130
rect 23266 20078 23278 20130
rect 16494 20066 16546 20078
rect 23886 20066 23938 20078
rect 24110 20130 24162 20142
rect 24110 20066 24162 20078
rect 24222 20130 24274 20142
rect 26226 20078 26238 20130
rect 26290 20078 26302 20130
rect 29026 20078 29038 20130
rect 29090 20078 29102 20130
rect 24222 20066 24274 20078
rect 14030 20018 14082 20030
rect 19070 20018 19122 20030
rect 22878 20018 22930 20030
rect 17266 19966 17278 20018
rect 17330 19966 17342 20018
rect 18386 19966 18398 20018
rect 18450 19966 18462 20018
rect 20514 19966 20526 20018
rect 20578 19966 20590 20018
rect 14030 19954 14082 19966
rect 19070 19954 19122 19966
rect 22878 19954 22930 19966
rect 24334 20018 24386 20030
rect 24546 19966 24558 20018
rect 24610 19966 24622 20018
rect 25442 19966 25454 20018
rect 25506 19966 25518 20018
rect 28802 19966 28814 20018
rect 28866 19966 28878 20018
rect 24334 19954 24386 19966
rect 13134 19906 13186 19918
rect 13806 19906 13858 19918
rect 13346 19854 13358 19906
rect 13410 19854 13422 19906
rect 15810 19854 15822 19906
rect 15874 19854 15886 19906
rect 17938 19854 17950 19906
rect 18002 19854 18014 19906
rect 20962 19854 20974 19906
rect 21026 19854 21038 19906
rect 28354 19854 28366 19906
rect 28418 19854 28430 19906
rect 13134 19842 13186 19854
rect 13806 19842 13858 19854
rect 15374 19794 15426 19806
rect 14354 19742 14366 19794
rect 14418 19742 14430 19794
rect 15374 19730 15426 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 17166 19458 17218 19470
rect 17166 19394 17218 19406
rect 17838 19458 17890 19470
rect 17838 19394 17890 19406
rect 18174 19458 18226 19470
rect 18174 19394 18226 19406
rect 13582 19346 13634 19358
rect 10770 19294 10782 19346
rect 10834 19294 10846 19346
rect 12898 19294 12910 19346
rect 12962 19294 12974 19346
rect 13582 19282 13634 19294
rect 25118 19346 25170 19358
rect 25118 19282 25170 19294
rect 40014 19346 40066 19358
rect 40014 19282 40066 19294
rect 18510 19234 18562 19246
rect 22206 19234 22258 19246
rect 10098 19182 10110 19234
rect 10162 19182 10174 19234
rect 14130 19182 14142 19234
rect 14194 19182 14206 19234
rect 15362 19182 15374 19234
rect 15426 19182 15438 19234
rect 15810 19182 15822 19234
rect 15874 19182 15886 19234
rect 16482 19182 16494 19234
rect 16546 19182 16558 19234
rect 18162 19182 18174 19234
rect 18226 19182 18238 19234
rect 19282 19182 19294 19234
rect 19346 19182 19358 19234
rect 20066 19182 20078 19234
rect 20130 19182 20142 19234
rect 20514 19182 20526 19234
rect 20578 19182 20590 19234
rect 18510 19170 18562 19182
rect 22206 19170 22258 19182
rect 22430 19234 22482 19246
rect 22430 19170 22482 19182
rect 22766 19234 22818 19246
rect 22766 19170 22818 19182
rect 25454 19234 25506 19246
rect 37650 19182 37662 19234
rect 37714 19182 37726 19234
rect 25454 19170 25506 19182
rect 20862 19122 20914 19134
rect 14354 19070 14366 19122
rect 14418 19070 14430 19122
rect 18834 19070 18846 19122
rect 18898 19070 18910 19122
rect 19394 19070 19406 19122
rect 19458 19070 19470 19122
rect 20862 19058 20914 19070
rect 25902 19122 25954 19134
rect 25902 19058 25954 19070
rect 26126 19122 26178 19134
rect 26126 19058 26178 19070
rect 26462 19122 26514 19134
rect 26462 19058 26514 19070
rect 26574 19122 26626 19134
rect 26574 19058 26626 19070
rect 15934 19010 15986 19022
rect 17278 19010 17330 19022
rect 16706 18958 16718 19010
rect 16770 18958 16782 19010
rect 15934 18946 15986 18958
rect 17278 18946 17330 18958
rect 17390 19010 17442 19022
rect 17390 18946 17442 18958
rect 22318 19010 22370 19022
rect 22318 18946 22370 18958
rect 25790 19010 25842 19022
rect 25790 18946 25842 18958
rect 26798 19010 26850 19022
rect 26798 18946 26850 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 20414 18674 20466 18686
rect 18386 18622 18398 18674
rect 18450 18622 18462 18674
rect 18834 18622 18846 18674
rect 18898 18622 18910 18674
rect 20414 18610 20466 18622
rect 24670 18674 24722 18686
rect 24670 18610 24722 18622
rect 16158 18562 16210 18574
rect 16158 18498 16210 18510
rect 16606 18562 16658 18574
rect 16606 18498 16658 18510
rect 16718 18562 16770 18574
rect 19966 18562 20018 18574
rect 17714 18510 17726 18562
rect 17778 18510 17790 18562
rect 16718 18498 16770 18510
rect 19966 18498 20018 18510
rect 20302 18562 20354 18574
rect 22082 18510 22094 18562
rect 22146 18510 22158 18562
rect 26114 18510 26126 18562
rect 26178 18510 26190 18562
rect 20302 18498 20354 18510
rect 14478 18450 14530 18462
rect 14478 18386 14530 18398
rect 14702 18450 14754 18462
rect 14702 18386 14754 18398
rect 15038 18450 15090 18462
rect 19182 18450 19234 18462
rect 17378 18398 17390 18450
rect 17442 18398 17454 18450
rect 18274 18398 18286 18450
rect 18338 18398 18350 18450
rect 15038 18386 15090 18398
rect 19182 18386 19234 18398
rect 19630 18450 19682 18462
rect 21410 18398 21422 18450
rect 21474 18398 21486 18450
rect 25330 18398 25342 18450
rect 25394 18398 25406 18450
rect 19630 18386 19682 18398
rect 14590 18338 14642 18350
rect 24210 18286 24222 18338
rect 24274 18286 24286 18338
rect 28242 18286 28254 18338
rect 28306 18286 28318 18338
rect 14590 18274 14642 18286
rect 16270 18226 16322 18238
rect 16270 18162 16322 18174
rect 16718 18226 16770 18238
rect 16718 18162 16770 18174
rect 20414 18226 20466 18238
rect 20414 18162 20466 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 20190 17890 20242 17902
rect 17154 17838 17166 17890
rect 17218 17887 17230 17890
rect 17714 17887 17726 17890
rect 17218 17841 17726 17887
rect 17218 17838 17230 17841
rect 17714 17838 17726 17841
rect 17778 17838 17790 17890
rect 20190 17826 20242 17838
rect 17390 17778 17442 17790
rect 25006 17778 25058 17790
rect 14242 17726 14254 17778
rect 14306 17726 14318 17778
rect 16370 17726 16382 17778
rect 16434 17726 16446 17778
rect 19842 17726 19854 17778
rect 19906 17726 19918 17778
rect 22306 17726 22318 17778
rect 22370 17726 22382 17778
rect 17390 17714 17442 17726
rect 25006 17714 25058 17726
rect 16942 17666 16994 17678
rect 19518 17666 19570 17678
rect 22766 17666 22818 17678
rect 13570 17614 13582 17666
rect 13634 17614 13646 17666
rect 18162 17614 18174 17666
rect 18226 17614 18238 17666
rect 21970 17614 21982 17666
rect 22034 17614 22046 17666
rect 16942 17602 16994 17614
rect 19518 17602 19570 17614
rect 22766 17602 22818 17614
rect 22990 17666 23042 17678
rect 22990 17602 23042 17614
rect 23438 17666 23490 17678
rect 23438 17602 23490 17614
rect 19966 17554 20018 17566
rect 17938 17502 17950 17554
rect 18002 17502 18014 17554
rect 19966 17490 20018 17502
rect 21758 17554 21810 17566
rect 22082 17502 22094 17554
rect 22146 17502 22158 17554
rect 21758 17490 21810 17502
rect 16606 17442 16658 17454
rect 16606 17378 16658 17390
rect 16830 17442 16882 17454
rect 21534 17442 21586 17454
rect 19170 17390 19182 17442
rect 19234 17390 19246 17442
rect 16830 17378 16882 17390
rect 21534 17378 21586 17390
rect 23102 17442 23154 17454
rect 23102 17378 23154 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 18286 17106 18338 17118
rect 25342 17106 25394 17118
rect 18610 17054 18622 17106
rect 18674 17054 18686 17106
rect 27234 17054 27246 17106
rect 27298 17054 27310 17106
rect 18286 17042 18338 17054
rect 25342 17042 25394 17054
rect 15150 16994 15202 17006
rect 15150 16930 15202 16942
rect 23886 16994 23938 17006
rect 23886 16930 23938 16942
rect 24110 16994 24162 17006
rect 24110 16930 24162 16942
rect 26686 16994 26738 17006
rect 26686 16930 26738 16942
rect 23550 16882 23602 16894
rect 4274 16830 4286 16882
rect 4338 16830 4350 16882
rect 14802 16830 14814 16882
rect 14866 16830 14878 16882
rect 23550 16818 23602 16830
rect 25790 16882 25842 16894
rect 25790 16818 25842 16830
rect 26014 16882 26066 16894
rect 37874 16830 37886 16882
rect 37938 16830 37950 16882
rect 26014 16818 26066 16830
rect 15038 16770 15090 16782
rect 39890 16718 39902 16770
rect 39954 16718 39966 16770
rect 15038 16706 15090 16718
rect 1934 16658 1986 16670
rect 1934 16594 1986 16606
rect 23774 16658 23826 16670
rect 26910 16658 26962 16670
rect 26338 16606 26350 16658
rect 26402 16606 26414 16658
rect 23774 16594 23826 16606
rect 26910 16594 26962 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 15598 16322 15650 16334
rect 15598 16258 15650 16270
rect 40014 16210 40066 16222
rect 18610 16158 18622 16210
rect 18674 16158 18686 16210
rect 22866 16158 22878 16210
rect 22930 16158 22942 16210
rect 24994 16158 25006 16210
rect 25058 16158 25070 16210
rect 28354 16158 28366 16210
rect 28418 16158 28430 16210
rect 40014 16146 40066 16158
rect 15374 16098 15426 16110
rect 15138 16046 15150 16098
rect 15202 16046 15214 16098
rect 22194 16046 22206 16098
rect 22258 16046 22270 16098
rect 25442 16046 25454 16098
rect 25506 16046 25518 16098
rect 37650 16046 37662 16098
rect 37714 16046 37726 16098
rect 15374 16034 15426 16046
rect 18734 15986 18786 15998
rect 18734 15922 18786 15934
rect 18958 15986 19010 15998
rect 26226 15934 26238 15986
rect 26290 15934 26302 15986
rect 18958 15922 19010 15934
rect 15262 15874 15314 15886
rect 15262 15810 15314 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 15486 15538 15538 15550
rect 15486 15474 15538 15486
rect 16382 15538 16434 15550
rect 16382 15474 16434 15486
rect 17502 15538 17554 15550
rect 17502 15474 17554 15486
rect 18622 15538 18674 15550
rect 18622 15474 18674 15486
rect 19070 15538 19122 15550
rect 19070 15474 19122 15486
rect 19182 15538 19234 15550
rect 19182 15474 19234 15486
rect 19518 15538 19570 15550
rect 19518 15474 19570 15486
rect 25342 15538 25394 15550
rect 25342 15474 25394 15486
rect 26014 15538 26066 15550
rect 26014 15474 26066 15486
rect 19966 15426 20018 15438
rect 14242 15374 14254 15426
rect 14306 15374 14318 15426
rect 19966 15362 20018 15374
rect 20974 15426 21026 15438
rect 20974 15362 21026 15374
rect 21086 15426 21138 15438
rect 21086 15362 21138 15374
rect 26350 15426 26402 15438
rect 27794 15374 27806 15426
rect 27858 15374 27870 15426
rect 26350 15362 26402 15374
rect 18174 15314 18226 15326
rect 15026 15262 15038 15314
rect 15090 15262 15102 15314
rect 18174 15250 18226 15262
rect 18398 15314 18450 15326
rect 18398 15250 18450 15262
rect 19294 15314 19346 15326
rect 19294 15250 19346 15262
rect 20302 15314 20354 15326
rect 20302 15250 20354 15262
rect 20526 15314 20578 15326
rect 20526 15250 20578 15262
rect 20750 15314 20802 15326
rect 27570 15262 27582 15314
rect 27634 15262 27646 15314
rect 20750 15250 20802 15262
rect 16606 15202 16658 15214
rect 12114 15150 12126 15202
rect 12178 15150 12190 15202
rect 16258 15150 16270 15202
rect 16322 15150 16334 15202
rect 16606 15138 16658 15150
rect 18286 15202 18338 15214
rect 18286 15138 18338 15150
rect 20414 15202 20466 15214
rect 20414 15138 20466 15150
rect 17266 15038 17278 15090
rect 17330 15087 17342 15090
rect 17938 15087 17950 15090
rect 17330 15041 17950 15087
rect 17330 15038 17342 15041
rect 17938 15038 17950 15041
rect 18002 15038 18014 15090
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 14914 14590 14926 14642
rect 14978 14590 14990 14642
rect 17042 14590 17054 14642
rect 17106 14590 17118 14642
rect 18162 14590 18174 14642
rect 18226 14590 18238 14642
rect 20290 14590 20302 14642
rect 20354 14590 20366 14642
rect 14242 14478 14254 14530
rect 14306 14478 14318 14530
rect 17378 14478 17390 14530
rect 17442 14478 17454 14530
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 17614 13970 17666 13982
rect 17614 13906 17666 13918
rect 19954 13806 19966 13858
rect 20018 13806 20030 13858
rect 22542 13746 22594 13758
rect 19282 13694 19294 13746
rect 19346 13694 19358 13746
rect 22542 13682 22594 13694
rect 22082 13582 22094 13634
rect 22146 13582 22158 13634
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 22318 5234 22370 5246
rect 22318 5170 22370 5182
rect 21298 5070 21310 5122
rect 21362 5070 21374 5122
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 21858 4286 21870 4338
rect 21922 4286 21934 4338
rect 22766 4114 22818 4126
rect 22766 4050 22818 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 18622 3666 18674 3678
rect 18622 3602 18674 3614
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 17602 3502 17614 3554
rect 17666 3502 17678 3554
rect 23538 3502 23550 3554
rect 23602 3502 23614 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 22194 3390 22206 3442
rect 22258 3390 22270 3442
rect 7646 3330 7698 3342
rect 7646 3266 7698 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 25566 38222 25618 38274
rect 18846 38110 18898 38162
rect 22206 38110 22258 38162
rect 17838 37998 17890 38050
rect 23662 37998 23714 38050
rect 24558 37998 24610 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 18734 37438 18786 37490
rect 22094 37438 22146 37490
rect 27470 37438 27522 37490
rect 17726 37214 17778 37266
rect 21534 37214 21586 37266
rect 26462 37214 26514 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 40238 36318 40290 36370
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 21534 28590 21586 28642
rect 21310 28366 21362 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 17502 28030 17554 28082
rect 20750 27918 20802 27970
rect 25230 27918 25282 27970
rect 17278 27806 17330 27858
rect 17614 27806 17666 27858
rect 19966 27806 20018 27858
rect 23438 27806 23490 27858
rect 25454 27806 25506 27858
rect 22878 27694 22930 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 20750 27246 20802 27298
rect 15934 27134 15986 27186
rect 24334 27134 24386 27186
rect 26462 27134 26514 27186
rect 40014 27134 40066 27186
rect 18846 27022 18898 27074
rect 19294 27022 19346 27074
rect 20190 27022 20242 27074
rect 20414 27022 20466 27074
rect 21422 27022 21474 27074
rect 21758 27022 21810 27074
rect 23550 27022 23602 27074
rect 28254 27022 28306 27074
rect 37662 27022 37714 27074
rect 18062 26910 18114 26962
rect 21982 26910 22034 26962
rect 22430 26910 22482 26962
rect 26910 26910 26962 26962
rect 28478 26910 28530 26962
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 24670 26462 24722 26514
rect 17950 26350 18002 26402
rect 4062 26238 4114 26290
rect 14030 26238 14082 26290
rect 17838 26238 17890 26290
rect 23886 26238 23938 26290
rect 24110 26238 24162 26290
rect 24222 26238 24274 26290
rect 25342 26238 25394 26290
rect 25790 26238 25842 26290
rect 37886 26238 37938 26290
rect 14702 26126 14754 26178
rect 16830 26126 16882 26178
rect 17614 26126 17666 26178
rect 26462 26126 26514 26178
rect 28590 26126 28642 26178
rect 39902 26126 39954 26178
rect 1934 26014 1986 26066
rect 17278 26014 17330 26066
rect 17502 26014 17554 26066
rect 17950 26014 18002 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 24334 25678 24386 25730
rect 2046 25566 2098 25618
rect 13470 25566 13522 25618
rect 20750 25566 20802 25618
rect 21982 25566 22034 25618
rect 24894 25566 24946 25618
rect 26686 25566 26738 25618
rect 27582 25566 27634 25618
rect 4286 25454 4338 25506
rect 16382 25454 16434 25506
rect 16606 25454 16658 25506
rect 16942 25454 16994 25506
rect 17278 25454 17330 25506
rect 17614 25454 17666 25506
rect 17950 25454 18002 25506
rect 24670 25454 24722 25506
rect 26126 25454 26178 25506
rect 12910 25342 12962 25394
rect 15598 25342 15650 25394
rect 16830 25342 16882 25394
rect 17390 25342 17442 25394
rect 18622 25342 18674 25394
rect 21422 25342 21474 25394
rect 21534 25342 21586 25394
rect 26798 25342 26850 25394
rect 12798 25230 12850 25282
rect 21198 25230 21250 25282
rect 23438 25230 23490 25282
rect 23774 25230 23826 25282
rect 26574 25230 26626 25282
rect 27470 25230 27522 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 15486 24894 15538 24946
rect 15598 24894 15650 24946
rect 16606 24894 16658 24946
rect 17614 24894 17666 24946
rect 19966 24894 20018 24946
rect 12798 24782 12850 24834
rect 12126 24670 12178 24722
rect 15262 24670 15314 24722
rect 15710 24670 15762 24722
rect 15934 24670 15986 24722
rect 17838 24670 17890 24722
rect 19854 24670 19906 24722
rect 20078 24670 20130 24722
rect 20526 24670 20578 24722
rect 14926 24558 14978 24610
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 13918 24110 13970 24162
rect 15150 23998 15202 24050
rect 25342 23998 25394 24050
rect 28590 23998 28642 24050
rect 40014 23998 40066 24050
rect 14590 23886 14642 23938
rect 22318 23886 22370 23938
rect 25678 23886 25730 23938
rect 37886 23886 37938 23938
rect 14030 23774 14082 23826
rect 14254 23774 14306 23826
rect 14478 23774 14530 23826
rect 21982 23774 22034 23826
rect 26462 23774 26514 23826
rect 13918 23662 13970 23714
rect 22094 23662 22146 23714
rect 22654 23662 22706 23714
rect 22990 23662 23042 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 15598 23326 15650 23378
rect 17390 23326 17442 23378
rect 19742 23326 19794 23378
rect 23550 23326 23602 23378
rect 26014 23326 26066 23378
rect 17950 23214 18002 23266
rect 18734 23214 18786 23266
rect 19518 23214 19570 23266
rect 24110 23214 24162 23266
rect 24222 23214 24274 23266
rect 12350 23102 12402 23154
rect 17838 23102 17890 23154
rect 18062 23102 18114 23154
rect 18510 23102 18562 23154
rect 20302 23102 20354 23154
rect 24446 23102 24498 23154
rect 26350 23102 26402 23154
rect 37662 23102 37714 23154
rect 13022 22990 13074 23042
rect 15150 22990 15202 23042
rect 18846 22990 18898 23042
rect 20974 22990 21026 23042
rect 23102 22990 23154 23042
rect 27134 22990 27186 23042
rect 29262 22990 29314 23042
rect 19854 22878 19906 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 20190 22542 20242 22594
rect 27134 22542 27186 22594
rect 14142 22430 14194 22482
rect 16270 22430 16322 22482
rect 20638 22430 20690 22482
rect 26350 22430 26402 22482
rect 27470 22430 27522 22482
rect 27918 22430 27970 22482
rect 40014 22430 40066 22482
rect 17390 22318 17442 22370
rect 18846 22318 18898 22370
rect 19070 22318 19122 22370
rect 19966 22318 20018 22370
rect 21870 22318 21922 22370
rect 28142 22318 28194 22370
rect 37662 22318 37714 22370
rect 16382 22206 16434 22258
rect 17726 22206 17778 22258
rect 18062 22206 18114 22258
rect 20526 22206 20578 22258
rect 20750 22206 20802 22258
rect 27806 22206 27858 22258
rect 13806 22094 13858 22146
rect 14030 22094 14082 22146
rect 14254 22094 14306 22146
rect 14702 22094 14754 22146
rect 17054 22094 17106 22146
rect 18398 22094 18450 22146
rect 18958 22094 19010 22146
rect 27246 22094 27298 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 15038 21758 15090 21810
rect 24446 21758 24498 21810
rect 27134 21758 27186 21810
rect 27246 21758 27298 21810
rect 14478 21646 14530 21698
rect 15150 21646 15202 21698
rect 16158 21646 16210 21698
rect 16830 21646 16882 21698
rect 21870 21646 21922 21698
rect 11006 21534 11058 21586
rect 14814 21534 14866 21586
rect 15934 21534 15986 21586
rect 16606 21534 16658 21586
rect 17502 21534 17554 21586
rect 18510 21534 18562 21586
rect 23998 21534 24050 21586
rect 24222 21534 24274 21586
rect 26014 21534 26066 21586
rect 26238 21534 26290 21586
rect 26686 21534 26738 21586
rect 37886 21534 37938 21586
rect 11790 21422 11842 21474
rect 13918 21422 13970 21474
rect 14366 21422 14418 21474
rect 17838 21422 17890 21474
rect 24110 21422 24162 21474
rect 26126 21422 26178 21474
rect 26462 21422 26514 21474
rect 27022 21422 27074 21474
rect 39902 21422 39954 21474
rect 14254 21310 14306 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 20638 20974 20690 21026
rect 21422 20974 21474 21026
rect 15262 20862 15314 20914
rect 22206 20862 22258 20914
rect 23438 20862 23490 20914
rect 25566 20862 25618 20914
rect 26238 20862 26290 20914
rect 26686 20862 26738 20914
rect 40014 20862 40066 20914
rect 20078 20750 20130 20802
rect 22094 20750 22146 20802
rect 22430 20750 22482 20802
rect 22766 20750 22818 20802
rect 37662 20750 37714 20802
rect 14478 20638 14530 20690
rect 20526 20638 20578 20690
rect 21310 20638 21362 20690
rect 21870 20638 21922 20690
rect 25902 20638 25954 20690
rect 14142 20526 14194 20578
rect 20638 20526 20690 20578
rect 21422 20526 21474 20578
rect 26126 20526 26178 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 19182 20190 19234 20242
rect 15262 20078 15314 20130
rect 15374 20078 15426 20130
rect 15934 20078 15986 20130
rect 16158 20078 16210 20130
rect 16494 20078 16546 20130
rect 16830 20078 16882 20130
rect 18174 20078 18226 20130
rect 19294 20078 19346 20130
rect 19854 20078 19906 20130
rect 20862 20078 20914 20130
rect 23214 20078 23266 20130
rect 23886 20078 23938 20130
rect 24110 20078 24162 20130
rect 24222 20078 24274 20130
rect 26238 20078 26290 20130
rect 29038 20078 29090 20130
rect 14030 19966 14082 20018
rect 17278 19966 17330 20018
rect 18398 19966 18450 20018
rect 19070 19966 19122 20018
rect 20526 19966 20578 20018
rect 22878 19966 22930 20018
rect 24334 19966 24386 20018
rect 24558 19966 24610 20018
rect 25454 19966 25506 20018
rect 28814 19966 28866 20018
rect 13134 19854 13186 19906
rect 13358 19854 13410 19906
rect 13806 19854 13858 19906
rect 15822 19854 15874 19906
rect 17950 19854 18002 19906
rect 20974 19854 21026 19906
rect 28366 19854 28418 19906
rect 14366 19742 14418 19794
rect 15374 19742 15426 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 17166 19406 17218 19458
rect 17838 19406 17890 19458
rect 18174 19406 18226 19458
rect 10782 19294 10834 19346
rect 12910 19294 12962 19346
rect 13582 19294 13634 19346
rect 25118 19294 25170 19346
rect 40014 19294 40066 19346
rect 10110 19182 10162 19234
rect 14142 19182 14194 19234
rect 15374 19182 15426 19234
rect 15822 19182 15874 19234
rect 16494 19182 16546 19234
rect 18174 19182 18226 19234
rect 18510 19182 18562 19234
rect 19294 19182 19346 19234
rect 20078 19182 20130 19234
rect 20526 19182 20578 19234
rect 22206 19182 22258 19234
rect 22430 19182 22482 19234
rect 22766 19182 22818 19234
rect 25454 19182 25506 19234
rect 37662 19182 37714 19234
rect 14366 19070 14418 19122
rect 18846 19070 18898 19122
rect 19406 19070 19458 19122
rect 20862 19070 20914 19122
rect 25902 19070 25954 19122
rect 26126 19070 26178 19122
rect 26462 19070 26514 19122
rect 26574 19070 26626 19122
rect 15934 18958 15986 19010
rect 16718 18958 16770 19010
rect 17278 18958 17330 19010
rect 17390 18958 17442 19010
rect 22318 18958 22370 19010
rect 25790 18958 25842 19010
rect 26798 18958 26850 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 18398 18622 18450 18674
rect 18846 18622 18898 18674
rect 20414 18622 20466 18674
rect 24670 18622 24722 18674
rect 16158 18510 16210 18562
rect 16606 18510 16658 18562
rect 16718 18510 16770 18562
rect 17726 18510 17778 18562
rect 19966 18510 20018 18562
rect 20302 18510 20354 18562
rect 22094 18510 22146 18562
rect 26126 18510 26178 18562
rect 14478 18398 14530 18450
rect 14702 18398 14754 18450
rect 15038 18398 15090 18450
rect 17390 18398 17442 18450
rect 18286 18398 18338 18450
rect 19182 18398 19234 18450
rect 19630 18398 19682 18450
rect 21422 18398 21474 18450
rect 25342 18398 25394 18450
rect 14590 18286 14642 18338
rect 24222 18286 24274 18338
rect 28254 18286 28306 18338
rect 16270 18174 16322 18226
rect 16718 18174 16770 18226
rect 20414 18174 20466 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 17166 17838 17218 17890
rect 17726 17838 17778 17890
rect 20190 17838 20242 17890
rect 14254 17726 14306 17778
rect 16382 17726 16434 17778
rect 17390 17726 17442 17778
rect 19854 17726 19906 17778
rect 22318 17726 22370 17778
rect 25006 17726 25058 17778
rect 13582 17614 13634 17666
rect 16942 17614 16994 17666
rect 18174 17614 18226 17666
rect 19518 17614 19570 17666
rect 21982 17614 22034 17666
rect 22766 17614 22818 17666
rect 22990 17614 23042 17666
rect 23438 17614 23490 17666
rect 17950 17502 18002 17554
rect 19966 17502 20018 17554
rect 21758 17502 21810 17554
rect 22094 17502 22146 17554
rect 16606 17390 16658 17442
rect 16830 17390 16882 17442
rect 19182 17390 19234 17442
rect 21534 17390 21586 17442
rect 23102 17390 23154 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 18286 17054 18338 17106
rect 18622 17054 18674 17106
rect 25342 17054 25394 17106
rect 27246 17054 27298 17106
rect 15150 16942 15202 16994
rect 23886 16942 23938 16994
rect 24110 16942 24162 16994
rect 26686 16942 26738 16994
rect 4286 16830 4338 16882
rect 14814 16830 14866 16882
rect 23550 16830 23602 16882
rect 25790 16830 25842 16882
rect 26014 16830 26066 16882
rect 37886 16830 37938 16882
rect 15038 16718 15090 16770
rect 39902 16718 39954 16770
rect 1934 16606 1986 16658
rect 23774 16606 23826 16658
rect 26350 16606 26402 16658
rect 26910 16606 26962 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 15598 16270 15650 16322
rect 18622 16158 18674 16210
rect 22878 16158 22930 16210
rect 25006 16158 25058 16210
rect 28366 16158 28418 16210
rect 40014 16158 40066 16210
rect 15150 16046 15202 16098
rect 15374 16046 15426 16098
rect 22206 16046 22258 16098
rect 25454 16046 25506 16098
rect 37662 16046 37714 16098
rect 18734 15934 18786 15986
rect 18958 15934 19010 15986
rect 26238 15934 26290 15986
rect 15262 15822 15314 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 15486 15486 15538 15538
rect 16382 15486 16434 15538
rect 17502 15486 17554 15538
rect 18622 15486 18674 15538
rect 19070 15486 19122 15538
rect 19182 15486 19234 15538
rect 19518 15486 19570 15538
rect 25342 15486 25394 15538
rect 26014 15486 26066 15538
rect 14254 15374 14306 15426
rect 19966 15374 20018 15426
rect 20974 15374 21026 15426
rect 21086 15374 21138 15426
rect 26350 15374 26402 15426
rect 27806 15374 27858 15426
rect 15038 15262 15090 15314
rect 18174 15262 18226 15314
rect 18398 15262 18450 15314
rect 19294 15262 19346 15314
rect 20302 15262 20354 15314
rect 20526 15262 20578 15314
rect 20750 15262 20802 15314
rect 27582 15262 27634 15314
rect 12126 15150 12178 15202
rect 16270 15150 16322 15202
rect 16606 15150 16658 15202
rect 18286 15150 18338 15202
rect 20414 15150 20466 15202
rect 17278 15038 17330 15090
rect 17950 15038 18002 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 14926 14590 14978 14642
rect 17054 14590 17106 14642
rect 18174 14590 18226 14642
rect 20302 14590 20354 14642
rect 14254 14478 14306 14530
rect 17390 14478 17442 14530
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 17614 13918 17666 13970
rect 19966 13806 20018 13858
rect 19294 13694 19346 13746
rect 22542 13694 22594 13746
rect 22094 13582 22146 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 22318 5182 22370 5234
rect 21310 5070 21362 5122
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 21870 4286 21922 4338
rect 22766 4062 22818 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18622 3614 18674 3666
rect 25566 3614 25618 3666
rect 17614 3502 17666 3554
rect 23550 3502 23602 3554
rect 24558 3502 24610 3554
rect 22206 3390 22258 3442
rect 7646 3278 7698 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 17472 41200 17584 42000
rect 18816 41200 18928 42000
rect 20832 41200 20944 42000
rect 22176 41200 22288 42000
rect 22848 41200 22960 42000
rect 26208 41200 26320 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 17500 37492 17556 41200
rect 18844 38162 18900 41200
rect 18844 38110 18846 38162
rect 18898 38110 18900 38162
rect 18844 38098 18900 38110
rect 17500 37426 17556 37436
rect 17836 38050 17892 38062
rect 17836 37998 17838 38050
rect 17890 37998 17892 38050
rect 17724 37266 17780 37278
rect 17724 37214 17726 37266
rect 17778 37214 17780 37266
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 17724 34580 17780 37214
rect 17500 34524 17780 34580
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 15932 28084 15988 28094
rect 17500 28084 17556 34524
rect 17836 32004 17892 37998
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 18732 37492 18788 37502
rect 18732 37398 18788 37436
rect 20860 37492 20916 41200
rect 22204 38162 22260 41200
rect 22876 38276 22932 41200
rect 22876 38210 22932 38220
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 22204 38110 22206 38162
rect 22258 38110 22260 38162
rect 22204 38098 22260 38110
rect 23660 38050 23716 38062
rect 23660 37998 23662 38050
rect 23714 37998 23716 38050
rect 20860 37426 20916 37436
rect 22092 37492 22148 37502
rect 22092 37398 22148 37436
rect 21532 37268 21588 37278
rect 21532 37266 21700 37268
rect 21532 37214 21534 37266
rect 21586 37214 21700 37266
rect 21532 37212 21700 37214
rect 21532 37202 21588 37212
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 17724 31948 17892 32004
rect 4172 27636 4228 27646
rect 4060 26290 4116 26302
rect 4060 26238 4062 26290
rect 4114 26238 4116 26290
rect 1932 26066 1988 26078
rect 1932 26014 1934 26066
rect 1986 26014 1988 26066
rect 1932 25620 1988 26014
rect 1932 25554 1988 25564
rect 2044 25618 2100 25630
rect 2044 25566 2046 25618
rect 2098 25566 2100 25618
rect 2044 24948 2100 25566
rect 2044 24882 2100 24892
rect 4060 24612 4116 26238
rect 4060 24546 4116 24556
rect 4172 22148 4228 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 15932 27186 15988 28028
rect 15932 27134 15934 27186
rect 15986 27134 15988 27186
rect 15932 27122 15988 27134
rect 16828 28082 17556 28084
rect 16828 28030 17502 28082
rect 17554 28030 17556 28082
rect 16828 28028 17556 28030
rect 14028 26290 14084 26302
rect 14028 26238 14030 26290
rect 14082 26238 14084 26290
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 13468 25618 13524 25630
rect 13468 25566 13470 25618
rect 13522 25566 13524 25618
rect 4284 25508 4340 25518
rect 4284 25414 4340 25452
rect 13468 25508 13524 25566
rect 13468 25442 13524 25452
rect 14028 25508 14084 26238
rect 14700 26180 14756 26190
rect 14700 26086 14756 26124
rect 16380 26180 16436 26190
rect 14028 25442 14084 25452
rect 15148 25508 15204 25518
rect 12908 25394 12964 25406
rect 12908 25342 12910 25394
rect 12962 25342 12964 25394
rect 12796 25282 12852 25294
rect 12796 25230 12798 25282
rect 12850 25230 12852 25282
rect 12796 24834 12852 25230
rect 12908 24948 12964 25342
rect 12908 24882 12964 24892
rect 13916 25396 13972 25406
rect 12796 24782 12798 24834
rect 12850 24782 12852 24834
rect 12796 24770 12852 24782
rect 12124 24722 12180 24734
rect 12124 24670 12126 24722
rect 12178 24670 12180 24722
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 12124 23492 12180 24670
rect 13916 24162 13972 25340
rect 13916 24110 13918 24162
rect 13970 24110 13972 24162
rect 13916 24098 13972 24110
rect 14476 25284 14532 25294
rect 14028 23828 14084 23838
rect 14252 23828 14308 23838
rect 14028 23826 14308 23828
rect 14028 23774 14030 23826
rect 14082 23774 14254 23826
rect 14306 23774 14308 23826
rect 14028 23772 14308 23774
rect 14028 23762 14084 23772
rect 14252 23762 14308 23772
rect 14476 23826 14532 25228
rect 14588 25060 14644 25070
rect 14588 23938 14644 25004
rect 14924 24612 14980 24622
rect 14924 24518 14980 24556
rect 14588 23886 14590 23938
rect 14642 23886 14644 23938
rect 14588 23874 14644 23886
rect 15148 24050 15204 25452
rect 16380 25508 16436 26124
rect 16828 26178 16884 28028
rect 17500 28018 17556 28028
rect 17612 31892 17780 31948
rect 17612 28084 17668 31892
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 21532 28644 21588 28654
rect 21420 28642 21588 28644
rect 21420 28590 21534 28642
rect 21586 28590 21588 28642
rect 21420 28588 21588 28590
rect 21308 28420 21364 28430
rect 20748 28418 21364 28420
rect 20748 28366 21310 28418
rect 21362 28366 21364 28418
rect 20748 28364 21364 28366
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 17612 28018 17668 28028
rect 20748 27970 20804 28364
rect 21308 28354 21364 28364
rect 20748 27918 20750 27970
rect 20802 27918 20804 27970
rect 20748 27906 20804 27918
rect 17276 27860 17332 27870
rect 16828 26126 16830 26178
rect 16882 26126 16884 26178
rect 16828 26114 16884 26126
rect 16940 27858 17332 27860
rect 16940 27806 17278 27858
rect 17330 27806 17332 27858
rect 16940 27804 17332 27806
rect 16604 26068 16660 26078
rect 16436 25452 16548 25508
rect 16380 25414 16436 25452
rect 15596 25396 15652 25406
rect 15596 25302 15652 25340
rect 15484 25060 15540 25070
rect 15484 24946 15540 25004
rect 15484 24894 15486 24946
rect 15538 24894 15540 24946
rect 15484 24882 15540 24894
rect 15596 24948 15652 24958
rect 16492 24948 16548 25452
rect 16604 25506 16660 26012
rect 16940 25956 16996 27804
rect 17276 27794 17332 27804
rect 17388 27860 17444 27870
rect 17612 27860 17668 27870
rect 16604 25454 16606 25506
rect 16658 25454 16660 25506
rect 16604 25442 16660 25454
rect 16828 25900 16996 25956
rect 17052 26964 17108 26974
rect 16828 25394 16884 25900
rect 16940 25508 16996 25518
rect 17052 25508 17108 26908
rect 16940 25506 17108 25508
rect 16940 25454 16942 25506
rect 16994 25454 17108 25506
rect 16940 25452 17108 25454
rect 17276 26066 17332 26078
rect 17276 26014 17278 26066
rect 17330 26014 17332 26066
rect 17276 25506 17332 26014
rect 17276 25454 17278 25506
rect 17330 25454 17332 25506
rect 16940 25442 16996 25452
rect 17276 25442 17332 25454
rect 16828 25342 16830 25394
rect 16882 25342 16884 25394
rect 16828 25330 16884 25342
rect 17388 25394 17444 27804
rect 17388 25342 17390 25394
rect 17442 25342 17444 25394
rect 17388 25330 17444 25342
rect 17500 27858 17668 27860
rect 17500 27806 17614 27858
rect 17666 27806 17668 27858
rect 17500 27804 17668 27806
rect 17500 26066 17556 27804
rect 17612 27794 17668 27804
rect 19964 27860 20020 27870
rect 18172 27076 18228 27086
rect 18060 26962 18116 26974
rect 18060 26910 18062 26962
rect 18114 26910 18116 26962
rect 17948 26404 18004 26414
rect 17948 26310 18004 26348
rect 17836 26292 17892 26302
rect 17724 26290 17892 26292
rect 17724 26238 17838 26290
rect 17890 26238 17892 26290
rect 17724 26236 17892 26238
rect 17612 26180 17668 26190
rect 17612 26086 17668 26124
rect 17500 26014 17502 26066
rect 17554 26014 17556 26066
rect 17500 25060 17556 26014
rect 17612 25508 17668 25518
rect 17724 25508 17780 26236
rect 17836 26226 17892 26236
rect 17948 26068 18004 26078
rect 18060 26068 18116 26910
rect 17948 26066 18116 26068
rect 17948 26014 17950 26066
rect 18002 26014 18116 26066
rect 17948 26012 18116 26014
rect 17948 26002 18004 26012
rect 17612 25506 17780 25508
rect 17612 25454 17614 25506
rect 17666 25454 17780 25506
rect 17612 25452 17780 25454
rect 17948 25508 18004 25518
rect 18172 25508 18228 27020
rect 18844 27076 18900 27086
rect 18844 26982 18900 27020
rect 19292 27076 19348 27086
rect 19292 26982 19348 27020
rect 19964 27076 20020 27804
rect 21420 27748 21476 28588
rect 21532 28578 21588 28588
rect 20748 27692 21476 27748
rect 20748 27298 20804 27692
rect 20748 27246 20750 27298
rect 20802 27246 20804 27298
rect 20748 27234 20804 27246
rect 19964 27010 20020 27020
rect 20188 27074 20244 27086
rect 20188 27022 20190 27074
rect 20242 27022 20244 27074
rect 18396 26964 18452 26974
rect 17948 25506 18228 25508
rect 17948 25454 17950 25506
rect 18002 25454 18228 25506
rect 17948 25452 18228 25454
rect 18284 26404 18340 26414
rect 17612 25442 17668 25452
rect 17948 25442 18004 25452
rect 16604 24948 16660 24958
rect 16492 24946 16660 24948
rect 16492 24894 16606 24946
rect 16658 24894 16660 24946
rect 16492 24892 16660 24894
rect 17500 24948 17556 25004
rect 17612 24948 17668 24958
rect 17500 24946 17668 24948
rect 17500 24894 17614 24946
rect 17666 24894 17668 24946
rect 17500 24892 17668 24894
rect 15596 24854 15652 24892
rect 16604 24882 16660 24892
rect 17612 24882 17668 24892
rect 15260 24724 15316 24734
rect 15260 24630 15316 24668
rect 15708 24722 15764 24734
rect 15708 24670 15710 24722
rect 15762 24670 15764 24722
rect 15148 23998 15150 24050
rect 15202 23998 15204 24050
rect 14476 23774 14478 23826
rect 14530 23774 14532 23826
rect 14476 23762 14532 23774
rect 13916 23716 13972 23726
rect 13804 23714 13972 23716
rect 13804 23662 13918 23714
rect 13970 23662 13972 23714
rect 13804 23660 13972 23662
rect 12348 23492 12404 23502
rect 12124 23436 12348 23492
rect 12348 23154 12404 23436
rect 12348 23102 12350 23154
rect 12402 23102 12404 23154
rect 12348 23090 12404 23102
rect 13020 23044 13076 23054
rect 13020 22950 13076 22988
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4172 22082 4228 22092
rect 13804 22146 13860 23660
rect 13916 23650 13972 23660
rect 14588 23604 14644 23614
rect 14140 23044 14196 23054
rect 14140 22482 14196 22988
rect 14140 22430 14142 22482
rect 14194 22430 14196 22482
rect 14140 22418 14196 22430
rect 13804 22094 13806 22146
rect 13858 22094 13860 22146
rect 13804 21700 13860 22094
rect 14028 22146 14084 22158
rect 14028 22094 14030 22146
rect 14082 22094 14084 22146
rect 13916 21700 13972 21710
rect 13804 21644 13916 21700
rect 13916 21634 13972 21644
rect 11004 21586 11060 21598
rect 11004 21534 11006 21586
rect 11058 21534 11060 21586
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 10780 19460 10836 19470
rect 10108 19348 10164 19358
rect 10108 19234 10164 19292
rect 10780 19346 10836 19404
rect 10780 19294 10782 19346
rect 10834 19294 10836 19346
rect 10780 19282 10836 19294
rect 11004 19348 11060 21534
rect 11788 21476 11844 21486
rect 13916 21476 13972 21486
rect 11788 21382 11844 21420
rect 13692 21474 13972 21476
rect 13692 21422 13918 21474
rect 13970 21422 13972 21474
rect 13692 21420 13972 21422
rect 13692 20356 13748 21420
rect 13916 21410 13972 21420
rect 14028 20804 14084 22094
rect 14028 20738 14084 20748
rect 14252 22146 14308 22158
rect 14252 22094 14254 22146
rect 14306 22094 14308 22146
rect 14252 21812 14308 22094
rect 14252 21362 14308 21756
rect 14476 21700 14532 21710
rect 14476 21606 14532 21644
rect 14364 21476 14420 21486
rect 14364 21382 14420 21420
rect 14252 21310 14254 21362
rect 14306 21310 14308 21362
rect 14140 20580 14196 20590
rect 13692 20290 13748 20300
rect 13804 20578 14196 20580
rect 13804 20526 14142 20578
rect 14194 20526 14196 20578
rect 13804 20524 14196 20526
rect 13132 19908 13188 19918
rect 11004 19282 11060 19292
rect 12908 19348 12964 19358
rect 13132 19348 13188 19852
rect 12908 19346 13188 19348
rect 12908 19294 12910 19346
rect 12962 19294 13188 19346
rect 12908 19292 13188 19294
rect 13356 19906 13412 19918
rect 13356 19854 13358 19906
rect 13410 19854 13412 19906
rect 13356 19460 13412 19854
rect 13804 19908 13860 20524
rect 14140 20514 14196 20524
rect 14028 20356 14084 20366
rect 14028 20018 14084 20300
rect 14028 19966 14030 20018
rect 14082 19966 14084 20018
rect 14028 19954 14084 19966
rect 13804 19814 13860 19852
rect 12908 19282 12964 19292
rect 10108 19182 10110 19234
rect 10162 19182 10164 19234
rect 10108 19170 10164 19182
rect 13356 18788 13412 19404
rect 14140 19796 14196 19806
rect 13356 18722 13412 18732
rect 13580 19348 13636 19358
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 13580 17666 13636 19292
rect 14140 19236 14196 19740
rect 14140 19142 14196 19180
rect 14252 19124 14308 21310
rect 14476 20692 14532 20702
rect 14588 20692 14644 23548
rect 15148 23492 15204 23998
rect 15708 23604 15764 24670
rect 15708 23538 15764 23548
rect 15932 24722 15988 24734
rect 15932 24670 15934 24722
rect 15986 24670 15988 24722
rect 15204 23436 15652 23492
rect 15148 23426 15204 23436
rect 15148 23042 15204 23054
rect 15148 22990 15150 23042
rect 15202 22990 15204 23042
rect 15148 22484 15204 22990
rect 15148 22418 15204 22428
rect 14700 22146 14756 22158
rect 14700 22094 14702 22146
rect 14754 22094 14756 22146
rect 14700 22036 14756 22094
rect 14700 21970 14756 21980
rect 15260 22036 15316 23436
rect 15596 23378 15652 23436
rect 15596 23326 15598 23378
rect 15650 23326 15652 23378
rect 15596 23314 15652 23326
rect 15932 23380 15988 24670
rect 17836 24722 17892 24734
rect 17836 24670 17838 24722
rect 17890 24670 17892 24722
rect 17836 23492 17892 24670
rect 17836 23426 17892 23436
rect 18172 23828 18228 23838
rect 15932 23314 15988 23324
rect 17388 23380 17444 23390
rect 17388 23286 17444 23324
rect 15484 23268 15540 23278
rect 15148 21924 15204 21934
rect 15036 21812 15092 21822
rect 15036 21718 15092 21756
rect 15148 21698 15204 21868
rect 15148 21646 15150 21698
rect 15202 21646 15204 21698
rect 15148 21634 15204 21646
rect 14812 21588 14868 21598
rect 14812 21494 14868 21532
rect 15260 20916 15316 21980
rect 14476 20690 14644 20692
rect 14476 20638 14478 20690
rect 14530 20638 14644 20690
rect 14476 20636 14644 20638
rect 15148 20914 15316 20916
rect 15148 20862 15262 20914
rect 15314 20862 15316 20914
rect 15148 20860 15316 20862
rect 14476 20626 14532 20636
rect 14364 19796 14420 19806
rect 14364 19702 14420 19740
rect 15148 19348 15204 20860
rect 15260 20850 15316 20860
rect 15372 22260 15428 22270
rect 15372 20692 15428 22204
rect 15260 20636 15428 20692
rect 15260 20130 15316 20636
rect 15260 20078 15262 20130
rect 15314 20078 15316 20130
rect 15260 20066 15316 20078
rect 15372 20132 15428 20142
rect 15484 20132 15540 23212
rect 17948 23268 18004 23278
rect 17948 23174 18004 23212
rect 17836 23156 17892 23166
rect 17612 23100 17836 23156
rect 16044 22484 16100 22494
rect 16268 22484 16324 22494
rect 16100 22482 16324 22484
rect 16100 22430 16270 22482
rect 16322 22430 16324 22482
rect 16100 22428 16324 22430
rect 15932 21924 15988 21934
rect 15820 21868 15932 21924
rect 15372 20130 15540 20132
rect 15372 20078 15374 20130
rect 15426 20078 15540 20130
rect 15372 20076 15540 20078
rect 15596 20580 15652 20590
rect 15372 20066 15428 20076
rect 15596 20020 15652 20524
rect 15484 19964 15652 20020
rect 15372 19796 15428 19806
rect 15372 19702 15428 19740
rect 14364 19124 14420 19134
rect 14252 19122 14756 19124
rect 14252 19070 14366 19122
rect 14418 19070 14756 19122
rect 14252 19068 14756 19070
rect 14364 19058 14420 19068
rect 14476 18452 14532 18462
rect 14476 18358 14532 18396
rect 14700 18450 14756 19068
rect 15148 18564 15204 19292
rect 15372 19236 15428 19246
rect 15372 19142 15428 19180
rect 15148 18498 15204 18508
rect 14700 18398 14702 18450
rect 14754 18398 14756 18450
rect 14700 18386 14756 18398
rect 15036 18450 15092 18462
rect 15036 18398 15038 18450
rect 15090 18398 15092 18450
rect 14588 18338 14644 18350
rect 14588 18286 14590 18338
rect 14642 18286 14644 18338
rect 14252 17780 14308 17790
rect 14588 17780 14644 18286
rect 15036 18116 15092 18398
rect 15036 18050 15092 18060
rect 14252 17778 14644 17780
rect 14252 17726 14254 17778
rect 14306 17726 14644 17778
rect 14252 17724 14644 17726
rect 14252 17714 14308 17724
rect 13580 17614 13582 17666
rect 13634 17614 13636 17666
rect 13580 17602 13636 17614
rect 15148 16996 15204 17006
rect 15484 16996 15540 19964
rect 15820 19906 15876 21868
rect 15932 21858 15988 21868
rect 15932 21588 15988 21598
rect 16044 21588 16100 22428
rect 16268 22418 16324 22428
rect 17388 22370 17444 22382
rect 17388 22318 17390 22370
rect 17442 22318 17444 22370
rect 16380 22260 16436 22270
rect 16380 22166 16436 22204
rect 17052 22148 17108 22158
rect 17052 22054 17108 22092
rect 16940 22036 16996 22046
rect 15932 21586 16100 21588
rect 15932 21534 15934 21586
rect 15986 21534 16100 21586
rect 15932 21532 16100 21534
rect 16156 21698 16212 21710
rect 16156 21646 16158 21698
rect 16210 21646 16212 21698
rect 15932 21522 15988 21532
rect 15820 19854 15822 19906
rect 15874 19854 15876 19906
rect 15820 19842 15876 19854
rect 15932 20130 15988 20142
rect 15932 20078 15934 20130
rect 15986 20078 15988 20130
rect 15820 19236 15876 19246
rect 15932 19236 15988 20078
rect 16156 20132 16212 21646
rect 16828 21700 16884 21710
rect 16940 21700 16996 21980
rect 17388 21924 17444 22318
rect 17388 21858 17444 21868
rect 17500 22260 17556 22270
rect 17612 22260 17668 23100
rect 17836 23062 17892 23100
rect 18060 23154 18116 23166
rect 18060 23102 18062 23154
rect 18114 23102 18116 23154
rect 18060 22484 18116 23102
rect 17836 22428 18060 22484
rect 17556 22204 17668 22260
rect 17724 22260 17780 22270
rect 17836 22260 17892 22428
rect 18060 22418 18116 22428
rect 17724 22258 17892 22260
rect 17724 22206 17726 22258
rect 17778 22206 17892 22258
rect 17724 22204 17892 22206
rect 18060 22258 18116 22270
rect 18060 22206 18062 22258
rect 18114 22206 18116 22258
rect 16828 21698 16996 21700
rect 16828 21646 16830 21698
rect 16882 21646 16996 21698
rect 16828 21644 16996 21646
rect 16828 21634 16884 21644
rect 16604 21588 16660 21598
rect 16604 20356 16660 21532
rect 16604 20290 16660 20300
rect 16492 20132 16548 20142
rect 16156 20130 16660 20132
rect 16156 20078 16158 20130
rect 16210 20078 16494 20130
rect 16546 20078 16660 20130
rect 16156 20076 16660 20078
rect 16156 20066 16212 20076
rect 16492 20066 16548 20076
rect 16604 20020 16660 20076
rect 16492 19236 16548 19246
rect 15820 19234 15988 19236
rect 15820 19182 15822 19234
rect 15874 19182 15988 19234
rect 15820 19180 15988 19182
rect 16156 19180 16492 19236
rect 15820 18788 15876 19180
rect 15820 18722 15876 18732
rect 15932 19010 15988 19022
rect 15932 18958 15934 19010
rect 15986 18958 15988 19010
rect 15932 18340 15988 18958
rect 16156 18562 16212 19180
rect 16156 18510 16158 18562
rect 16210 18510 16212 18562
rect 16156 18498 16212 18510
rect 15988 18284 16212 18340
rect 15932 18274 15988 18284
rect 15148 16994 15540 16996
rect 15148 16942 15150 16994
rect 15202 16942 15540 16994
rect 15148 16940 15540 16942
rect 15596 17444 15652 17454
rect 15148 16930 15204 16940
rect 4284 16884 4340 16894
rect 4284 16790 4340 16828
rect 12124 16884 12180 16894
rect 1932 16658 1988 16670
rect 1932 16606 1934 16658
rect 1986 16606 1988 16658
rect 1932 16212 1988 16606
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 1932 16146 1988 16156
rect 12124 15202 12180 16828
rect 14812 16884 14868 16894
rect 14812 16790 14868 16828
rect 15036 16770 15092 16782
rect 15036 16718 15038 16770
rect 15090 16718 15092 16770
rect 15036 16100 15092 16718
rect 15596 16322 15652 17388
rect 16156 17332 16212 18284
rect 16268 18226 16324 18238
rect 16268 18174 16270 18226
rect 16322 18174 16324 18226
rect 16268 17668 16324 18174
rect 16380 17778 16436 19180
rect 16492 19142 16548 19180
rect 16604 18562 16660 19964
rect 16828 20130 16884 20142
rect 16828 20078 16830 20130
rect 16882 20078 16884 20130
rect 16828 19460 16884 20078
rect 16940 19460 16996 21644
rect 17500 21586 17556 22204
rect 17612 22036 17668 22046
rect 17724 22036 17780 22204
rect 17668 21980 17780 22036
rect 17612 21970 17668 21980
rect 17500 21534 17502 21586
rect 17554 21534 17556 21586
rect 17500 21522 17556 21534
rect 17836 21474 17892 21486
rect 17836 21422 17838 21474
rect 17890 21422 17892 21474
rect 17836 20580 17892 21422
rect 17836 20514 17892 20524
rect 17276 20018 17332 20030
rect 17276 19966 17278 20018
rect 17330 19966 17332 20018
rect 17164 19460 17220 19470
rect 16940 19458 17220 19460
rect 16940 19406 17166 19458
rect 17218 19406 17220 19458
rect 16940 19404 17220 19406
rect 16828 19394 16884 19404
rect 17164 19394 17220 19404
rect 17276 19236 17332 19966
rect 17948 20020 18004 20030
rect 17948 19906 18004 19964
rect 17948 19854 17950 19906
rect 18002 19854 18004 19906
rect 17948 19842 18004 19854
rect 17276 19170 17332 19180
rect 17724 19796 17780 19806
rect 16716 19010 16772 19022
rect 16716 18958 16718 19010
rect 16770 18958 16772 19010
rect 16716 18788 16772 18958
rect 17276 19012 17332 19022
rect 17276 18918 17332 18956
rect 17388 19010 17444 19022
rect 17388 18958 17390 19010
rect 17442 18958 17444 19010
rect 17388 18900 17444 18958
rect 17388 18834 17444 18844
rect 16716 18722 16772 18732
rect 16604 18510 16606 18562
rect 16658 18510 16660 18562
rect 16604 18498 16660 18510
rect 16716 18564 16772 18574
rect 17052 18564 17108 18574
rect 16716 18562 17052 18564
rect 16716 18510 16718 18562
rect 16770 18510 17052 18562
rect 16716 18508 17052 18510
rect 16716 18498 16772 18508
rect 17052 18498 17108 18508
rect 17724 18562 17780 19740
rect 17836 19460 17892 19470
rect 17836 19366 17892 19404
rect 18060 18900 18116 22206
rect 18172 20130 18228 23772
rect 18284 21476 18340 26348
rect 18396 22146 18452 26908
rect 20188 26908 20244 27022
rect 20412 27076 20468 27086
rect 21420 27076 21476 27086
rect 20412 27074 21476 27076
rect 20412 27022 20414 27074
rect 20466 27022 21422 27074
rect 21474 27022 21476 27074
rect 20412 27020 21476 27022
rect 20412 27010 20468 27020
rect 21420 27010 21476 27020
rect 21644 26908 21700 37212
rect 21980 27860 22036 27870
rect 23436 27860 23492 27870
rect 22036 27804 22148 27860
rect 21980 27794 22036 27804
rect 21756 27076 21812 27086
rect 21756 26982 21812 27020
rect 21980 26964 22036 26974
rect 20188 26852 20468 26908
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20412 26292 20468 26852
rect 18620 25396 18676 25406
rect 18620 25394 19684 25396
rect 18620 25342 18622 25394
rect 18674 25342 19684 25394
rect 18620 25340 19684 25342
rect 18620 25330 18676 25340
rect 19628 24948 19684 25340
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19964 24948 20020 24958
rect 19628 24946 20020 24948
rect 19628 24894 19966 24946
rect 20018 24894 20020 24946
rect 19628 24892 20020 24894
rect 19964 24882 20020 24892
rect 19852 24724 19908 24734
rect 19852 24630 19908 24668
rect 20076 24722 20132 24734
rect 20076 24670 20078 24722
rect 20130 24670 20132 24722
rect 20076 23716 20132 24670
rect 20412 24724 20468 26236
rect 21420 26852 21700 26908
rect 21868 26962 22036 26964
rect 21868 26910 21982 26962
rect 22034 26910 22036 26962
rect 21868 26908 22036 26910
rect 20748 25620 20804 25630
rect 21420 25620 21476 26852
rect 20748 25618 21476 25620
rect 20748 25566 20750 25618
rect 20802 25566 21476 25618
rect 20748 25564 21476 25566
rect 20748 25554 20804 25564
rect 21420 25394 21476 25564
rect 21420 25342 21422 25394
rect 21474 25342 21476 25394
rect 21420 25330 21476 25342
rect 21532 25394 21588 25406
rect 21532 25342 21534 25394
rect 21586 25342 21588 25394
rect 21196 25284 21252 25294
rect 20300 23716 20356 23726
rect 19628 23660 20132 23716
rect 20188 23660 20300 23716
rect 19068 23604 19124 23614
rect 18844 23492 18900 23502
rect 18732 23266 18788 23278
rect 18732 23214 18734 23266
rect 18786 23214 18788 23266
rect 18508 23156 18564 23166
rect 18508 23062 18564 23100
rect 18396 22094 18398 22146
rect 18450 22094 18452 22146
rect 18396 21812 18452 22094
rect 18396 21746 18452 21756
rect 18508 22148 18564 22158
rect 18284 21410 18340 21420
rect 18396 21588 18452 21598
rect 18172 20078 18174 20130
rect 18226 20078 18228 20130
rect 18172 20066 18228 20078
rect 18284 20132 18340 20142
rect 18172 19460 18228 19470
rect 18172 19366 18228 19404
rect 18060 18834 18116 18844
rect 18172 19236 18228 19246
rect 18284 19236 18340 20076
rect 18172 19234 18340 19236
rect 18172 19182 18174 19234
rect 18226 19182 18340 19234
rect 18172 19180 18340 19182
rect 18396 20018 18452 21532
rect 18508 21586 18564 22092
rect 18508 21534 18510 21586
rect 18562 21534 18564 21586
rect 18508 21522 18564 21534
rect 18732 20132 18788 23214
rect 18844 23156 18900 23436
rect 18844 23042 18900 23100
rect 18844 22990 18846 23042
rect 18898 22990 18900 23042
rect 18844 22978 18900 22990
rect 18844 22484 18900 22494
rect 18844 22370 18900 22428
rect 18844 22318 18846 22370
rect 18898 22318 18900 22370
rect 18844 22306 18900 22318
rect 19068 22370 19124 23548
rect 19628 23604 19684 23660
rect 19628 23380 19684 23548
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19740 23380 19796 23390
rect 19628 23378 19796 23380
rect 19628 23326 19742 23378
rect 19794 23326 19796 23378
rect 19628 23324 19796 23326
rect 19740 23314 19796 23324
rect 19964 23380 20020 23390
rect 19516 23268 19572 23278
rect 19572 23212 19684 23268
rect 19516 23174 19572 23212
rect 19068 22318 19070 22370
rect 19122 22318 19124 22370
rect 19068 22306 19124 22318
rect 18956 22146 19012 22158
rect 18956 22094 18958 22146
rect 19010 22094 19012 22146
rect 18956 21700 19012 22094
rect 19012 21644 19124 21700
rect 18956 21634 19012 21644
rect 18732 20066 18788 20076
rect 18396 19966 18398 20018
rect 18450 19966 18452 20018
rect 18396 19236 18452 19966
rect 19068 20020 19124 21644
rect 19180 21476 19236 21486
rect 19180 20692 19236 21420
rect 19180 20242 19236 20636
rect 19180 20190 19182 20242
rect 19234 20190 19236 20242
rect 19180 20178 19236 20190
rect 19292 20132 19348 20142
rect 19292 20038 19348 20076
rect 19068 19926 19124 19964
rect 19404 19572 19460 19582
rect 19460 19516 19572 19572
rect 19404 19506 19460 19516
rect 18508 19236 18564 19246
rect 18396 19234 18564 19236
rect 18396 19182 18510 19234
rect 18562 19182 18564 19234
rect 18396 19180 18564 19182
rect 18172 18676 18228 19180
rect 18508 19170 18564 19180
rect 18844 19236 18900 19246
rect 18844 19122 18900 19180
rect 18844 19070 18846 19122
rect 18898 19070 18900 19122
rect 18844 19058 18900 19070
rect 19292 19234 19348 19246
rect 19292 19182 19294 19234
rect 19346 19182 19348 19234
rect 19292 18900 19348 19182
rect 19292 18834 19348 18844
rect 19404 19122 19460 19134
rect 19404 19070 19406 19122
rect 19458 19070 19460 19122
rect 18844 18788 18900 18798
rect 17724 18510 17726 18562
rect 17778 18510 17780 18562
rect 16492 18452 16548 18462
rect 16492 18228 16548 18396
rect 17164 18452 17220 18462
rect 17220 18396 17332 18452
rect 17164 18386 17220 18396
rect 16716 18228 16772 18238
rect 16492 18172 16716 18228
rect 16772 18172 16996 18228
rect 16716 18134 16772 18172
rect 16380 17726 16382 17778
rect 16434 17726 16436 17778
rect 16380 17714 16436 17726
rect 16268 17602 16324 17612
rect 16940 17666 16996 18172
rect 17164 17892 17220 17902
rect 16940 17614 16942 17666
rect 16994 17614 16996 17666
rect 16940 17602 16996 17614
rect 17052 17890 17220 17892
rect 17052 17838 17166 17890
rect 17218 17838 17220 17890
rect 17052 17836 17220 17838
rect 16604 17444 16660 17454
rect 16604 17350 16660 17388
rect 16828 17444 16884 17454
rect 17052 17444 17108 17836
rect 17164 17826 17220 17836
rect 16828 17442 17108 17444
rect 16828 17390 16830 17442
rect 16882 17390 17108 17442
rect 16828 17388 17108 17390
rect 17276 17780 17332 18396
rect 17388 18450 17444 18462
rect 17388 18398 17390 18450
rect 17442 18398 17444 18450
rect 17388 18228 17444 18398
rect 17388 18162 17444 18172
rect 17724 17890 17780 18510
rect 17724 17838 17726 17890
rect 17778 17838 17780 17890
rect 17724 17826 17780 17838
rect 17948 18620 18228 18676
rect 18396 18674 18452 18686
rect 18396 18622 18398 18674
rect 18450 18622 18452 18674
rect 17948 18564 18004 18620
rect 17388 17780 17444 17790
rect 17276 17778 17444 17780
rect 17276 17726 17390 17778
rect 17442 17726 17444 17778
rect 17276 17724 17444 17726
rect 16828 17378 16884 17388
rect 16156 17276 16436 17332
rect 15596 16270 15598 16322
rect 15650 16270 15652 16322
rect 15596 16258 15652 16270
rect 15148 16100 15204 16110
rect 15036 16098 15204 16100
rect 15036 16046 15150 16098
rect 15202 16046 15204 16098
rect 15036 16044 15204 16046
rect 15148 16034 15204 16044
rect 15372 16100 15428 16110
rect 15372 16006 15428 16044
rect 14252 15876 14308 15886
rect 14252 15426 14308 15820
rect 15260 15876 15316 15886
rect 15260 15782 15316 15820
rect 14252 15374 14254 15426
rect 14306 15374 14308 15426
rect 14252 15362 14308 15374
rect 14364 15540 14420 15550
rect 12124 15150 12126 15202
rect 12178 15150 12180 15202
rect 12124 15138 12180 15150
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 14252 14532 14308 14542
rect 14364 14532 14420 15484
rect 15036 15540 15092 15550
rect 15036 15314 15092 15484
rect 15484 15540 15540 15550
rect 15484 15446 15540 15484
rect 16380 15538 16436 17276
rect 16380 15486 16382 15538
rect 16434 15486 16436 15538
rect 16380 15474 16436 15486
rect 17276 15540 17332 17724
rect 17388 17714 17444 17724
rect 17948 17554 18004 18508
rect 18396 18564 18452 18622
rect 18844 18674 18900 18732
rect 18844 18622 18846 18674
rect 18898 18622 18900 18674
rect 18844 18610 18900 18622
rect 19180 18676 19236 18686
rect 18396 18498 18452 18508
rect 18284 18450 18340 18462
rect 18284 18398 18286 18450
rect 18338 18398 18340 18450
rect 18284 18340 18340 18398
rect 19180 18450 19236 18620
rect 19180 18398 19182 18450
rect 19234 18398 19236 18450
rect 19180 18386 19236 18398
rect 18284 18274 18340 18284
rect 18172 17668 18228 17678
rect 19404 17668 19460 19070
rect 18228 17612 18340 17668
rect 18172 17574 18228 17612
rect 17948 17502 17950 17554
rect 18002 17502 18004 17554
rect 17948 17490 18004 17502
rect 18284 17106 18340 17612
rect 18284 17054 18286 17106
rect 18338 17054 18340 17106
rect 18284 17042 18340 17054
rect 18620 17612 19460 17668
rect 19516 17666 19572 19516
rect 19628 18788 19684 23212
rect 19852 22930 19908 22942
rect 19852 22878 19854 22930
rect 19906 22878 19908 22930
rect 19852 22260 19908 22878
rect 19964 22370 20020 23324
rect 20188 22594 20244 23660
rect 20300 23650 20356 23660
rect 20300 23380 20356 23390
rect 20300 23154 20356 23324
rect 20300 23102 20302 23154
rect 20354 23102 20356 23154
rect 20300 23090 20356 23102
rect 20188 22542 20190 22594
rect 20242 22542 20244 22594
rect 20188 22530 20244 22542
rect 19964 22318 19966 22370
rect 20018 22318 20020 22370
rect 19964 22306 20020 22318
rect 19852 22194 19908 22204
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20076 21700 20132 21710
rect 20076 20802 20132 21644
rect 20412 21028 20468 24668
rect 20524 25282 21252 25284
rect 20524 25230 21198 25282
rect 21250 25230 21252 25282
rect 20524 25228 21252 25230
rect 20524 24722 20580 25228
rect 21196 25218 21252 25228
rect 20524 24670 20526 24722
rect 20578 24670 20580 24722
rect 20524 24658 20580 24670
rect 21532 23492 21588 25342
rect 21868 25284 21924 26908
rect 21980 26898 22036 26908
rect 21980 25620 22036 25630
rect 22092 25620 22148 27804
rect 22428 27748 22484 27758
rect 22428 26962 22484 27692
rect 22876 27748 22932 27758
rect 22876 27654 22932 27692
rect 23436 27076 23492 27804
rect 23548 27076 23604 27086
rect 23436 27074 23604 27076
rect 23436 27022 23550 27074
rect 23602 27022 23604 27074
rect 23436 27020 23604 27022
rect 22428 26910 22430 26962
rect 22482 26910 22484 26962
rect 22428 26898 22484 26910
rect 23548 26908 23604 27020
rect 23436 26852 23604 26908
rect 23436 26786 23492 26796
rect 21980 25618 22148 25620
rect 21980 25566 21982 25618
rect 22034 25566 22148 25618
rect 21980 25564 22148 25566
rect 21980 25554 22036 25564
rect 23436 25396 23492 25406
rect 23436 25284 23492 25340
rect 21868 23828 21924 25228
rect 23324 25282 23492 25284
rect 23324 25230 23438 25282
rect 23490 25230 23492 25282
rect 23324 25228 23492 25230
rect 22316 23940 22372 23950
rect 22316 23846 22372 23884
rect 23100 23940 23156 23950
rect 21980 23828 22036 23838
rect 21868 23772 21980 23828
rect 21980 23734 22036 23772
rect 22092 23716 22148 23726
rect 22092 23622 22148 23660
rect 22652 23714 22708 23726
rect 22652 23662 22654 23714
rect 22706 23662 22708 23714
rect 21532 23156 21588 23436
rect 22652 23268 22708 23662
rect 22652 23202 22708 23212
rect 22988 23714 23044 23726
rect 22988 23662 22990 23714
rect 23042 23662 23044 23714
rect 21532 23090 21588 23100
rect 20972 23042 21028 23054
rect 20972 22990 20974 23042
rect 21026 22990 21028 23042
rect 20636 22484 20692 22494
rect 20972 22484 21028 22990
rect 20636 22482 21028 22484
rect 20636 22430 20638 22482
rect 20690 22430 21028 22482
rect 20636 22428 21028 22430
rect 20636 22418 20692 22428
rect 21868 22370 21924 22382
rect 21868 22318 21870 22370
rect 21922 22318 21924 22370
rect 20524 22260 20580 22270
rect 20524 22166 20580 22204
rect 20748 22260 20804 22270
rect 20748 22258 21476 22260
rect 20748 22206 20750 22258
rect 20802 22206 21476 22258
rect 20748 22204 21476 22206
rect 20748 22194 20804 22204
rect 20636 21028 20692 21038
rect 20412 21026 20692 21028
rect 20412 20974 20638 21026
rect 20690 20974 20692 21026
rect 20412 20972 20692 20974
rect 20636 20962 20692 20972
rect 21420 21026 21476 22204
rect 21868 21700 21924 22318
rect 22988 22148 23044 23662
rect 23100 23042 23156 23884
rect 23100 22990 23102 23042
rect 23154 22990 23156 23042
rect 23100 22978 23156 22990
rect 22876 22092 22988 22148
rect 21868 21606 21924 21644
rect 22092 21812 22148 21822
rect 21420 20974 21422 21026
rect 21474 20974 21476 21026
rect 21420 20962 21476 20974
rect 20076 20750 20078 20802
rect 20130 20750 20132 20802
rect 20076 20738 20132 20750
rect 22092 20802 22148 21756
rect 22764 21812 22820 21822
rect 22092 20750 22094 20802
rect 22146 20750 22148 20802
rect 22092 20738 22148 20750
rect 22204 20914 22260 20926
rect 22204 20862 22206 20914
rect 22258 20862 22260 20914
rect 20524 20692 20580 20702
rect 20412 20690 20580 20692
rect 20412 20638 20526 20690
rect 20578 20638 20580 20690
rect 20412 20636 20580 20638
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19852 20130 19908 20142
rect 19852 20078 19854 20130
rect 19906 20078 19908 20130
rect 19852 19572 19908 20078
rect 19852 19506 19908 19516
rect 20412 19460 20468 20636
rect 20524 20626 20580 20636
rect 21308 20690 21364 20702
rect 21308 20638 21310 20690
rect 21362 20638 21364 20690
rect 20636 20580 20692 20590
rect 20860 20580 20916 20590
rect 20636 20578 20804 20580
rect 20636 20526 20638 20578
rect 20690 20526 20804 20578
rect 20636 20524 20804 20526
rect 20636 20514 20692 20524
rect 20524 20020 20580 20030
rect 20524 19926 20580 19964
rect 20076 19236 20132 19246
rect 20076 19142 20132 19180
rect 20300 19012 20356 19022
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 18450 19684 18732
rect 19628 18398 19630 18450
rect 19682 18398 19684 18450
rect 19628 18386 19684 18398
rect 19964 18562 20020 18574
rect 20300 18564 20356 18956
rect 20412 18674 20468 19404
rect 20524 19572 20580 19582
rect 20524 19234 20580 19516
rect 20524 19182 20526 19234
rect 20578 19182 20580 19234
rect 20524 19170 20580 19182
rect 20636 19236 20692 19246
rect 20748 19236 20804 20524
rect 20860 20130 20916 20524
rect 21308 20580 21364 20638
rect 21868 20692 21924 20702
rect 21868 20598 21924 20636
rect 21308 20514 21364 20524
rect 21420 20578 21476 20590
rect 21420 20526 21422 20578
rect 21474 20526 21476 20578
rect 20860 20078 20862 20130
rect 20914 20078 20916 20130
rect 20860 20066 20916 20078
rect 20972 20244 21028 20254
rect 20692 19180 20804 19236
rect 20972 19906 21028 20188
rect 20972 19854 20974 19906
rect 21026 19854 21028 19906
rect 20636 19170 20692 19180
rect 20860 19124 20916 19134
rect 20860 19030 20916 19068
rect 20412 18622 20414 18674
rect 20466 18622 20468 18674
rect 20412 18610 20468 18622
rect 19964 18510 19966 18562
rect 20018 18510 20020 18562
rect 19852 17780 19908 17790
rect 19516 17614 19518 17666
rect 19570 17614 19572 17666
rect 18620 17106 18676 17612
rect 18620 17054 18622 17106
rect 18674 17054 18676 17106
rect 18620 17042 18676 17054
rect 18620 16212 18676 16222
rect 18508 16210 18676 16212
rect 18508 16158 18622 16210
rect 18674 16158 18676 16210
rect 18508 16156 18676 16158
rect 17500 15540 17556 15550
rect 17332 15538 17556 15540
rect 17332 15486 17502 15538
rect 17554 15486 17556 15538
rect 17332 15484 17556 15486
rect 17276 15474 17332 15484
rect 15036 15262 15038 15314
rect 15090 15262 15092 15314
rect 15036 15250 15092 15262
rect 14924 15204 14980 15214
rect 14924 14642 14980 15148
rect 16268 15204 16324 15242
rect 16268 15138 16324 15148
rect 16604 15204 16660 15242
rect 16604 15138 16660 15148
rect 17276 15090 17332 15102
rect 17276 15038 17278 15090
rect 17330 15038 17332 15090
rect 14924 14590 14926 14642
rect 14978 14590 14980 14642
rect 14924 14578 14980 14590
rect 17052 14644 17108 14654
rect 17276 14644 17332 15038
rect 17052 14642 17332 14644
rect 17052 14590 17054 14642
rect 17106 14590 17332 14642
rect 17052 14588 17332 14590
rect 14252 14530 14420 14532
rect 14252 14478 14254 14530
rect 14306 14478 14420 14530
rect 14252 14476 14420 14478
rect 14252 14466 14308 14476
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 17052 8428 17108 14588
rect 17388 14532 17444 15484
rect 17500 15474 17556 15484
rect 18060 15484 18452 15540
rect 17948 15092 18004 15102
rect 18060 15092 18116 15484
rect 18172 15316 18228 15326
rect 18172 15222 18228 15260
rect 18396 15314 18452 15484
rect 18396 15262 18398 15314
rect 18450 15262 18452 15314
rect 18396 15250 18452 15262
rect 18284 15204 18340 15242
rect 18284 15138 18340 15148
rect 18508 15092 18564 16156
rect 18620 16146 18676 16156
rect 18732 16100 18788 16110
rect 18732 15986 18788 16044
rect 18732 15934 18734 15986
rect 18786 15934 18788 15986
rect 18732 15922 18788 15934
rect 18620 15540 18676 15550
rect 18844 15540 18900 17612
rect 19516 17602 19572 17614
rect 19628 17778 19908 17780
rect 19628 17726 19854 17778
rect 19906 17726 19908 17778
rect 19628 17724 19908 17726
rect 19180 17444 19236 17454
rect 19236 17388 19460 17444
rect 19180 17350 19236 17388
rect 18956 15988 19012 15998
rect 18956 15986 19236 15988
rect 18956 15934 18958 15986
rect 19010 15934 19236 15986
rect 18956 15932 19236 15934
rect 18956 15922 19012 15932
rect 19068 15540 19124 15550
rect 18844 15538 19124 15540
rect 18844 15486 19070 15538
rect 19122 15486 19124 15538
rect 18844 15484 19124 15486
rect 18620 15446 18676 15484
rect 19068 15428 19124 15484
rect 19180 15538 19236 15932
rect 19180 15486 19182 15538
rect 19234 15486 19236 15538
rect 19180 15474 19236 15486
rect 19404 15540 19460 17388
rect 19628 16100 19684 17724
rect 19852 17714 19908 17724
rect 19964 17668 20020 18510
rect 20188 18562 20356 18564
rect 20188 18510 20302 18562
rect 20354 18510 20356 18562
rect 20188 18508 20356 18510
rect 20188 17890 20244 18508
rect 20300 18498 20356 18508
rect 20412 18228 20468 18238
rect 20412 18134 20468 18172
rect 20972 18004 21028 19854
rect 21420 19236 21476 20526
rect 21420 19170 21476 19180
rect 21756 19236 21812 19246
rect 20188 17838 20190 17890
rect 20242 17838 20244 17890
rect 20188 17826 20244 17838
rect 20300 17948 21028 18004
rect 21420 18450 21476 18462
rect 21420 18398 21422 18450
rect 21474 18398 21476 18450
rect 19964 17554 20020 17612
rect 19964 17502 19966 17554
rect 20018 17502 20020 17554
rect 19964 17490 20020 17502
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 16034 19684 16044
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19516 15540 19572 15550
rect 19460 15538 19572 15540
rect 19460 15486 19518 15538
rect 19570 15486 19572 15538
rect 19460 15484 19572 15486
rect 19404 15446 19460 15484
rect 19516 15474 19572 15484
rect 19068 15362 19124 15372
rect 19964 15428 20020 15438
rect 19964 15334 20020 15372
rect 17948 15090 18116 15092
rect 17948 15038 17950 15090
rect 18002 15038 18116 15090
rect 17948 15036 18116 15038
rect 18396 15036 18564 15092
rect 19292 15314 19348 15326
rect 19292 15262 19294 15314
rect 19346 15262 19348 15314
rect 17948 15026 18004 15036
rect 18396 14980 18452 15036
rect 18172 14924 18452 14980
rect 18172 14642 18228 14924
rect 18172 14590 18174 14642
rect 18226 14590 18228 14642
rect 18172 14578 18228 14590
rect 19292 14644 19348 15262
rect 20300 15314 20356 17948
rect 21084 17444 21140 17454
rect 20972 15428 21028 15438
rect 20972 15334 21028 15372
rect 21084 15426 21140 17388
rect 21420 16884 21476 18398
rect 21756 17554 21812 19180
rect 22204 19234 22260 20862
rect 22428 20804 22484 20814
rect 22428 20710 22484 20748
rect 22764 20802 22820 21756
rect 22764 20750 22766 20802
rect 22818 20750 22820 20802
rect 22764 20738 22820 20750
rect 22876 20580 22932 22092
rect 22988 22082 23044 22092
rect 23324 20804 23380 25228
rect 23436 25218 23492 25228
rect 23660 23940 23716 37998
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 24332 27972 24388 27982
rect 24332 27186 24388 27916
rect 24556 27748 24612 37998
rect 26236 37492 26292 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 26236 37426 26292 37436
rect 27468 37492 27524 37502
rect 27468 37398 27524 37436
rect 26460 37266 26516 37278
rect 26460 37214 26462 37266
rect 26514 37214 26516 37266
rect 25228 27972 25284 27982
rect 25228 27878 25284 27916
rect 24556 27682 24612 27692
rect 24668 27860 24724 27870
rect 24332 27134 24334 27186
rect 24386 27134 24388 27186
rect 24332 27122 24388 27134
rect 24668 26514 24724 27804
rect 25452 27860 25508 27870
rect 25452 27766 25508 27804
rect 24668 26462 24670 26514
rect 24722 26462 24724 26514
rect 24668 26450 24724 26462
rect 24892 27188 24948 27198
rect 23884 26292 23940 26302
rect 23884 26198 23940 26236
rect 24108 26290 24164 26302
rect 24108 26238 24110 26290
rect 24162 26238 24164 26290
rect 23772 25284 23828 25294
rect 23772 25190 23828 25228
rect 23660 23874 23716 23884
rect 24108 23716 24164 26238
rect 24220 26290 24276 26302
rect 24220 26238 24222 26290
rect 24274 26238 24276 26290
rect 24220 25732 24276 26238
rect 24332 25732 24388 25742
rect 24220 25730 24388 25732
rect 24220 25678 24334 25730
rect 24386 25678 24388 25730
rect 24220 25676 24388 25678
rect 24332 25666 24388 25676
rect 24892 25618 24948 27132
rect 26460 27188 26516 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 40236 36372 40292 36382
rect 40236 36278 40292 36316
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 26460 27094 26516 27132
rect 40012 27186 40068 27198
rect 40012 27134 40014 27186
rect 40066 27134 40068 27186
rect 28252 27074 28308 27086
rect 28252 27022 28254 27074
rect 28306 27022 28308 27074
rect 26908 26962 26964 26974
rect 26908 26910 26910 26962
rect 26962 26910 26964 26962
rect 25788 26852 25844 26862
rect 24892 25566 24894 25618
rect 24946 25566 24948 25618
rect 24892 25554 24948 25566
rect 25340 26292 25396 26302
rect 25788 26292 25844 26796
rect 26908 26852 26964 26910
rect 26908 26786 26964 26796
rect 27580 26852 27636 26862
rect 25340 26290 25844 26292
rect 25340 26238 25342 26290
rect 25394 26238 25790 26290
rect 25842 26238 25844 26290
rect 25340 26236 25844 26238
rect 24668 25506 24724 25518
rect 24668 25454 24670 25506
rect 24722 25454 24724 25506
rect 24668 25284 24724 25454
rect 24668 25218 24724 25228
rect 23772 23660 24164 23716
rect 25340 24052 25396 26236
rect 25788 26226 25844 26236
rect 26124 26292 26180 26302
rect 26124 25506 26180 26236
rect 26460 26180 26516 26190
rect 26460 26178 26740 26180
rect 26460 26126 26462 26178
rect 26514 26126 26740 26178
rect 26460 26124 26740 26126
rect 26460 26114 26516 26124
rect 26684 25618 26740 26124
rect 26684 25566 26686 25618
rect 26738 25566 26740 25618
rect 26684 25554 26740 25566
rect 27580 25618 27636 26796
rect 28252 26852 28308 27022
rect 37660 27074 37716 27086
rect 37660 27022 37662 27074
rect 37714 27022 37716 27074
rect 28476 26964 28532 26974
rect 28476 26870 28532 26908
rect 28252 26786 28308 26796
rect 28588 26852 28644 26862
rect 28588 26178 28644 26796
rect 37660 26852 37716 27022
rect 37660 26786 37716 26796
rect 37884 26964 37940 26974
rect 37884 26290 37940 26908
rect 37884 26238 37886 26290
rect 37938 26238 37940 26290
rect 37884 26226 37940 26238
rect 39900 26852 39956 26862
rect 28588 26126 28590 26178
rect 28642 26126 28644 26178
rect 28588 26114 28644 26126
rect 39900 26178 39956 26796
rect 40012 26292 40068 27134
rect 40012 26226 40068 26236
rect 39900 26126 39902 26178
rect 39954 26126 39956 26178
rect 39900 26114 39956 26126
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 27580 25566 27582 25618
rect 27634 25566 27636 25618
rect 27580 25554 27636 25566
rect 26124 25454 26126 25506
rect 26178 25454 26180 25506
rect 26124 25442 26180 25454
rect 26796 25396 26852 25406
rect 26796 25302 26852 25340
rect 26572 25284 26628 25294
rect 26572 25190 26628 25228
rect 27468 25284 27524 25294
rect 27468 25190 27524 25228
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 25340 24050 25732 24052
rect 25340 23998 25342 24050
rect 25394 23998 25732 24050
rect 25340 23996 25732 23998
rect 23548 23380 23604 23390
rect 23548 21812 23604 23324
rect 23548 21746 23604 21756
rect 23548 21588 23604 21598
rect 23436 21476 23492 21486
rect 23436 20914 23492 21420
rect 23436 20862 23438 20914
rect 23490 20862 23492 20914
rect 23436 20850 23492 20862
rect 23324 20738 23380 20748
rect 22764 20524 22932 20580
rect 22204 19182 22206 19234
rect 22258 19182 22260 19234
rect 22204 19170 22260 19182
rect 22428 19234 22484 19246
rect 22428 19182 22430 19234
rect 22482 19182 22484 19234
rect 22316 19010 22372 19022
rect 22316 18958 22318 19010
rect 22370 18958 22372 19010
rect 22316 18676 22372 18958
rect 22092 18620 22372 18676
rect 22092 18562 22148 18620
rect 22092 18510 22094 18562
rect 22146 18510 22148 18562
rect 22092 18498 22148 18510
rect 22316 17780 22372 17790
rect 22428 17780 22484 19182
rect 22316 17778 22484 17780
rect 22316 17726 22318 17778
rect 22370 17726 22484 17778
rect 22316 17724 22484 17726
rect 22764 19234 22820 20524
rect 23548 20244 23604 21532
rect 23212 20132 23268 20142
rect 23212 20038 23268 20076
rect 22764 19182 22766 19234
rect 22818 19182 22820 19234
rect 22316 17714 22372 17724
rect 21756 17502 21758 17554
rect 21810 17502 21812 17554
rect 21756 17490 21812 17502
rect 21980 17668 22036 17678
rect 21532 17444 21588 17454
rect 21532 17350 21588 17388
rect 21980 16996 22036 17612
rect 22764 17666 22820 19182
rect 22876 20018 22932 20030
rect 22876 19966 22878 20018
rect 22930 19966 22932 20018
rect 22876 18676 22932 19966
rect 22876 18610 22932 18620
rect 22764 17614 22766 17666
rect 22818 17614 22820 17666
rect 22764 17602 22820 17614
rect 22988 18228 23044 18238
rect 22988 17666 23044 18172
rect 22988 17614 22990 17666
rect 23042 17614 23044 17666
rect 22988 17602 23044 17614
rect 23436 17666 23492 17678
rect 23436 17614 23438 17666
rect 23490 17614 23492 17666
rect 22092 17556 22148 17566
rect 22092 17462 22148 17500
rect 23324 17556 23380 17566
rect 21980 16930 22036 16940
rect 23100 17442 23156 17454
rect 23100 17390 23102 17442
rect 23154 17390 23156 17442
rect 21420 16818 21476 16828
rect 22204 16884 22260 16894
rect 22204 16100 22260 16828
rect 23100 16772 23156 17390
rect 22876 16716 23156 16772
rect 22876 16210 22932 16716
rect 23324 16548 23380 17500
rect 23436 16660 23492 17614
rect 23548 16882 23604 20188
rect 23772 19124 23828 23660
rect 24108 23492 24164 23502
rect 24108 23266 24164 23436
rect 25340 23380 25396 23996
rect 25676 23938 25732 23996
rect 25676 23886 25678 23938
rect 25730 23886 25732 23938
rect 25676 23874 25732 23886
rect 28588 24050 28644 24062
rect 28588 23998 28590 24050
rect 28642 23998 28644 24050
rect 26460 23828 26516 23838
rect 26460 23826 26852 23828
rect 26460 23774 26462 23826
rect 26514 23774 26852 23826
rect 26460 23772 26852 23774
rect 26460 23762 26516 23772
rect 25340 23314 25396 23324
rect 26012 23380 26068 23390
rect 26068 23324 26404 23380
rect 26012 23286 26068 23324
rect 24108 23214 24110 23266
rect 24162 23214 24164 23266
rect 24108 23202 24164 23214
rect 24220 23268 24276 23278
rect 24220 23174 24276 23212
rect 25564 23268 25620 23278
rect 24444 23154 24500 23166
rect 24444 23102 24446 23154
rect 24498 23102 24500 23154
rect 23884 22260 23940 22270
rect 23884 20130 23940 22204
rect 24444 21810 24500 23102
rect 24444 21758 24446 21810
rect 24498 21758 24500 21810
rect 24444 21746 24500 21758
rect 23996 21588 24052 21598
rect 23996 21494 24052 21532
rect 24220 21586 24276 21598
rect 24220 21534 24222 21586
rect 24274 21534 24276 21586
rect 24108 21476 24164 21486
rect 24108 21382 24164 21420
rect 24220 20916 24276 21534
rect 25452 20916 25508 20926
rect 24220 20860 24500 20916
rect 23884 20078 23886 20130
rect 23938 20078 23940 20130
rect 23884 20066 23940 20078
rect 23996 20692 24052 20702
rect 23996 20132 24052 20636
rect 24220 20692 24276 20702
rect 24108 20132 24164 20142
rect 23996 20130 24164 20132
rect 23996 20078 24110 20130
rect 24162 20078 24164 20130
rect 23996 20076 24164 20078
rect 24108 20066 24164 20076
rect 24220 20130 24276 20636
rect 24220 20078 24222 20130
rect 24274 20078 24276 20130
rect 24220 20066 24276 20078
rect 24444 20132 24500 20860
rect 24556 20132 24612 20142
rect 24444 20076 24556 20132
rect 24332 20020 24388 20030
rect 24332 19926 24388 19964
rect 24556 20018 24612 20076
rect 25452 20020 25508 20860
rect 25564 20914 25620 23212
rect 26348 23154 26404 23324
rect 26348 23102 26350 23154
rect 26402 23102 26404 23154
rect 26348 22484 26404 23102
rect 26348 22482 26628 22484
rect 26348 22430 26350 22482
rect 26402 22430 26628 22482
rect 26348 22428 26628 22430
rect 26348 22418 26404 22428
rect 26460 21812 26516 21822
rect 26012 21588 26068 21598
rect 26012 21494 26068 21532
rect 26236 21588 26292 21598
rect 26236 21586 26404 21588
rect 26236 21534 26238 21586
rect 26290 21534 26404 21586
rect 26236 21532 26404 21534
rect 26236 21522 26292 21532
rect 26124 21476 26180 21486
rect 26124 21382 26180 21420
rect 25564 20862 25566 20914
rect 25618 20862 25620 20914
rect 25564 20850 25620 20862
rect 26236 20914 26292 20926
rect 26236 20862 26238 20914
rect 26290 20862 26292 20914
rect 25900 20692 25956 20702
rect 25900 20598 25956 20636
rect 24556 19966 24558 20018
rect 24610 19966 24612 20018
rect 24556 19954 24612 19966
rect 25116 20018 25508 20020
rect 25116 19966 25454 20018
rect 25506 19966 25508 20018
rect 25116 19964 25508 19966
rect 25116 19348 25172 19964
rect 24668 19346 25172 19348
rect 24668 19294 25118 19346
rect 25170 19294 25172 19346
rect 24668 19292 25172 19294
rect 23884 19124 23940 19134
rect 23772 19068 23884 19124
rect 23884 19058 23940 19068
rect 24668 18674 24724 19292
rect 24668 18622 24670 18674
rect 24722 18622 24724 18674
rect 24668 18610 24724 18622
rect 24220 18338 24276 18350
rect 24220 18286 24222 18338
rect 24274 18286 24276 18338
rect 24220 17556 24276 18286
rect 25004 17778 25060 19292
rect 25116 19282 25172 19292
rect 25004 17726 25006 17778
rect 25058 17726 25060 17778
rect 25004 17714 25060 17726
rect 25340 18450 25396 19964
rect 25452 19954 25508 19964
rect 26124 20578 26180 20590
rect 26124 20526 26126 20578
rect 26178 20526 26180 20578
rect 25452 19234 25508 19246
rect 25452 19182 25454 19234
rect 25506 19182 25508 19234
rect 25452 19124 25508 19182
rect 25452 19058 25508 19068
rect 25900 19124 25956 19134
rect 25900 19030 25956 19068
rect 26124 19124 26180 20526
rect 26236 20130 26292 20862
rect 26236 20078 26238 20130
rect 26290 20078 26292 20130
rect 26236 20066 26292 20078
rect 26348 20132 26404 21532
rect 26460 21474 26516 21756
rect 26460 21422 26462 21474
rect 26514 21422 26516 21474
rect 26460 20804 26516 21422
rect 26572 20916 26628 22428
rect 26796 22372 26852 23772
rect 27132 23042 27188 23054
rect 27132 22990 27134 23042
rect 27186 22990 27188 23042
rect 27132 22594 27188 22990
rect 27132 22542 27134 22594
rect 27186 22542 27188 22594
rect 27132 22530 27188 22542
rect 28140 23044 28196 23054
rect 27468 22484 27524 22494
rect 27916 22484 27972 22494
rect 27468 22482 27972 22484
rect 27468 22430 27470 22482
rect 27522 22430 27918 22482
rect 27970 22430 27972 22482
rect 27468 22428 27972 22430
rect 27468 22418 27524 22428
rect 27916 22418 27972 22428
rect 26796 22316 27188 22372
rect 27132 21810 27188 22316
rect 28140 22370 28196 22988
rect 28140 22318 28142 22370
rect 28194 22318 28196 22370
rect 28140 22306 28196 22318
rect 28588 22372 28644 23998
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 37884 23938 37940 23950
rect 37884 23886 37886 23938
rect 37938 23886 37940 23938
rect 37660 23156 37716 23166
rect 37660 23062 37716 23100
rect 29260 23044 29316 23054
rect 29260 22950 29316 22988
rect 37884 23044 37940 23886
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 37884 22978 37940 22988
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 27804 22258 27860 22270
rect 27804 22206 27806 22258
rect 27858 22206 27860 22258
rect 27132 21758 27134 21810
rect 27186 21758 27188 21810
rect 27132 21746 27188 21758
rect 27244 22148 27300 22158
rect 27244 21810 27300 22092
rect 27244 21758 27246 21810
rect 27298 21758 27300 21810
rect 27244 21746 27300 21758
rect 27804 21812 27860 22206
rect 27804 21746 27860 21756
rect 26684 21588 26740 21598
rect 26684 21494 26740 21532
rect 28588 21588 28644 22316
rect 37660 22372 37716 22382
rect 37660 22278 37716 22316
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 28588 21522 28644 21532
rect 37884 21586 37940 21598
rect 37884 21534 37886 21586
rect 37938 21534 37940 21586
rect 27020 21476 27076 21486
rect 27020 21382 27076 21420
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 26684 20916 26740 20926
rect 26628 20914 26740 20916
rect 26628 20862 26686 20914
rect 26738 20862 26740 20914
rect 26628 20860 26740 20862
rect 26572 20822 26628 20860
rect 26684 20850 26740 20860
rect 26460 20738 26516 20748
rect 37660 20802 37716 20814
rect 37660 20750 37662 20802
rect 37714 20750 37716 20802
rect 26348 19236 26404 20076
rect 29036 20132 29092 20142
rect 29036 20038 29092 20076
rect 37660 20132 37716 20750
rect 37660 20066 37716 20076
rect 28364 20020 28420 20030
rect 28364 19906 28420 19964
rect 28812 20020 28868 20030
rect 28812 19926 28868 19964
rect 37884 20020 37940 21534
rect 39900 21474 39956 21486
rect 39900 21422 39902 21474
rect 39954 21422 39956 21474
rect 39900 20916 39956 21422
rect 39900 20850 39956 20860
rect 40012 20914 40068 20926
rect 40012 20862 40014 20914
rect 40066 20862 40068 20914
rect 40012 20244 40068 20862
rect 40012 20178 40068 20188
rect 37884 19954 37940 19964
rect 28364 19854 28366 19906
rect 28418 19854 28420 19906
rect 28364 19842 28420 19854
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 40012 19346 40068 19358
rect 40012 19294 40014 19346
rect 40066 19294 40068 19346
rect 26572 19236 26628 19246
rect 26348 19180 26516 19236
rect 26124 19122 26292 19124
rect 26124 19070 26126 19122
rect 26178 19070 26292 19122
rect 26124 19068 26292 19070
rect 26124 19058 26180 19068
rect 25788 19010 25844 19022
rect 25788 18958 25790 19010
rect 25842 18958 25844 19010
rect 25788 18676 25844 18958
rect 25788 18620 26180 18676
rect 26124 18562 26180 18620
rect 26124 18510 26126 18562
rect 26178 18510 26180 18562
rect 26124 18498 26180 18510
rect 26236 18564 26292 19068
rect 26460 19122 26516 19180
rect 26460 19070 26462 19122
rect 26514 19070 26516 19122
rect 26460 19058 26516 19070
rect 26572 19122 26628 19180
rect 28252 19236 28308 19246
rect 26572 19070 26574 19122
rect 26626 19070 26628 19122
rect 26572 19058 26628 19070
rect 26684 19124 26740 19134
rect 26684 19012 26740 19068
rect 26796 19012 26852 19022
rect 26684 19010 26852 19012
rect 26684 18958 26798 19010
rect 26850 18958 26852 19010
rect 26684 18956 26852 18958
rect 26796 18946 26852 18956
rect 26236 18498 26292 18508
rect 26684 18564 26740 18574
rect 25340 18398 25342 18450
rect 25394 18398 25396 18450
rect 24220 17490 24276 17500
rect 25340 17106 25396 18398
rect 25340 17054 25342 17106
rect 25394 17054 25396 17106
rect 23884 16996 23940 17006
rect 23884 16902 23940 16940
rect 24108 16996 24164 17006
rect 24108 16994 25060 16996
rect 24108 16942 24110 16994
rect 24162 16942 25060 16994
rect 24108 16940 25060 16942
rect 24108 16930 24164 16940
rect 23548 16830 23550 16882
rect 23602 16830 23604 16882
rect 23548 16818 23604 16830
rect 23772 16660 23828 16670
rect 23436 16658 23828 16660
rect 23436 16606 23774 16658
rect 23826 16606 23828 16658
rect 23436 16604 23828 16606
rect 23772 16594 23828 16604
rect 23324 16492 23604 16548
rect 22876 16158 22878 16210
rect 22930 16158 22932 16210
rect 22876 16146 22932 16158
rect 21084 15374 21086 15426
rect 21138 15374 21140 15426
rect 21084 15362 21140 15374
rect 22092 15428 22148 15438
rect 20300 15262 20302 15314
rect 20354 15262 20356 15314
rect 20300 15250 20356 15262
rect 20524 15316 20580 15326
rect 20748 15316 20804 15326
rect 20524 15314 20804 15316
rect 20524 15262 20526 15314
rect 20578 15262 20750 15314
rect 20802 15262 20804 15314
rect 20524 15260 20804 15262
rect 20524 15250 20580 15260
rect 20748 15250 20804 15260
rect 20412 15202 20468 15214
rect 20412 15150 20414 15202
rect 20466 15150 20468 15202
rect 20412 15148 20468 15150
rect 19292 14578 19348 14588
rect 20076 15092 20468 15148
rect 17388 14530 17668 14532
rect 17388 14478 17390 14530
rect 17442 14478 17668 14530
rect 17388 14476 17668 14478
rect 17388 14466 17444 14476
rect 17612 13970 17668 14476
rect 20076 14308 20132 15092
rect 20300 14644 20356 14654
rect 20300 14550 20356 14588
rect 21308 14644 21364 14654
rect 20076 14252 20244 14308
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20188 13972 20244 14252
rect 17612 13918 17614 13970
rect 17666 13918 17668 13970
rect 17612 13906 17668 13918
rect 19964 13916 20244 13972
rect 19964 13858 20020 13916
rect 19964 13806 19966 13858
rect 20018 13806 20020 13858
rect 19964 13794 20020 13806
rect 19292 13748 19348 13758
rect 19292 13654 19348 13692
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 17052 8372 17668 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 17612 3554 17668 8372
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20188 5236 20244 5246
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 18620 3668 18676 3678
rect 17612 3502 17614 3554
rect 17666 3502 17668 3554
rect 17612 3490 17668 3502
rect 18172 3666 18676 3668
rect 18172 3614 18622 3666
rect 18674 3614 18676 3666
rect 18172 3612 18676 3614
rect 7644 3332 7700 3342
rect 7420 3330 7700 3332
rect 7420 3278 7646 3330
rect 7698 3278 7700 3330
rect 7420 3276 7700 3278
rect 7420 800 7476 3276
rect 7644 3266 7700 3276
rect 18172 800 18228 3612
rect 18620 3602 18676 3612
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 800 20244 5180
rect 21308 5122 21364 14588
rect 22092 13634 22148 15372
rect 22204 13748 22260 16044
rect 22204 13682 22260 13692
rect 22540 13748 22596 13758
rect 22540 13654 22596 13692
rect 22092 13582 22094 13634
rect 22146 13582 22148 13634
rect 22092 8428 22148 13582
rect 21308 5070 21310 5122
rect 21362 5070 21364 5122
rect 21308 5058 21364 5070
rect 21868 8372 22148 8428
rect 21868 4338 21924 8372
rect 22316 5236 22372 5246
rect 22316 5142 22372 5180
rect 21868 4286 21870 4338
rect 21922 4286 21924 4338
rect 21868 4274 21924 4286
rect 21532 4116 21588 4126
rect 21532 800 21588 4060
rect 22764 4116 22820 4126
rect 22764 4022 22820 4060
rect 23548 3554 23604 16492
rect 25004 16210 25060 16940
rect 25004 16158 25006 16210
rect 25058 16158 25060 16210
rect 25004 8428 25060 16158
rect 25340 16100 25396 17054
rect 26460 17108 26516 17118
rect 26012 16996 26068 17006
rect 25788 16884 25844 16894
rect 25788 16790 25844 16828
rect 26012 16882 26068 16940
rect 26012 16830 26014 16882
rect 26066 16830 26068 16882
rect 26012 16818 26068 16830
rect 26348 16660 26404 16670
rect 26348 16566 26404 16604
rect 25452 16100 25508 16110
rect 25396 16098 25508 16100
rect 25396 16046 25454 16098
rect 25506 16046 25508 16098
rect 25396 16044 25508 16046
rect 25340 15538 25396 16044
rect 25452 16034 25508 16044
rect 26236 15988 26292 15998
rect 25340 15486 25342 15538
rect 25394 15486 25396 15538
rect 25340 15474 25396 15486
rect 26012 15986 26292 15988
rect 26012 15934 26238 15986
rect 26290 15934 26292 15986
rect 26012 15932 26292 15934
rect 26012 15538 26068 15932
rect 26236 15922 26292 15932
rect 26012 15486 26014 15538
rect 26066 15486 26068 15538
rect 26012 15474 26068 15486
rect 26348 15428 26404 15438
rect 26460 15428 26516 17052
rect 26684 16994 26740 18508
rect 28252 18338 28308 19180
rect 37660 19236 37716 19246
rect 37660 19142 37716 19180
rect 40012 18900 40068 19294
rect 40012 18834 40068 18844
rect 28252 18286 28254 18338
rect 28306 18286 28308 18338
rect 28252 18274 28308 18286
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 27244 17108 27300 17118
rect 27244 17014 27300 17052
rect 26684 16942 26686 16994
rect 26738 16942 26740 16994
rect 26684 16930 26740 16942
rect 27580 16884 27636 16894
rect 26908 16660 26964 16670
rect 26908 16566 26964 16604
rect 26348 15426 26516 15428
rect 26348 15374 26350 15426
rect 26402 15374 26516 15426
rect 26348 15372 26516 15374
rect 27580 16212 27636 16828
rect 37884 16882 37940 16894
rect 37884 16830 37886 16882
rect 37938 16830 37940 16882
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 26348 15362 26404 15372
rect 27580 15314 27636 16156
rect 28364 16212 28420 16222
rect 28364 16118 28420 16156
rect 37660 16100 37716 16110
rect 37660 16006 37716 16044
rect 27804 15428 27860 15438
rect 27804 15334 27860 15372
rect 37884 15428 37940 16830
rect 39900 16770 39956 16782
rect 39900 16718 39902 16770
rect 39954 16718 39956 16770
rect 39900 16212 39956 16718
rect 39900 16146 39956 16156
rect 40012 16210 40068 16222
rect 40012 16158 40014 16210
rect 40066 16158 40068 16210
rect 40012 15540 40068 16158
rect 40012 15474 40068 15484
rect 37884 15362 37940 15372
rect 27580 15262 27582 15314
rect 27634 15262 27636 15314
rect 27580 15250 27636 15262
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 24556 8372 25060 8428
rect 23548 3502 23550 3554
rect 23602 3502 23604 3554
rect 23548 3490 23604 3502
rect 24220 3668 24276 3678
rect 22204 3442 22260 3454
rect 22204 3390 22206 3442
rect 22258 3390 22260 3442
rect 22204 800 22260 3390
rect 24220 800 24276 3612
rect 24556 3554 24612 8372
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 7392 0 7504 800
rect 18144 0 18256 800
rect 20160 0 20272 800
rect 21504 0 21616 800
rect 22176 0 22288 800
rect 24192 0 24304 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 17500 37436 17556 37492
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 18732 37490 18788 37492
rect 18732 37438 18734 37490
rect 18734 37438 18786 37490
rect 18786 37438 18788 37490
rect 18732 37436 18788 37438
rect 22876 38220 22932 38276
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 20860 37436 20916 37492
rect 22092 37490 22148 37492
rect 22092 37438 22094 37490
rect 22094 37438 22146 37490
rect 22146 37438 22148 37490
rect 22092 37436 22148 37438
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 15932 28028 15988 28084
rect 4172 27580 4228 27636
rect 1932 25564 1988 25620
rect 2044 24892 2100 24948
rect 4060 24556 4116 24612
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4284 25506 4340 25508
rect 4284 25454 4286 25506
rect 4286 25454 4338 25506
rect 4338 25454 4340 25506
rect 4284 25452 4340 25454
rect 13468 25452 13524 25508
rect 14700 26178 14756 26180
rect 14700 26126 14702 26178
rect 14702 26126 14754 26178
rect 14754 26126 14756 26178
rect 14700 26124 14756 26126
rect 16380 26124 16436 26180
rect 14028 25452 14084 25508
rect 15148 25452 15204 25508
rect 12908 24892 12964 24948
rect 13916 25340 13972 25396
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 14476 25228 14532 25284
rect 14588 25004 14644 25060
rect 14924 24610 14980 24612
rect 14924 24558 14926 24610
rect 14926 24558 14978 24610
rect 14978 24558 14980 24610
rect 14924 24556 14980 24558
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 17612 28028 17668 28084
rect 16604 26012 16660 26068
rect 16380 25506 16436 25508
rect 16380 25454 16382 25506
rect 16382 25454 16434 25506
rect 16434 25454 16436 25506
rect 16380 25452 16436 25454
rect 15596 25394 15652 25396
rect 15596 25342 15598 25394
rect 15598 25342 15650 25394
rect 15650 25342 15652 25394
rect 15596 25340 15652 25342
rect 15484 25004 15540 25060
rect 15596 24946 15652 24948
rect 15596 24894 15598 24946
rect 15598 24894 15650 24946
rect 15650 24894 15652 24946
rect 15596 24892 15652 24894
rect 17388 27804 17444 27860
rect 17052 26908 17108 26964
rect 19964 27858 20020 27860
rect 19964 27806 19966 27858
rect 19966 27806 20018 27858
rect 20018 27806 20020 27858
rect 19964 27804 20020 27806
rect 18172 27020 18228 27076
rect 17948 26402 18004 26404
rect 17948 26350 17950 26402
rect 17950 26350 18002 26402
rect 18002 26350 18004 26402
rect 17948 26348 18004 26350
rect 17612 26178 17668 26180
rect 17612 26126 17614 26178
rect 17614 26126 17666 26178
rect 17666 26126 17668 26178
rect 17612 26124 17668 26126
rect 18844 27074 18900 27076
rect 18844 27022 18846 27074
rect 18846 27022 18898 27074
rect 18898 27022 18900 27074
rect 18844 27020 18900 27022
rect 19292 27074 19348 27076
rect 19292 27022 19294 27074
rect 19294 27022 19346 27074
rect 19346 27022 19348 27074
rect 19292 27020 19348 27022
rect 19964 27020 20020 27076
rect 18396 26908 18452 26964
rect 18284 26348 18340 26404
rect 17500 25004 17556 25060
rect 15260 24722 15316 24724
rect 15260 24670 15262 24722
rect 15262 24670 15314 24722
rect 15314 24670 15316 24722
rect 15260 24668 15316 24670
rect 12348 23436 12404 23492
rect 13020 23042 13076 23044
rect 13020 22990 13022 23042
rect 13022 22990 13074 23042
rect 13074 22990 13076 23042
rect 13020 22988 13076 22990
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4172 22092 4228 22148
rect 14588 23548 14644 23604
rect 14140 22988 14196 23044
rect 13916 21644 13972 21700
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 10780 19404 10836 19460
rect 10108 19292 10164 19348
rect 11788 21474 11844 21476
rect 11788 21422 11790 21474
rect 11790 21422 11842 21474
rect 11842 21422 11844 21474
rect 11788 21420 11844 21422
rect 14028 20748 14084 20804
rect 14252 21756 14308 21812
rect 14476 21698 14532 21700
rect 14476 21646 14478 21698
rect 14478 21646 14530 21698
rect 14530 21646 14532 21698
rect 14476 21644 14532 21646
rect 14364 21474 14420 21476
rect 14364 21422 14366 21474
rect 14366 21422 14418 21474
rect 14418 21422 14420 21474
rect 14364 21420 14420 21422
rect 13692 20300 13748 20356
rect 13132 19906 13188 19908
rect 13132 19854 13134 19906
rect 13134 19854 13186 19906
rect 13186 19854 13188 19906
rect 13132 19852 13188 19854
rect 11004 19292 11060 19348
rect 14028 20300 14084 20356
rect 13804 19906 13860 19908
rect 13804 19854 13806 19906
rect 13806 19854 13858 19906
rect 13858 19854 13860 19906
rect 13804 19852 13860 19854
rect 13356 19404 13412 19460
rect 14140 19740 14196 19796
rect 13356 18732 13412 18788
rect 13580 19346 13636 19348
rect 13580 19294 13582 19346
rect 13582 19294 13634 19346
rect 13634 19294 13636 19346
rect 13580 19292 13636 19294
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 14140 19234 14196 19236
rect 14140 19182 14142 19234
rect 14142 19182 14194 19234
rect 14194 19182 14196 19234
rect 14140 19180 14196 19182
rect 15708 23548 15764 23604
rect 15148 23436 15204 23492
rect 15148 22428 15204 22484
rect 14700 21980 14756 22036
rect 17836 23436 17892 23492
rect 18172 23772 18228 23828
rect 15932 23324 15988 23380
rect 17388 23378 17444 23380
rect 17388 23326 17390 23378
rect 17390 23326 17442 23378
rect 17442 23326 17444 23378
rect 17388 23324 17444 23326
rect 15484 23212 15540 23268
rect 15260 21980 15316 22036
rect 15148 21868 15204 21924
rect 15036 21810 15092 21812
rect 15036 21758 15038 21810
rect 15038 21758 15090 21810
rect 15090 21758 15092 21810
rect 15036 21756 15092 21758
rect 14812 21586 14868 21588
rect 14812 21534 14814 21586
rect 14814 21534 14866 21586
rect 14866 21534 14868 21586
rect 14812 21532 14868 21534
rect 14364 19794 14420 19796
rect 14364 19742 14366 19794
rect 14366 19742 14418 19794
rect 14418 19742 14420 19794
rect 14364 19740 14420 19742
rect 15372 22204 15428 22260
rect 17948 23266 18004 23268
rect 17948 23214 17950 23266
rect 17950 23214 18002 23266
rect 18002 23214 18004 23266
rect 17948 23212 18004 23214
rect 17836 23154 17892 23156
rect 17836 23102 17838 23154
rect 17838 23102 17890 23154
rect 17890 23102 17892 23154
rect 17836 23100 17892 23102
rect 16044 22428 16100 22484
rect 15932 21868 15988 21924
rect 15596 20524 15652 20580
rect 15372 19794 15428 19796
rect 15372 19742 15374 19794
rect 15374 19742 15426 19794
rect 15426 19742 15428 19794
rect 15372 19740 15428 19742
rect 15148 19292 15204 19348
rect 14476 18450 14532 18452
rect 14476 18398 14478 18450
rect 14478 18398 14530 18450
rect 14530 18398 14532 18450
rect 14476 18396 14532 18398
rect 15372 19234 15428 19236
rect 15372 19182 15374 19234
rect 15374 19182 15426 19234
rect 15426 19182 15428 19234
rect 15372 19180 15428 19182
rect 15148 18508 15204 18564
rect 15036 18060 15092 18116
rect 16380 22258 16436 22260
rect 16380 22206 16382 22258
rect 16382 22206 16434 22258
rect 16434 22206 16436 22258
rect 16380 22204 16436 22206
rect 17052 22146 17108 22148
rect 17052 22094 17054 22146
rect 17054 22094 17106 22146
rect 17106 22094 17108 22146
rect 17052 22092 17108 22094
rect 16940 21980 16996 22036
rect 17388 21868 17444 21924
rect 18060 22428 18116 22484
rect 17500 22204 17556 22260
rect 16604 21586 16660 21588
rect 16604 21534 16606 21586
rect 16606 21534 16658 21586
rect 16658 21534 16660 21586
rect 16604 21532 16660 21534
rect 16604 20300 16660 20356
rect 16604 19964 16660 20020
rect 16492 19234 16548 19236
rect 16492 19182 16494 19234
rect 16494 19182 16546 19234
rect 16546 19182 16548 19234
rect 16492 19180 16548 19182
rect 15820 18732 15876 18788
rect 15932 18284 15988 18340
rect 15596 17388 15652 17444
rect 4284 16882 4340 16884
rect 4284 16830 4286 16882
rect 4286 16830 4338 16882
rect 4338 16830 4340 16882
rect 4284 16828 4340 16830
rect 12124 16828 12180 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 1932 16156 1988 16212
rect 14812 16882 14868 16884
rect 14812 16830 14814 16882
rect 14814 16830 14866 16882
rect 14866 16830 14868 16882
rect 14812 16828 14868 16830
rect 16828 19404 16884 19460
rect 17612 21980 17668 22036
rect 17836 20524 17892 20580
rect 17948 19964 18004 20020
rect 17276 19180 17332 19236
rect 17724 19740 17780 19796
rect 17276 19010 17332 19012
rect 17276 18958 17278 19010
rect 17278 18958 17330 19010
rect 17330 18958 17332 19010
rect 17276 18956 17332 18958
rect 17388 18844 17444 18900
rect 16716 18732 16772 18788
rect 17052 18508 17108 18564
rect 17836 19458 17892 19460
rect 17836 19406 17838 19458
rect 17838 19406 17890 19458
rect 17890 19406 17892 19458
rect 17836 19404 17892 19406
rect 21980 27804 22036 27860
rect 21756 27074 21812 27076
rect 21756 27022 21758 27074
rect 21758 27022 21810 27074
rect 21810 27022 21812 27074
rect 21756 27020 21812 27022
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20412 26236 20468 26292
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19852 24722 19908 24724
rect 19852 24670 19854 24722
rect 19854 24670 19906 24722
rect 19906 24670 19908 24722
rect 19852 24668 19908 24670
rect 20412 24668 20468 24724
rect 20300 23660 20356 23716
rect 19068 23548 19124 23604
rect 18844 23436 18900 23492
rect 18508 23154 18564 23156
rect 18508 23102 18510 23154
rect 18510 23102 18562 23154
rect 18562 23102 18564 23154
rect 18508 23100 18564 23102
rect 18396 21756 18452 21812
rect 18508 22092 18564 22148
rect 18284 21420 18340 21476
rect 18396 21532 18452 21588
rect 18284 20076 18340 20132
rect 18172 19458 18228 19460
rect 18172 19406 18174 19458
rect 18174 19406 18226 19458
rect 18226 19406 18228 19458
rect 18172 19404 18228 19406
rect 18060 18844 18116 18900
rect 18844 23100 18900 23156
rect 18844 22428 18900 22484
rect 19628 23548 19684 23604
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19964 23324 20020 23380
rect 19516 23266 19572 23268
rect 19516 23214 19518 23266
rect 19518 23214 19570 23266
rect 19570 23214 19572 23266
rect 19516 23212 19572 23214
rect 18956 21644 19012 21700
rect 18732 20076 18788 20132
rect 19180 21420 19236 21476
rect 19180 20636 19236 20692
rect 19292 20130 19348 20132
rect 19292 20078 19294 20130
rect 19294 20078 19346 20130
rect 19346 20078 19348 20130
rect 19292 20076 19348 20078
rect 19068 20018 19124 20020
rect 19068 19966 19070 20018
rect 19070 19966 19122 20018
rect 19122 19966 19124 20018
rect 19068 19964 19124 19966
rect 19404 19516 19460 19572
rect 18844 19180 18900 19236
rect 19292 18844 19348 18900
rect 18844 18732 18900 18788
rect 16492 18396 16548 18452
rect 17164 18396 17220 18452
rect 16716 18226 16772 18228
rect 16716 18174 16718 18226
rect 16718 18174 16770 18226
rect 16770 18174 16772 18226
rect 16716 18172 16772 18174
rect 16268 17612 16324 17668
rect 16604 17442 16660 17444
rect 16604 17390 16606 17442
rect 16606 17390 16658 17442
rect 16658 17390 16660 17442
rect 16604 17388 16660 17390
rect 17388 18172 17444 18228
rect 17948 18508 18004 18564
rect 15372 16098 15428 16100
rect 15372 16046 15374 16098
rect 15374 16046 15426 16098
rect 15426 16046 15428 16098
rect 15372 16044 15428 16046
rect 14252 15820 14308 15876
rect 15260 15874 15316 15876
rect 15260 15822 15262 15874
rect 15262 15822 15314 15874
rect 15314 15822 15316 15874
rect 15260 15820 15316 15822
rect 14364 15484 14420 15540
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 15036 15484 15092 15540
rect 15484 15538 15540 15540
rect 15484 15486 15486 15538
rect 15486 15486 15538 15538
rect 15538 15486 15540 15538
rect 15484 15484 15540 15486
rect 19180 18620 19236 18676
rect 18396 18508 18452 18564
rect 18284 18284 18340 18340
rect 18172 17666 18228 17668
rect 18172 17614 18174 17666
rect 18174 17614 18226 17666
rect 18226 17614 18228 17666
rect 18172 17612 18228 17614
rect 20300 23324 20356 23380
rect 19852 22204 19908 22260
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20076 21644 20132 21700
rect 23436 27858 23492 27860
rect 23436 27806 23438 27858
rect 23438 27806 23490 27858
rect 23490 27806 23492 27858
rect 23436 27804 23492 27806
rect 22428 27692 22484 27748
rect 22876 27746 22932 27748
rect 22876 27694 22878 27746
rect 22878 27694 22930 27746
rect 22930 27694 22932 27746
rect 22876 27692 22932 27694
rect 23436 26796 23492 26852
rect 23436 25340 23492 25396
rect 21868 25228 21924 25284
rect 22316 23938 22372 23940
rect 22316 23886 22318 23938
rect 22318 23886 22370 23938
rect 22370 23886 22372 23938
rect 22316 23884 22372 23886
rect 23100 23884 23156 23940
rect 21980 23826 22036 23828
rect 21980 23774 21982 23826
rect 21982 23774 22034 23826
rect 22034 23774 22036 23826
rect 21980 23772 22036 23774
rect 22092 23714 22148 23716
rect 22092 23662 22094 23714
rect 22094 23662 22146 23714
rect 22146 23662 22148 23714
rect 22092 23660 22148 23662
rect 21532 23436 21588 23492
rect 22652 23212 22708 23268
rect 21532 23100 21588 23156
rect 20524 22258 20580 22260
rect 20524 22206 20526 22258
rect 20526 22206 20578 22258
rect 20578 22206 20580 22258
rect 20524 22204 20580 22206
rect 22988 22092 23044 22148
rect 21868 21698 21924 21700
rect 21868 21646 21870 21698
rect 21870 21646 21922 21698
rect 21922 21646 21924 21698
rect 21868 21644 21924 21646
rect 22092 21756 22148 21812
rect 22764 21756 22820 21812
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19852 19516 19908 19572
rect 20524 20018 20580 20020
rect 20524 19966 20526 20018
rect 20526 19966 20578 20018
rect 20578 19966 20580 20018
rect 20524 19964 20580 19966
rect 20412 19404 20468 19460
rect 20076 19234 20132 19236
rect 20076 19182 20078 19234
rect 20078 19182 20130 19234
rect 20130 19182 20132 19234
rect 20076 19180 20132 19182
rect 20300 18956 20356 19012
rect 19628 18732 19684 18788
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20524 19516 20580 19572
rect 20860 20524 20916 20580
rect 21868 20690 21924 20692
rect 21868 20638 21870 20690
rect 21870 20638 21922 20690
rect 21922 20638 21924 20690
rect 21868 20636 21924 20638
rect 21308 20524 21364 20580
rect 20972 20188 21028 20244
rect 20636 19180 20692 19236
rect 20860 19122 20916 19124
rect 20860 19070 20862 19122
rect 20862 19070 20914 19122
rect 20914 19070 20916 19122
rect 20860 19068 20916 19070
rect 17276 15484 17332 15540
rect 14924 15148 14980 15204
rect 16268 15202 16324 15204
rect 16268 15150 16270 15202
rect 16270 15150 16322 15202
rect 16322 15150 16324 15202
rect 16268 15148 16324 15150
rect 16604 15202 16660 15204
rect 16604 15150 16606 15202
rect 16606 15150 16658 15202
rect 16658 15150 16660 15202
rect 16604 15148 16660 15150
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 18172 15314 18228 15316
rect 18172 15262 18174 15314
rect 18174 15262 18226 15314
rect 18226 15262 18228 15314
rect 18172 15260 18228 15262
rect 18284 15202 18340 15204
rect 18284 15150 18286 15202
rect 18286 15150 18338 15202
rect 18338 15150 18340 15202
rect 18284 15148 18340 15150
rect 18732 16044 18788 16100
rect 18620 15538 18676 15540
rect 18620 15486 18622 15538
rect 18622 15486 18674 15538
rect 18674 15486 18676 15538
rect 18620 15484 18676 15486
rect 19180 17442 19236 17444
rect 19180 17390 19182 17442
rect 19182 17390 19234 17442
rect 19234 17390 19236 17442
rect 19180 17388 19236 17390
rect 20412 18226 20468 18228
rect 20412 18174 20414 18226
rect 20414 18174 20466 18226
rect 20466 18174 20468 18226
rect 20412 18172 20468 18174
rect 21420 19180 21476 19236
rect 21756 19180 21812 19236
rect 19964 17612 20020 17668
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19628 16044 19684 16100
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19404 15484 19460 15540
rect 19068 15372 19124 15428
rect 19964 15426 20020 15428
rect 19964 15374 19966 15426
rect 19966 15374 20018 15426
rect 20018 15374 20020 15426
rect 19964 15372 20020 15374
rect 21084 17388 21140 17444
rect 20972 15426 21028 15428
rect 20972 15374 20974 15426
rect 20974 15374 21026 15426
rect 21026 15374 21028 15426
rect 20972 15372 21028 15374
rect 22428 20802 22484 20804
rect 22428 20750 22430 20802
rect 22430 20750 22482 20802
rect 22482 20750 22484 20802
rect 22428 20748 22484 20750
rect 24332 27916 24388 27972
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 26236 37436 26292 37492
rect 27468 37490 27524 37492
rect 27468 37438 27470 37490
rect 27470 37438 27522 37490
rect 27522 37438 27524 37490
rect 27468 37436 27524 37438
rect 25228 27970 25284 27972
rect 25228 27918 25230 27970
rect 25230 27918 25282 27970
rect 25282 27918 25284 27970
rect 25228 27916 25284 27918
rect 24556 27692 24612 27748
rect 24668 27804 24724 27860
rect 25452 27858 25508 27860
rect 25452 27806 25454 27858
rect 25454 27806 25506 27858
rect 25506 27806 25508 27858
rect 25452 27804 25508 27806
rect 24892 27132 24948 27188
rect 23884 26290 23940 26292
rect 23884 26238 23886 26290
rect 23886 26238 23938 26290
rect 23938 26238 23940 26290
rect 23884 26236 23940 26238
rect 23772 25282 23828 25284
rect 23772 25230 23774 25282
rect 23774 25230 23826 25282
rect 23826 25230 23828 25282
rect 23772 25228 23828 25230
rect 23660 23884 23716 23940
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 40236 36370 40292 36372
rect 40236 36318 40238 36370
rect 40238 36318 40290 36370
rect 40290 36318 40292 36370
rect 40236 36316 40292 36318
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 26460 27186 26516 27188
rect 26460 27134 26462 27186
rect 26462 27134 26514 27186
rect 26514 27134 26516 27186
rect 26460 27132 26516 27134
rect 25788 26796 25844 26852
rect 26908 26796 26964 26852
rect 27580 26796 27636 26852
rect 24668 25228 24724 25284
rect 26124 26236 26180 26292
rect 28476 26962 28532 26964
rect 28476 26910 28478 26962
rect 28478 26910 28530 26962
rect 28530 26910 28532 26962
rect 28476 26908 28532 26910
rect 28252 26796 28308 26852
rect 28588 26796 28644 26852
rect 37660 26796 37716 26852
rect 37884 26908 37940 26964
rect 39900 26796 39956 26852
rect 40012 26236 40068 26292
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 26796 25394 26852 25396
rect 26796 25342 26798 25394
rect 26798 25342 26850 25394
rect 26850 25342 26852 25394
rect 26796 25340 26852 25342
rect 26572 25282 26628 25284
rect 26572 25230 26574 25282
rect 26574 25230 26626 25282
rect 26626 25230 26628 25282
rect 26572 25228 26628 25230
rect 27468 25282 27524 25284
rect 27468 25230 27470 25282
rect 27470 25230 27522 25282
rect 27522 25230 27524 25282
rect 27468 25228 27524 25230
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 23548 23378 23604 23380
rect 23548 23326 23550 23378
rect 23550 23326 23602 23378
rect 23602 23326 23604 23378
rect 23548 23324 23604 23326
rect 23548 21756 23604 21812
rect 23548 21532 23604 21588
rect 23436 21420 23492 21476
rect 23324 20748 23380 20804
rect 23548 20188 23604 20244
rect 23212 20130 23268 20132
rect 23212 20078 23214 20130
rect 23214 20078 23266 20130
rect 23266 20078 23268 20130
rect 23212 20076 23268 20078
rect 21980 17666 22036 17668
rect 21980 17614 21982 17666
rect 21982 17614 22034 17666
rect 22034 17614 22036 17666
rect 21980 17612 22036 17614
rect 21532 17442 21588 17444
rect 21532 17390 21534 17442
rect 21534 17390 21586 17442
rect 21586 17390 21588 17442
rect 21532 17388 21588 17390
rect 22876 18620 22932 18676
rect 22988 18172 23044 18228
rect 22092 17554 22148 17556
rect 22092 17502 22094 17554
rect 22094 17502 22146 17554
rect 22146 17502 22148 17554
rect 22092 17500 22148 17502
rect 23324 17500 23380 17556
rect 21980 16940 22036 16996
rect 21420 16828 21476 16884
rect 22204 16828 22260 16884
rect 24108 23436 24164 23492
rect 25340 23324 25396 23380
rect 26012 23378 26068 23380
rect 26012 23326 26014 23378
rect 26014 23326 26066 23378
rect 26066 23326 26068 23378
rect 26012 23324 26068 23326
rect 24220 23266 24276 23268
rect 24220 23214 24222 23266
rect 24222 23214 24274 23266
rect 24274 23214 24276 23266
rect 24220 23212 24276 23214
rect 25564 23212 25620 23268
rect 23884 22204 23940 22260
rect 23996 21586 24052 21588
rect 23996 21534 23998 21586
rect 23998 21534 24050 21586
rect 24050 21534 24052 21586
rect 23996 21532 24052 21534
rect 24108 21474 24164 21476
rect 24108 21422 24110 21474
rect 24110 21422 24162 21474
rect 24162 21422 24164 21474
rect 24108 21420 24164 21422
rect 23996 20636 24052 20692
rect 24220 20636 24276 20692
rect 25452 20860 25508 20916
rect 24556 20076 24612 20132
rect 24332 20018 24388 20020
rect 24332 19966 24334 20018
rect 24334 19966 24386 20018
rect 24386 19966 24388 20018
rect 24332 19964 24388 19966
rect 26460 21756 26516 21812
rect 26012 21586 26068 21588
rect 26012 21534 26014 21586
rect 26014 21534 26066 21586
rect 26066 21534 26068 21586
rect 26012 21532 26068 21534
rect 26124 21474 26180 21476
rect 26124 21422 26126 21474
rect 26126 21422 26178 21474
rect 26178 21422 26180 21474
rect 26124 21420 26180 21422
rect 25900 20690 25956 20692
rect 25900 20638 25902 20690
rect 25902 20638 25954 20690
rect 25954 20638 25956 20690
rect 25900 20636 25956 20638
rect 23884 19068 23940 19124
rect 25452 19068 25508 19124
rect 25900 19122 25956 19124
rect 25900 19070 25902 19122
rect 25902 19070 25954 19122
rect 25954 19070 25956 19122
rect 25900 19068 25956 19070
rect 28140 22988 28196 23044
rect 37660 23154 37716 23156
rect 37660 23102 37662 23154
rect 37662 23102 37714 23154
rect 37714 23102 37716 23154
rect 37660 23100 37716 23102
rect 29260 23042 29316 23044
rect 29260 22990 29262 23042
rect 29262 22990 29314 23042
rect 29314 22990 29316 23042
rect 29260 22988 29316 22990
rect 40012 23548 40068 23604
rect 37884 22988 37940 23044
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 28588 22316 28644 22372
rect 27244 22146 27300 22148
rect 27244 22094 27246 22146
rect 27246 22094 27298 22146
rect 27298 22094 27300 22146
rect 27244 22092 27300 22094
rect 27804 21756 27860 21812
rect 26684 21586 26740 21588
rect 26684 21534 26686 21586
rect 26686 21534 26738 21586
rect 26738 21534 26740 21586
rect 26684 21532 26740 21534
rect 37660 22370 37716 22372
rect 37660 22318 37662 22370
rect 37662 22318 37714 22370
rect 37714 22318 37716 22370
rect 37660 22316 37716 22318
rect 40012 22204 40068 22260
rect 28588 21532 28644 21588
rect 27020 21474 27076 21476
rect 27020 21422 27022 21474
rect 27022 21422 27074 21474
rect 27074 21422 27076 21474
rect 27020 21420 27076 21422
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 26572 20860 26628 20916
rect 26460 20748 26516 20804
rect 26348 20076 26404 20132
rect 29036 20130 29092 20132
rect 29036 20078 29038 20130
rect 29038 20078 29090 20130
rect 29090 20078 29092 20130
rect 29036 20076 29092 20078
rect 37660 20076 37716 20132
rect 28364 19964 28420 20020
rect 28812 20018 28868 20020
rect 28812 19966 28814 20018
rect 28814 19966 28866 20018
rect 28866 19966 28868 20018
rect 28812 19964 28868 19966
rect 39900 20860 39956 20916
rect 40012 20188 40068 20244
rect 37884 19964 37940 20020
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 26572 19180 26628 19236
rect 28252 19180 28308 19236
rect 26684 19068 26740 19124
rect 26236 18508 26292 18564
rect 26684 18508 26740 18564
rect 24220 17500 24276 17556
rect 23884 16994 23940 16996
rect 23884 16942 23886 16994
rect 23886 16942 23938 16994
rect 23938 16942 23940 16994
rect 23884 16940 23940 16942
rect 22204 16098 22260 16100
rect 22204 16046 22206 16098
rect 22206 16046 22258 16098
rect 22258 16046 22260 16098
rect 22204 16044 22260 16046
rect 22092 15372 22148 15428
rect 19292 14588 19348 14644
rect 20300 14642 20356 14644
rect 20300 14590 20302 14642
rect 20302 14590 20354 14642
rect 20354 14590 20356 14642
rect 20300 14588 20356 14590
rect 21308 14588 21364 14644
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19292 13746 19348 13748
rect 19292 13694 19294 13746
rect 19294 13694 19346 13746
rect 19346 13694 19348 13746
rect 19292 13692 19348 13694
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 20188 5180 20244 5236
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 22204 13692 22260 13748
rect 22540 13746 22596 13748
rect 22540 13694 22542 13746
rect 22542 13694 22594 13746
rect 22594 13694 22596 13746
rect 22540 13692 22596 13694
rect 22316 5234 22372 5236
rect 22316 5182 22318 5234
rect 22318 5182 22370 5234
rect 22370 5182 22372 5234
rect 22316 5180 22372 5182
rect 21532 4060 21588 4116
rect 22764 4114 22820 4116
rect 22764 4062 22766 4114
rect 22766 4062 22818 4114
rect 22818 4062 22820 4114
rect 22764 4060 22820 4062
rect 26460 17052 26516 17108
rect 26012 16940 26068 16996
rect 25788 16882 25844 16884
rect 25788 16830 25790 16882
rect 25790 16830 25842 16882
rect 25842 16830 25844 16882
rect 25788 16828 25844 16830
rect 26348 16658 26404 16660
rect 26348 16606 26350 16658
rect 26350 16606 26402 16658
rect 26402 16606 26404 16658
rect 26348 16604 26404 16606
rect 25340 16044 25396 16100
rect 37660 19234 37716 19236
rect 37660 19182 37662 19234
rect 37662 19182 37714 19234
rect 37714 19182 37716 19234
rect 37660 19180 37716 19182
rect 40012 18844 40068 18900
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 27244 17106 27300 17108
rect 27244 17054 27246 17106
rect 27246 17054 27298 17106
rect 27298 17054 27300 17106
rect 27244 17052 27300 17054
rect 27580 16828 27636 16884
rect 26908 16658 26964 16660
rect 26908 16606 26910 16658
rect 26910 16606 26962 16658
rect 26962 16606 26964 16658
rect 26908 16604 26964 16606
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 27580 16156 27636 16212
rect 28364 16210 28420 16212
rect 28364 16158 28366 16210
rect 28366 16158 28418 16210
rect 28418 16158 28420 16210
rect 28364 16156 28420 16158
rect 37660 16098 37716 16100
rect 37660 16046 37662 16098
rect 37662 16046 37714 16098
rect 37714 16046 37716 16098
rect 37660 16044 37716 16046
rect 27804 15426 27860 15428
rect 27804 15374 27806 15426
rect 27806 15374 27858 15426
rect 27858 15374 27860 15426
rect 27804 15372 27860 15374
rect 39900 16156 39956 16212
rect 40012 15484 40068 15540
rect 37884 15372 37940 15428
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 24220 3612 24276 3668
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 22866 38220 22876 38276
rect 22932 38220 25564 38276
rect 25620 38220 25630 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 17490 37436 17500 37492
rect 17556 37436 18732 37492
rect 18788 37436 18798 37492
rect 20850 37436 20860 37492
rect 20916 37436 22092 37492
rect 22148 37436 22158 37492
rect 26226 37436 26236 37492
rect 26292 37436 27468 37492
rect 27524 37436 27534 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 41200 36372 42000 36400
rect 40226 36316 40236 36372
rect 40292 36316 42000 36372
rect 41200 36288 42000 36316
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 15922 28028 15932 28084
rect 15988 28028 17612 28084
rect 17668 28028 17678 28084
rect 17388 27860 17444 28028
rect 24322 27916 24332 27972
rect 24388 27916 25228 27972
rect 25284 27916 25294 27972
rect 17378 27804 17388 27860
rect 17444 27804 17454 27860
rect 19954 27804 19964 27860
rect 20020 27804 21980 27860
rect 22036 27804 23436 27860
rect 23492 27804 23502 27860
rect 24658 27804 24668 27860
rect 24724 27804 25452 27860
rect 25508 27804 25518 27860
rect 22418 27692 22428 27748
rect 22484 27692 22876 27748
rect 22932 27692 24556 27748
rect 24612 27692 24622 27748
rect 0 27636 800 27664
rect 0 27580 4172 27636
rect 4228 27580 4238 27636
rect 0 27552 800 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 24882 27132 24892 27188
rect 24948 27132 26460 27188
rect 26516 27132 26526 27188
rect 18162 27020 18172 27076
rect 18228 27020 18844 27076
rect 18900 27020 19292 27076
rect 19348 27020 19964 27076
rect 20020 27020 20030 27076
rect 20132 27020 21756 27076
rect 21812 27020 21822 27076
rect 20132 26964 20188 27020
rect 41200 26964 42000 26992
rect 17042 26908 17052 26964
rect 17108 26908 18396 26964
rect 18452 26908 20188 26964
rect 28466 26908 28476 26964
rect 28532 26908 37884 26964
rect 37940 26908 37950 26964
rect 39900 26908 42000 26964
rect 39900 26852 39956 26908
rect 41200 26880 42000 26908
rect 23426 26796 23436 26852
rect 23492 26796 25788 26852
rect 25844 26796 26908 26852
rect 26964 26796 26974 26852
rect 27570 26796 27580 26852
rect 27636 26796 28252 26852
rect 28308 26796 28588 26852
rect 28644 26796 37660 26852
rect 37716 26796 37726 26852
rect 39890 26796 39900 26852
rect 39956 26796 39966 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 17938 26348 17948 26404
rect 18004 26348 18284 26404
rect 18340 26348 18350 26404
rect 41200 26292 42000 26320
rect 20402 26236 20412 26292
rect 20468 26236 23884 26292
rect 23940 26236 26124 26292
rect 26180 26236 26190 26292
rect 40002 26236 40012 26292
rect 40068 26236 42000 26292
rect 41200 26208 42000 26236
rect 14690 26124 14700 26180
rect 14756 26124 15148 26180
rect 16370 26124 16380 26180
rect 16436 26124 17612 26180
rect 17668 26124 17678 26180
rect 15092 26068 15148 26124
rect 15092 26012 16604 26068
rect 16660 26012 16670 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 0 25620 800 25648
rect 0 25564 1932 25620
rect 1988 25564 1998 25620
rect 0 25536 800 25564
rect 4274 25452 4284 25508
rect 4340 25452 13468 25508
rect 13524 25452 13534 25508
rect 14018 25452 14028 25508
rect 14084 25452 15148 25508
rect 15204 25452 16380 25508
rect 16436 25452 16446 25508
rect 13468 25284 13524 25452
rect 13906 25340 13916 25396
rect 13972 25340 15596 25396
rect 15652 25340 15662 25396
rect 23426 25340 23436 25396
rect 23492 25340 26796 25396
rect 26852 25340 26862 25396
rect 13468 25228 14476 25284
rect 14532 25228 14542 25284
rect 21858 25228 21868 25284
rect 21924 25228 23772 25284
rect 23828 25228 24668 25284
rect 24724 25228 24734 25284
rect 26562 25228 26572 25284
rect 26628 25228 27468 25284
rect 27524 25228 27534 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 14578 25004 14588 25060
rect 14644 25004 15484 25060
rect 15540 25004 17500 25060
rect 17556 25004 17566 25060
rect 0 24948 800 24976
rect 0 24892 2044 24948
rect 2100 24892 2110 24948
rect 12898 24892 12908 24948
rect 12964 24892 15596 24948
rect 15652 24892 15662 24948
rect 0 24864 800 24892
rect 15092 24668 15260 24724
rect 15316 24668 15326 24724
rect 19842 24668 19852 24724
rect 19908 24668 20412 24724
rect 20468 24668 20478 24724
rect 15092 24612 15148 24668
rect 4050 24556 4060 24612
rect 4116 24556 14924 24612
rect 14980 24556 15148 24612
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 22306 23884 22316 23940
rect 22372 23884 23100 23940
rect 23156 23884 23660 23940
rect 23716 23884 23726 23940
rect 18162 23772 18172 23828
rect 18228 23772 21980 23828
rect 22036 23772 22046 23828
rect 20290 23660 20300 23716
rect 20356 23660 22092 23716
rect 22148 23660 22158 23716
rect 41200 23604 42000 23632
rect 14578 23548 14588 23604
rect 14644 23548 15708 23604
rect 15764 23548 19068 23604
rect 19124 23548 19628 23604
rect 19684 23548 19694 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 41200 23520 42000 23548
rect 12338 23436 12348 23492
rect 12404 23436 15148 23492
rect 15204 23436 15214 23492
rect 17826 23436 17836 23492
rect 17892 23436 18844 23492
rect 18900 23436 18910 23492
rect 21522 23436 21532 23492
rect 21588 23436 24108 23492
rect 24164 23436 24174 23492
rect 15922 23324 15932 23380
rect 15988 23324 17388 23380
rect 17444 23324 19964 23380
rect 20020 23324 20030 23380
rect 20290 23324 20300 23380
rect 20356 23324 23548 23380
rect 23604 23324 25340 23380
rect 25396 23324 26012 23380
rect 26068 23324 26078 23380
rect 19964 23268 20020 23324
rect 15474 23212 15484 23268
rect 15540 23212 17948 23268
rect 18004 23212 19516 23268
rect 19572 23212 19582 23268
rect 19964 23212 22652 23268
rect 22708 23212 22718 23268
rect 24210 23212 24220 23268
rect 24276 23212 25564 23268
rect 25620 23212 31948 23268
rect 31892 23156 31948 23212
rect 17826 23100 17836 23156
rect 17892 23100 18508 23156
rect 18564 23100 18574 23156
rect 18834 23100 18844 23156
rect 18900 23100 21532 23156
rect 21588 23100 21598 23156
rect 31892 23100 37660 23156
rect 37716 23100 37726 23156
rect 13010 22988 13020 23044
rect 13076 22988 14140 23044
rect 14196 22988 14206 23044
rect 28130 22988 28140 23044
rect 28196 22988 29260 23044
rect 29316 22988 37884 23044
rect 37940 22988 37950 23044
rect 41200 22932 42000 22960
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 41200 22848 42000 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 15138 22428 15148 22484
rect 15204 22428 16044 22484
rect 16100 22428 16110 22484
rect 18050 22428 18060 22484
rect 18116 22428 18844 22484
rect 18900 22428 18910 22484
rect 28578 22316 28588 22372
rect 28644 22316 37660 22372
rect 37716 22316 37726 22372
rect 41200 22260 42000 22288
rect 15362 22204 15372 22260
rect 15428 22204 16380 22260
rect 16436 22204 17500 22260
rect 17556 22204 17566 22260
rect 19842 22204 19852 22260
rect 19908 22204 20524 22260
rect 20580 22204 23884 22260
rect 23940 22204 23950 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 41200 22176 42000 22204
rect 4162 22092 4172 22148
rect 4228 22092 17052 22148
rect 17108 22092 18508 22148
rect 18564 22092 18574 22148
rect 22978 22092 22988 22148
rect 23044 22092 27244 22148
rect 27300 22092 27310 22148
rect 14690 21980 14700 22036
rect 14756 21980 15260 22036
rect 15316 21980 15326 22036
rect 16930 21980 16940 22036
rect 16996 21980 17612 22036
rect 17668 21980 17678 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 15138 21868 15148 21924
rect 15204 21868 15932 21924
rect 15988 21868 17388 21924
rect 17444 21868 17454 21924
rect 14242 21756 14252 21812
rect 14308 21756 15036 21812
rect 15092 21756 15102 21812
rect 18386 21756 18396 21812
rect 18452 21756 22092 21812
rect 22148 21756 22158 21812
rect 22754 21756 22764 21812
rect 22820 21756 23548 21812
rect 23604 21756 23614 21812
rect 26450 21756 26460 21812
rect 26516 21756 27804 21812
rect 27860 21756 27870 21812
rect 13906 21644 13916 21700
rect 13972 21644 13982 21700
rect 14466 21644 14476 21700
rect 14532 21644 18956 21700
rect 19012 21644 19022 21700
rect 20066 21644 20076 21700
rect 20132 21644 21868 21700
rect 21924 21644 21934 21700
rect 13916 21588 13972 21644
rect 13916 21532 14812 21588
rect 14868 21532 14878 21588
rect 16594 21532 16604 21588
rect 16660 21532 18396 21588
rect 18452 21532 18462 21588
rect 23538 21532 23548 21588
rect 23604 21532 23996 21588
rect 24052 21532 26012 21588
rect 26068 21532 26078 21588
rect 26674 21532 26684 21588
rect 26740 21532 28588 21588
rect 28644 21532 28654 21588
rect 11778 21420 11788 21476
rect 11844 21420 14364 21476
rect 14420 21420 14430 21476
rect 18274 21420 18284 21476
rect 18340 21420 19180 21476
rect 19236 21420 19246 21476
rect 23426 21420 23436 21476
rect 23492 21420 24108 21476
rect 24164 21420 24174 21476
rect 26114 21420 26124 21476
rect 26180 21420 27020 21476
rect 27076 21420 27086 21476
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 41200 20916 42000 20944
rect 25442 20860 25452 20916
rect 25508 20860 26572 20916
rect 26628 20860 26638 20916
rect 39890 20860 39900 20916
rect 39956 20860 42000 20916
rect 41200 20832 42000 20860
rect 14018 20748 14028 20804
rect 14084 20748 14094 20804
rect 22418 20748 22428 20804
rect 22484 20748 23324 20804
rect 23380 20748 26460 20804
rect 26516 20748 26526 20804
rect 14028 20580 14084 20748
rect 19170 20636 19180 20692
rect 19236 20636 21868 20692
rect 21924 20636 23996 20692
rect 24052 20636 24062 20692
rect 24210 20636 24220 20692
rect 24276 20636 25900 20692
rect 25956 20636 25966 20692
rect 14028 20524 15596 20580
rect 15652 20524 17836 20580
rect 17892 20524 20860 20580
rect 20916 20524 21308 20580
rect 21364 20524 21374 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 13682 20300 13692 20356
rect 13748 20300 14028 20356
rect 14084 20300 16604 20356
rect 16660 20300 16670 20356
rect 41200 20244 42000 20272
rect 20962 20188 20972 20244
rect 21028 20188 23548 20244
rect 23604 20188 23614 20244
rect 40002 20188 40012 20244
rect 40068 20188 42000 20244
rect 41200 20160 42000 20188
rect 18274 20076 18284 20132
rect 18340 20076 18732 20132
rect 18788 20076 19292 20132
rect 19348 20076 19358 20132
rect 23202 20076 23212 20132
rect 23268 20076 24556 20132
rect 24612 20076 26348 20132
rect 26404 20076 26414 20132
rect 29026 20076 29036 20132
rect 29092 20076 37660 20132
rect 37716 20076 37726 20132
rect 16594 19964 16604 20020
rect 16660 19964 17948 20020
rect 18004 19964 18014 20020
rect 19058 19964 19068 20020
rect 19124 19964 20524 20020
rect 20580 19964 20590 20020
rect 24322 19964 24332 20020
rect 24388 19964 28364 20020
rect 28420 19964 28812 20020
rect 28868 19964 37884 20020
rect 37940 19964 37950 20020
rect 13122 19852 13132 19908
rect 13188 19852 13804 19908
rect 13860 19852 13870 19908
rect 14130 19740 14140 19796
rect 14196 19740 14364 19796
rect 14420 19740 14430 19796
rect 15362 19740 15372 19796
rect 15428 19740 17724 19796
rect 17780 19740 17790 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 17836 19516 19404 19572
rect 19460 19516 19852 19572
rect 19908 19516 20524 19572
rect 20580 19516 20590 19572
rect 17836 19460 17892 19516
rect 10770 19404 10780 19460
rect 10836 19404 13356 19460
rect 13412 19404 13422 19460
rect 16818 19404 16828 19460
rect 16884 19404 17836 19460
rect 17892 19404 17902 19460
rect 18162 19404 18172 19460
rect 18228 19404 20412 19460
rect 20468 19404 20478 19460
rect 10098 19292 10108 19348
rect 10164 19292 11004 19348
rect 11060 19292 13580 19348
rect 13636 19292 15148 19348
rect 15204 19292 15214 19348
rect 14130 19180 14140 19236
rect 14196 19180 15372 19236
rect 15428 19180 15438 19236
rect 16482 19180 16492 19236
rect 16548 19180 17276 19236
rect 17332 19180 17342 19236
rect 18834 19180 18844 19236
rect 18900 19180 20076 19236
rect 20132 19180 20636 19236
rect 20692 19180 21420 19236
rect 21476 19180 21756 19236
rect 21812 19180 21822 19236
rect 26562 19180 26572 19236
rect 26628 19180 28252 19236
rect 28308 19180 37660 19236
rect 37716 19180 37726 19236
rect 20850 19068 20860 19124
rect 20916 19068 23884 19124
rect 23940 19068 25452 19124
rect 25508 19068 25518 19124
rect 25890 19068 25900 19124
rect 25956 19068 26684 19124
rect 26740 19068 26750 19124
rect 17266 18956 17276 19012
rect 17332 18956 20300 19012
rect 20356 18956 20366 19012
rect 41200 18900 42000 18928
rect 15092 18844 17388 18900
rect 17444 18844 18060 18900
rect 18116 18844 19292 18900
rect 19348 18844 19358 18900
rect 40002 18844 40012 18900
rect 40068 18844 42000 18900
rect 15092 18788 15148 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 41200 18816 42000 18844
rect 13346 18732 13356 18788
rect 13412 18732 15148 18788
rect 15810 18732 15820 18788
rect 15876 18732 16716 18788
rect 16772 18732 16782 18788
rect 18834 18732 18844 18788
rect 18900 18732 19628 18788
rect 19684 18732 19694 18788
rect 16716 18676 16772 18732
rect 16716 18620 19180 18676
rect 19236 18620 22876 18676
rect 22932 18620 22942 18676
rect 15138 18508 15148 18564
rect 15204 18508 16772 18564
rect 17042 18508 17052 18564
rect 17108 18508 17948 18564
rect 18004 18508 18014 18564
rect 18386 18508 18396 18564
rect 18452 18508 26236 18564
rect 26292 18508 26684 18564
rect 26740 18508 26750 18564
rect 16716 18452 16772 18508
rect 14466 18396 14476 18452
rect 14532 18396 16492 18452
rect 16548 18396 16558 18452
rect 16716 18396 17164 18452
rect 17220 18396 17230 18452
rect 15092 18284 15932 18340
rect 15988 18284 18284 18340
rect 18340 18284 18350 18340
rect 15026 18060 15036 18116
rect 15092 18060 15148 18284
rect 16706 18172 16716 18228
rect 16772 18172 17388 18228
rect 17444 18172 17454 18228
rect 20402 18172 20412 18228
rect 20468 18172 22988 18228
rect 23044 18172 23054 18228
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 16258 17612 16268 17668
rect 16324 17612 18172 17668
rect 18228 17612 18238 17668
rect 19954 17612 19964 17668
rect 20020 17612 21980 17668
rect 22036 17612 22046 17668
rect 22082 17500 22092 17556
rect 22148 17500 23324 17556
rect 23380 17500 24220 17556
rect 24276 17500 24286 17556
rect 15586 17388 15596 17444
rect 15652 17388 16604 17444
rect 16660 17388 16670 17444
rect 19170 17388 19180 17444
rect 19236 17388 21084 17444
rect 21140 17388 21532 17444
rect 21588 17388 21598 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 26450 17052 26460 17108
rect 26516 17052 27244 17108
rect 27300 17052 27310 17108
rect 21970 16940 21980 16996
rect 22036 16940 23884 16996
rect 23940 16940 26012 16996
rect 26068 16940 26078 16996
rect 4274 16828 4284 16884
rect 4340 16828 12124 16884
rect 12180 16828 14812 16884
rect 14868 16828 14878 16884
rect 21410 16828 21420 16884
rect 21476 16828 22204 16884
rect 22260 16828 22270 16884
rect 25778 16828 25788 16884
rect 25844 16828 27580 16884
rect 27636 16828 27646 16884
rect 26338 16604 26348 16660
rect 26404 16604 26908 16660
rect 26964 16604 26974 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 0 16212 800 16240
rect 41200 16212 42000 16240
rect 0 16156 1932 16212
rect 1988 16156 1998 16212
rect 27570 16156 27580 16212
rect 27636 16156 28364 16212
rect 28420 16156 31948 16212
rect 39890 16156 39900 16212
rect 39956 16156 42000 16212
rect 0 16128 800 16156
rect 31892 16100 31948 16156
rect 41200 16128 42000 16156
rect 15362 16044 15372 16100
rect 15428 16044 18732 16100
rect 18788 16044 19628 16100
rect 19684 16044 19694 16100
rect 22194 16044 22204 16100
rect 22260 16044 25340 16100
rect 25396 16044 25406 16100
rect 31892 16044 37660 16100
rect 37716 16044 37726 16100
rect 14242 15820 14252 15876
rect 14308 15820 15260 15876
rect 15316 15820 15326 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 41200 15540 42000 15568
rect 14354 15484 14364 15540
rect 14420 15484 15036 15540
rect 15092 15484 15484 15540
rect 15540 15484 17276 15540
rect 17332 15484 17342 15540
rect 18610 15484 18620 15540
rect 18676 15484 19404 15540
rect 19460 15484 19470 15540
rect 40002 15484 40012 15540
rect 40068 15484 42000 15540
rect 41200 15456 42000 15484
rect 19058 15372 19068 15428
rect 19124 15372 19964 15428
rect 20020 15372 20030 15428
rect 20962 15372 20972 15428
rect 21028 15372 22092 15428
rect 22148 15372 22158 15428
rect 27794 15372 27804 15428
rect 27860 15372 37884 15428
rect 37940 15372 37950 15428
rect 19068 15316 19124 15372
rect 18162 15260 18172 15316
rect 18228 15260 19124 15316
rect 14914 15148 14924 15204
rect 14980 15148 16268 15204
rect 16324 15148 16334 15204
rect 16594 15148 16604 15204
rect 16660 15148 18284 15204
rect 18340 15148 18350 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 19282 14588 19292 14644
rect 19348 14588 20300 14644
rect 20356 14588 21308 14644
rect 21364 14588 21374 14644
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 19282 13692 19292 13748
rect 19348 13692 22204 13748
rect 22260 13692 22540 13748
rect 22596 13692 22606 13748
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 20178 5180 20188 5236
rect 20244 5180 22316 5236
rect 22372 5180 22382 5236
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 21522 4060 21532 4116
rect 21588 4060 22764 4116
rect 22820 4060 22830 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 24210 3612 24220 3668
rect 24276 3612 25564 3668
rect 25620 3612 25630 3668
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _092_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16016 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _093_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18480 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _094_
timestamp 1698175906
transform 1 0 15680 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _095_
timestamp 1698175906
transform 1 0 16352 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _096_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17696 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _097_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12992 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _098_
timestamp 1698175906
transform 1 0 16352 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _099_
timestamp 1698175906
transform 1 0 17024 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _101_
timestamp 1698175906
transform 1 0 16240 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _102_
timestamp 1698175906
transform -1 0 19376 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19488 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _104_
timestamp 1698175906
transform 1 0 16128 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_
timestamp 1698175906
transform 1 0 14000 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18704 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20384 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23520 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18368 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _111_
timestamp 1698175906
transform 1 0 22512 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23520 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_
timestamp 1698175906
transform -1 0 19712 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _114_
timestamp 1698175906
transform -1 0 21280 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform 1 0 18144 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _116_
timestamp 1698175906
transform -1 0 20720 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13664 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _119_
timestamp 1698175906
transform 1 0 14112 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _120_
timestamp 1698175906
transform -1 0 16352 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _121_
timestamp 1698175906
transform -1 0 15344 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14448 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _123_
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _124_
timestamp 1698175906
transform -1 0 16240 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _125_
timestamp 1698175906
transform 1 0 14336 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _126_
timestamp 1698175906
transform 1 0 18032 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _127_
timestamp 1698175906
transform -1 0 16800 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698175906
transform 1 0 22736 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _129_
timestamp 1698175906
transform 1 0 26320 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _130_
timestamp 1698175906
transform 1 0 18368 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _131_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19152 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _132_
timestamp 1698175906
transform 1 0 15120 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18704 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _134_
timestamp 1698175906
transform 1 0 25424 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _135_
timestamp 1698175906
transform -1 0 20384 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _136_
timestamp 1698175906
transform 1 0 18928 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _137_
timestamp 1698175906
transform -1 0 19152 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18928 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _139_
timestamp 1698175906
transform 1 0 18368 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _140_
timestamp 1698175906
transform -1 0 18144 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _141_
timestamp 1698175906
transform 1 0 17136 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform 1 0 17696 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _143_
timestamp 1698175906
transform -1 0 14784 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _144_
timestamp 1698175906
transform -1 0 14224 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform -1 0 17808 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _146_
timestamp 1698175906
transform -1 0 18704 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _147_
timestamp 1698175906
transform -1 0 17136 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_
timestamp 1698175906
transform -1 0 17136 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _149_
timestamp 1698175906
transform -1 0 15344 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _150_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15008 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _151_
timestamp 1698175906
transform 1 0 23968 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _152_
timestamp 1698175906
transform 1 0 23856 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _153_
timestamp 1698175906
transform 1 0 25648 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _154_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26544 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _155_
timestamp 1698175906
transform -1 0 26544 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _156_
timestamp 1698175906
transform 1 0 19376 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _157_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23744 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _158_
timestamp 1698175906
transform 1 0 25760 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _159_
timestamp 1698175906
transform 1 0 20384 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform -1 0 21728 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _161_
timestamp 1698175906
transform 1 0 19712 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _162_
timestamp 1698175906
transform 1 0 15120 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _163_
timestamp 1698175906
transform -1 0 13104 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _164_
timestamp 1698175906
transform -1 0 27776 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _165_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _166_
timestamp 1698175906
transform -1 0 23968 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _167_
timestamp 1698175906
transform -1 0 26992 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _168_
timestamp 1698175906
transform -1 0 25088 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _169_
timestamp 1698175906
transform 1 0 23744 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _170_
timestamp 1698175906
transform -1 0 25760 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _171_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _172_
timestamp 1698175906
transform 1 0 20048 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _173_
timestamp 1698175906
transform -1 0 21840 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _174_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 26880 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _175_
timestamp 1698175906
transform 1 0 26880 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _176_
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _177_
timestamp 1698175906
transform 1 0 21840 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _178_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _179_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21392 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _180_
timestamp 1698175906
transform -1 0 22512 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _181_
timestamp 1698175906
transform 1 0 22064 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _182_
timestamp 1698175906
transform 1 0 27664 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _183_
timestamp 1698175906
transform -1 0 27664 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _184_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21952 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _185_
timestamp 1698175906
transform 1 0 19040 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _186_
timestamp 1698175906
transform 1 0 9856 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _187_
timestamp 1698175906
transform 1 0 10864 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _188_
timestamp 1698175906
transform 1 0 12096 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _189_
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _190_
timestamp 1698175906
transform 1 0 14000 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _191_
timestamp 1698175906
transform 1 0 25200 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _192_
timestamp 1698175906
transform 1 0 17248 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _193_
timestamp 1698175906
transform -1 0 19040 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_
timestamp 1698175906
transform -1 0 16576 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1698175906
transform 1 0 13776 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _196_
timestamp 1698175906
transform -1 0 15232 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _197_
timestamp 1698175906
transform 1 0 22512 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _198_
timestamp 1698175906
transform 1 0 25312 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _199_
timestamp 1698175906
transform 1 0 25312 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _200_
timestamp 1698175906
transform 1 0 17696 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1698175906
transform 1 0 11872 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_
timestamp 1698175906
transform 1 0 25536 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform 1 0 23408 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform 1 0 19824 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform 1 0 25536 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform 1 0 20048 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform 1 0 21168 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform 1 0 26208 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _211_
timestamp 1698175906
transform 1 0 27328 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _212_
timestamp 1698175906
transform 1 0 28000 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _213_
timestamp 1698175906
transform 1 0 28560 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25312 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__CLK
timestamp 1698175906
transform 1 0 22512 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__CLK
timestamp 1698175906
transform 1 0 13552 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__CLK
timestamp 1698175906
transform 1 0 14672 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__CLK
timestamp 1698175906
transform 1 0 15568 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__CLK
timestamp 1698175906
transform 1 0 17360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__CLK
timestamp 1698175906
transform -1 0 17696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__CLK
timestamp 1698175906
transform 1 0 24976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__CLK
timestamp 1698175906
transform 1 0 19264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__CLK
timestamp 1698175906
transform 1 0 16576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1698175906
transform -1 0 17696 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__CLK
timestamp 1698175906
transform 1 0 15456 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__CLK
timestamp 1698175906
transform 1 0 26656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__CLK
timestamp 1698175906
transform 1 0 25088 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__CLK
timestamp 1698175906
transform 1 0 21952 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__CLK
timestamp 1698175906
transform 1 0 15120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1698175906
transform 1 0 26880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform -1 0 23520 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 25312 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 23520 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 25984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 17024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18256 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 20384 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 21392 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_52 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7168 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_54 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7392 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_59 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7952 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698175906
transform 1 0 8848 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_174
timestamp 1698175906
transform 1 0 20832 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_178
timestamp 1698175906
transform 1 0 21280 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_180
timestamp 1698175906
transform 1 0 21504 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_203
timestamp 1698175906
transform 1 0 24080 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_235
timestamp 1698175906
transform 1 0 27664 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_243
timestamp 1698175906
transform 1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_146
timestamp 1698175906
transform 1 0 17696 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_154
timestamp 1698175906
transform 1 0 18592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_187
timestamp 1698175906
transform 1 0 22288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_191
timestamp 1698175906
transform 1 0 22736 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1698175906
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_111
timestamp 1698175906
transform 1 0 13776 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698175906
transform 1 0 20496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_88
timestamp 1698175906
transform 1 0 11200 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_92
timestamp 1698175906
transform 1 0 11648 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_94
timestamp 1698175906
transform 1 0 11872 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_124
timestamp 1698175906
transform 1 0 15232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_128
timestamp 1698175906
transform 1 0 15680 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698175906
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_146
timestamp 1698175906
transform 1 0 17696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_148
timestamp 1698175906
transform 1 0 17920 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_178
timestamp 1698175906
transform 1 0 21280 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_216
timestamp 1698175906
transform 1 0 25536 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_218
timestamp 1698175906
transform 1 0 25760 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_225
timestamp 1698175906
transform 1 0 26544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_229
timestamp 1698175906
transform 1 0 26992 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_231
timestamp 1698175906
transform 1 0 27216 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_238
timestamp 1698175906
transform 1 0 28000 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_270
timestamp 1698175906
transform 1 0 31584 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698175906
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_115
timestamp 1698175906
transform 1 0 14224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_119
timestamp 1698175906
transform 1 0 14672 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_121
timestamp 1698175906
transform 1 0 14896 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_130
timestamp 1698175906
transform 1 0 15904 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_146
timestamp 1698175906
transform 1 0 17696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_150
timestamp 1698175906
transform 1 0 18144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_152
timestamp 1698175906
transform 1 0 18368 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_159
timestamp 1698175906
transform 1 0 19152 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_181
timestamp 1698175906
transform 1 0 21616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_183
timestamp 1698175906
transform 1 0 21840 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_213
timestamp 1698175906
transform 1 0 25200 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 37296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 4480 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_104
timestamp 1698175906
transform 1 0 12992 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_112
timestamp 1698175906
transform 1 0 13888 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_116
timestamp 1698175906
transform 1 0 14336 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_118
timestamp 1698175906
transform 1 0 14560 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_125
timestamp 1698175906
transform 1 0 15344 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_133
timestamp 1698175906
transform 1 0 16240 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698175906
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_156
timestamp 1698175906
transform 1 0 18816 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_188
timestamp 1698175906
transform 1 0 22400 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_196
timestamp 1698175906
transform 1 0 23296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_205
timestamp 1698175906
transform 1 0 24304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_216
timestamp 1698175906
transform 1 0 25536 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_233
timestamp 1698175906
transform 1 0 27440 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_265
timestamp 1698175906
transform 1 0 31024 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_273
timestamp 1698175906
transform 1 0 31920 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698175906
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 36512 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 37408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_141
timestamp 1698175906
transform 1 0 17136 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_145
timestamp 1698175906
transform 1 0 17584 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_153
timestamp 1698175906
transform 1 0 18480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_157
timestamp 1698175906
transform 1 0 18928 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_170
timestamp 1698175906
transform 1 0 20384 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_189
timestamp 1698175906
transform 1 0 22512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_198
timestamp 1698175906
transform 1 0 23520 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_206
timestamp 1698175906
transform 1 0 24416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_210
timestamp 1698175906
transform 1 0 24864 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_213
timestamp 1698175906
transform 1 0 25200 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_104
timestamp 1698175906
transform 1 0 12992 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_112
timestamp 1698175906
transform 1 0 13888 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_124
timestamp 1698175906
transform 1 0 15232 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_128
timestamp 1698175906
transform 1 0 15680 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_130
timestamp 1698175906
transform 1 0 15904 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_161
timestamp 1698175906
transform 1 0 19376 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_173
timestamp 1698175906
transform 1 0 20720 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_206
timestamp 1698175906
transform 1 0 24416 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_242
timestamp 1698175906
transform 1 0 28448 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_274
timestamp 1698175906
transform 1 0 32032 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 40320 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 9072 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698175906
transform 1 0 9520 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_75
timestamp 1698175906
transform 1 0 9744 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_111
timestamp 1698175906
transform 1 0 13776 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_118
timestamp 1698175906
transform 1 0 14560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_122
timestamp 1698175906
transform 1 0 15008 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_139
timestamp 1698175906
transform 1 0 16912 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_158
timestamp 1698175906
transform 1 0 19040 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_193
timestamp 1698175906
transform 1 0 22960 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_209
timestamp 1698175906
transform 1 0 24752 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_211
timestamp 1698175906
transform 1 0 24976 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_214
timestamp 1698175906
transform 1 0 25312 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_228
timestamp 1698175906
transform 1 0 26880 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_118
timestamp 1698175906
transform 1 0 14560 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_122
timestamp 1698175906
transform 1 0 15008 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_179
timestamp 1698175906
transform 1 0 21392 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_187
timestamp 1698175906
transform 1 0 22288 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_197
timestamp 1698175906
transform 1 0 23408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_199
timestamp 1698175906
transform 1 0 23632 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_249
timestamp 1698175906
transform 1 0 29232 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_265
timestamp 1698175906
transform 1 0 31024 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_273
timestamp 1698175906
transform 1 0 31920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698175906
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 40320 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_111
timestamp 1698175906
transform 1 0 13776 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_119
timestamp 1698175906
transform 1 0 14672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_224
timestamp 1698175906
transform 1 0 26432 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_228
timestamp 1698175906
transform 1 0 26880 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_80
timestamp 1698175906
transform 1 0 10304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_84
timestamp 1698175906
transform 1 0 10752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_125
timestamp 1698175906
transform 1 0 15344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_127
timestamp 1698175906
transform 1 0 15568 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_150
timestamp 1698175906
transform 1 0 18144 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_216
timestamp 1698175906
transform 1 0 25536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_234
timestamp 1698175906
transform 1 0 27552 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_266
timestamp 1698175906
transform 1 0 31136 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_274
timestamp 1698175906
transform 1 0 32032 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_117
timestamp 1698175906
transform 1 0 14448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_121
timestamp 1698175906
transform 1 0 14896 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_129
timestamp 1698175906
transform 1 0 15792 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_131
timestamp 1698175906
transform 1 0 16016 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_136
timestamp 1698175906
transform 1 0 16576 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_241
timestamp 1698175906
transform 1 0 28336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_88
timestamp 1698175906
transform 1 0 11200 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_125
timestamp 1698175906
transform 1 0 15344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_129
timestamp 1698175906
transform 1 0 15792 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698175906
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_158
timestamp 1698175906
transform 1 0 19040 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_160
timestamp 1698175906
transform 1 0 19264 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_196
timestamp 1698175906
transform 1 0 23296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_200
timestamp 1698175906
transform 1 0 23744 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698175906
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_251
timestamp 1698175906
transform 1 0 29456 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_267
timestamp 1698175906
transform 1 0 31248 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_275
timestamp 1698175906
transform 1 0 32144 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_109
timestamp 1698175906
transform 1 0 13552 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_120
timestamp 1698175906
transform 1 0 14784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_122
timestamp 1698175906
transform 1 0 15008 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_125
timestamp 1698175906
transform 1 0 15344 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_157
timestamp 1698175906
transform 1 0 18928 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_173
timestamp 1698175906
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_181
timestamp 1698175906
transform 1 0 21616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_195
timestamp 1698175906
transform 1 0 23184 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_211
timestamp 1698175906
transform 1 0 24976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_213
timestamp 1698175906
transform 1 0 25200 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_88
timestamp 1698175906
transform 1 0 11200 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_92
timestamp 1698175906
transform 1 0 11648 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_132
timestamp 1698175906
transform 1 0 16128 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_150
timestamp 1698175906
transform 1 0 18144 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_158
timestamp 1698175906
transform 1 0 19040 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_162
timestamp 1698175906
transform 1 0 19488 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_172
timestamp 1698175906
transform 1 0 20608 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_204
timestamp 1698175906
transform 1 0 24192 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698175906
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_182
timestamp 1698175906
transform 1 0 21728 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_186
timestamp 1698175906
transform 1 0 22176 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_194
timestamp 1698175906
transform 1 0 23072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_202
timestamp 1698175906
transform 1 0 23968 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_212
timestamp 1698175906
transform 1 0 25088 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_220
timestamp 1698175906
transform 1 0 25984 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_229
timestamp 1698175906
transform 1 0 26992 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_231
timestamp 1698175906
transform 1 0 27216 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_236
timestamp 1698175906
transform 1 0 27776 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 4480 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_104
timestamp 1698175906
transform 1 0 12992 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_108
timestamp 1698175906
transform 1 0 13440 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_110
timestamp 1698175906
transform 1 0 13664 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_151
timestamp 1698175906
transform 1 0 18256 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_183
timestamp 1698175906
transform 1 0 21840 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_199
timestamp 1698175906
transform 1 0 23632 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_245
timestamp 1698175906
transform 1 0 28784 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 32368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 36512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 37408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_123
timestamp 1698175906
transform 1 0 15120 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_127
timestamp 1698175906
transform 1 0 15568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_158
timestamp 1698175906
transform 1 0 19040 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_162
timestamp 1698175906
transform 1 0 19488 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_166
timestamp 1698175906
transform 1 0 19936 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_192
timestamp 1698175906
transform 1 0 22848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_196
timestamp 1698175906
transform 1 0 23296 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_226
timestamp 1698175906
transform 1 0 26656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_230
timestamp 1698175906
transform 1 0 27104 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_147
timestamp 1698175906
transform 1 0 17808 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_163
timestamp 1698175906
transform 1 0 19600 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_194
timestamp 1698175906
transform 1 0 23072 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_198
timestamp 1698175906
transform 1 0 23520 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698175906
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_218
timestamp 1698175906
transform 1 0 25760 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_250
timestamp 1698175906
transform 1 0 29344 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_266
timestamp 1698175906
transform 1 0 31136 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_274
timestamp 1698175906
transform 1 0 32032 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_278
timestamp 1698175906
transform 1 0 32480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_183
timestamp 1698175906
transform 1 0 21840 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_215
timestamp 1698175906
transform 1 0 25424 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_231
timestamp 1698175906
transform 1 0 27216 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_239
timestamp 1698175906
transform 1 0 28112 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_243
timestamp 1698175906
transform 1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_333
timestamp 1698175906
transform 1 0 38640 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_341
timestamp 1698175906
transform 1 0 39536 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_144
timestamp 1698175906
transform 1 0 17472 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_171
timestamp 1698175906
transform 1 0 20496 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_201
timestamp 1698175906
transform 1 0 23856 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_220
timestamp 1698175906
transform 1 0 25984 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_222
timestamp 1698175906
transform 1 0 26208 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_249
timestamp 1698175906
transform 1 0 29232 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_265
timestamp 1698175906
transform 1 0 31024 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_273
timestamp 1698175906
transform 1 0 31920 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_277
timestamp 1698175906
transform 1 0 32368 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita37_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 39984 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita37_26
timestamp 1698175906
transform -1 0 7952 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37520 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform -1 0 24192 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform -1 0 24192 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 37520 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 37520 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 37520 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 26320 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 20944 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform -1 0 4480 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 4480 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 17584 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 37520 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 17472 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 21616 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 41200 16128 42000 16240 0 FreeSans 448 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 41200 36288 42000 36400 0 FreeSans 448 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 41200 26880 42000 26992 0 FreeSans 448 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 41200 15456 42000 15568 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 41200 26208 42000 26320 0 FreeSans 448 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 41200 20160 42000 20272 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 26208 41200 26320 42000 0 FreeSans 448 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 22848 41200 22960 42000 0 FreeSans 448 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 20832 41200 20944 42000 0 FreeSans 448 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 17472 41200 17584 42000 0 FreeSans 448 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 18816 41200 18928 42000 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 41200 18816 42000 18928 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 20776 28168 20776 28168 0 _000_
rlabel metal2 27160 22064 27160 22064 0 _001_
rlabel metal2 21000 22736 21000 22736 0 _002_
rlabel metal2 22120 18592 22120 18592 0 _003_
rlabel metal2 27160 22792 27160 22792 0 _004_
rlabel metal2 22904 16464 22904 16464 0 _005_
rlabel metal2 20216 14112 20216 14112 0 _006_
rlabel metal2 13384 19656 13384 19656 0 _007_
rlabel metal3 13104 21448 13104 21448 0 _008_
rlabel metal2 14168 22736 14168 22736 0 _009_
rlabel metal2 14448 17752 14448 17752 0 _010_
rlabel metal2 14952 14896 14952 14896 0 _011_
rlabel metal2 26152 18592 26152 18592 0 _012_
rlabel metal2 18200 14784 18200 14784 0 _013_
rlabel metal2 18032 26040 18032 26040 0 _014_
rlabel metal2 13944 24752 13944 24752 0 _015_
rlabel metal3 14924 26152 14924 26152 0 _016_
rlabel metal2 14280 15624 14280 15624 0 _017_
rlabel metal2 23464 21168 23464 21168 0 _018_
rlabel metal2 26040 15736 26040 15736 0 _019_
rlabel metal2 26264 20496 26264 20496 0 _020_
rlabel metal2 19824 24920 19824 24920 0 _021_
rlabel metal2 12824 25032 12824 25032 0 _022_
rlabel metal2 26712 25872 26712 25872 0 _023_
rlabel metal2 24360 27552 24360 27552 0 _024_
rlabel metal2 17696 25480 17696 25480 0 _025_
rlabel metal2 14168 23800 14168 23800 0 _026_
rlabel metal2 17136 27832 17136 27832 0 _027_
rlabel metal3 20972 27048 20972 27048 0 _028_
rlabel metal2 15624 16856 15624 16856 0 _029_
rlabel metal2 15064 16408 15064 16408 0 _030_
rlabel metal2 24472 22456 24472 22456 0 _031_
rlabel metal3 26656 16632 26656 16632 0 _032_
rlabel metal2 26488 16240 26488 16240 0 _033_
rlabel metal3 22232 22232 22232 22232 0 _034_
rlabel metal2 24248 20384 24248 20384 0 _035_
rlabel metal2 20216 26964 20216 26964 0 _036_
rlabel metal2 20552 24976 20552 24976 0 _037_
rlabel metal2 12936 25144 12936 25144 0 _038_
rlabel metal3 27048 25256 27048 25256 0 _039_
rlabel metal2 21952 26936 21952 26936 0 _040_
rlabel metal2 27832 22008 27832 22008 0 _041_
rlabel metal2 24304 25704 24304 25704 0 _042_
rlabel metal3 25088 27832 25088 27832 0 _043_
rlabel metal2 20944 27048 20944 27048 0 _044_
rlabel metal2 20776 27496 20776 27496 0 _045_
rlabel metal3 26600 21448 26600 21448 0 _046_
rlabel metal2 21448 21616 21448 21616 0 _047_
rlabel metal2 20216 23128 20216 23128 0 _048_
rlabel metal2 22400 17752 22400 17752 0 _049_
rlabel metal2 22232 20048 22232 20048 0 _050_
rlabel metal2 27720 22456 27720 22456 0 _051_
rlabel metal3 17248 17640 17248 17640 0 _052_
rlabel metal3 19040 20104 19040 20104 0 _053_
rlabel metal2 16184 20888 16184 20888 0 _054_
rlabel metal3 17360 19432 17360 19432 0 _055_
rlabel metal2 20440 19656 20440 19656 0 _056_
rlabel metal2 16912 21672 16912 21672 0 _057_
rlabel metal2 20328 18760 20328 18760 0 _058_
rlabel metal2 23016 17920 23016 17920 0 _059_
rlabel metal2 19208 18536 19208 18536 0 _060_
rlabel metal3 18760 23240 18760 23240 0 _061_
rlabel metal3 24976 16968 24976 16968 0 _062_
rlabel metal3 15904 22232 15904 22232 0 _063_
rlabel metal2 14056 21448 14056 21448 0 _064_
rlabel metal2 14616 22120 14616 22120 0 _065_
rlabel metal2 18984 21896 18984 21896 0 _066_
rlabel metal2 21000 18928 21000 18928 0 _067_
rlabel metal2 23464 17136 23464 17136 0 _068_
rlabel metal3 16688 23352 16688 23352 0 _069_
rlabel metal2 27272 21952 27272 21952 0 _070_
rlabel metal3 20384 17416 20384 17416 0 _071_
rlabel metal2 20664 15288 20664 15288 0 _072_
rlabel metal2 18648 17360 18648 17360 0 _073_
rlabel metal3 14280 19768 14280 19768 0 _074_
rlabel metal2 14280 21728 14280 21728 0 _075_
rlabel metal2 15176 21784 15176 21784 0 _076_
rlabel metal2 13832 21896 13832 21896 0 _077_
rlabel metal2 16632 18200 16632 18200 0 _078_
rlabel metal2 15064 18256 15064 18256 0 _079_
rlabel metal3 17472 15176 17472 15176 0 _080_
rlabel metal2 26320 21560 26320 21560 0 _081_
rlabel metal2 26768 18984 26768 18984 0 _082_
rlabel metal3 20944 19208 20944 19208 0 _083_
rlabel metal2 25480 19152 25480 19152 0 _084_
rlabel metal2 17752 19152 17752 19152 0 _085_
rlabel metal2 26208 19096 26208 19096 0 _086_
rlabel metal2 18760 16016 18760 16016 0 _087_
rlabel metal2 19208 15736 19208 15736 0 _088_
rlabel metal2 19208 20832 19208 20832 0 _089_
rlabel metal2 21560 24416 21560 24416 0 _090_
rlabel metal2 17584 27832 17584 27832 0 _091_
rlabel metal3 2478 27608 2478 27608 0 clk
rlabel metal2 21896 22008 21896 22008 0 clknet_0_clk
rlabel metal2 14728 22064 14728 22064 0 clknet_1_0__leaf_clk
rlabel metal2 23520 27048 23520 27048 0 clknet_1_1__leaf_clk
rlabel metal2 14000 20552 14000 20552 0 dut37.count\[0\]
rlabel metal2 13832 21448 13832 21448 0 dut37.count\[1\]
rlabel metal2 16184 22456 16184 22456 0 dut37.count\[2\]
rlabel metal3 16912 19208 16912 19208 0 dut37.count\[3\]
rlabel metal2 37912 16128 37912 16128 0 net1
rlabel metal2 28392 19936 28392 19936 0 net10
rlabel metal3 25704 27160 25704 27160 0 net11
rlabel metal3 23744 27720 23744 27720 0 net12
rlabel metal3 31920 23184 31920 23184 0 net13
rlabel metal2 21616 37240 21616 37240 0 net14
rlabel metal2 4088 25424 4088 25424 0 net15
rlabel metal2 12152 16016 12152 16016 0 net16
rlabel metal2 17192 28056 17192 28056 0 net17
rlabel metal2 13496 25536 13496 25536 0 net18
rlabel metal2 15960 27608 15960 27608 0 net19
rlabel metal2 28616 22792 28616 22792 0 net2
rlabel metal2 21336 9856 21336 9856 0 net20
rlabel metal2 28280 18760 28280 18760 0 net21
rlabel metal2 17640 5964 17640 5964 0 net22
rlabel metal2 21896 6356 21896 6356 0 net23
rlabel metal2 24584 5964 24584 5964 0 net24
rlabel metal3 40754 36344 40754 36344 0 net25
rlabel metal2 7448 2030 7448 2030 0 net26
rlabel metal3 23016 23912 23016 23912 0 net3
rlabel metal3 22736 17528 22736 17528 0 net4
rlabel metal2 28168 22680 28168 22680 0 net5
rlabel metal2 37912 26600 37912 26600 0 net6
rlabel metal2 27608 15736 27608 15736 0 net7
rlabel metal2 28280 26936 28280 26936 0 net8
rlabel metal3 33376 20104 33376 20104 0 net9
rlabel metal2 39928 16464 39928 16464 0 segm[0]
rlabel metal2 40040 22344 40040 22344 0 segm[10]
rlabel metal2 22232 39690 22232 39690 0 segm[11]
rlabel metal2 22232 2086 22232 2086 0 segm[12]
rlabel metal2 40040 23800 40040 23800 0 segm[13]
rlabel metal2 39928 26488 39928 26488 0 segm[2]
rlabel metal2 40040 15848 40040 15848 0 segm[3]
rlabel metal2 40040 26712 40040 26712 0 segm[5]
rlabel metal2 40040 20552 40040 20552 0 segm[6]
rlabel metal2 39928 21168 39928 21168 0 segm[7]
rlabel metal2 26264 39354 26264 39354 0 segm[8]
rlabel metal2 22904 39746 22904 39746 0 segm[9]
rlabel metal3 40642 22904 40642 22904 0 sel[0]
rlabel metal2 20888 39354 20888 39354 0 sel[10]
rlabel metal3 1358 25592 1358 25592 0 sel[11]
rlabel metal3 1358 16184 1358 16184 0 sel[1]
rlabel metal2 17528 39354 17528 39354 0 sel[2]
rlabel metal3 1414 24920 1414 24920 0 sel[3]
rlabel metal2 18872 39690 18872 39690 0 sel[4]
rlabel metal2 20216 2982 20216 2982 0 sel[5]
rlabel metal2 40040 19096 40040 19096 0 sel[6]
rlabel metal2 18200 2198 18200 2198 0 sel[7]
rlabel metal2 21560 2422 21560 2422 0 sel[8]
rlabel metal2 24248 2198 24248 2198 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
