magic
tech gf180mcuD
magscale 1 5
timestamp 1699643551
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9311 19137 9337 19143
rect 9311 19105 9337 19111
rect 11215 19137 11241 19143
rect 11215 19105 11241 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 8801 18999 8807 19025
rect 8833 18999 8839 19025
rect 10873 18999 10879 19025
rect 10905 18999 10911 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 11383 18745 11409 18751
rect 11383 18713 11409 18719
rect 13119 18745 13145 18751
rect 13119 18713 13145 18719
rect 10481 18607 10487 18633
rect 10513 18607 10519 18633
rect 10929 18607 10935 18633
rect 10961 18607 10967 18633
rect 12665 18607 12671 18633
rect 12697 18607 12703 18633
rect 10033 18551 10039 18577
rect 10065 18551 10071 18577
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 8695 18353 8721 18359
rect 8695 18321 8721 18327
rect 11159 18353 11185 18359
rect 11159 18321 11185 18327
rect 13063 18353 13089 18359
rect 13063 18321 13089 18327
rect 8185 18215 8191 18241
rect 8217 18215 8223 18241
rect 10649 18215 10655 18241
rect 10681 18215 10687 18241
rect 12553 18215 12559 18241
rect 12585 18215 12591 18241
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 20119 17345 20145 17351
rect 20119 17313 20145 17319
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 10655 14321 10681 14327
rect 11097 14295 11103 14321
rect 11129 14295 11135 14321
rect 10655 14289 10681 14295
rect 10817 14239 10823 14265
rect 10849 14239 10855 14265
rect 10985 14239 10991 14265
rect 11017 14239 11023 14265
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 10761 14015 10767 14041
rect 10793 14015 10799 14041
rect 7009 13903 7015 13929
rect 7041 13903 7047 13929
rect 9305 13903 9311 13929
rect 9337 13903 9343 13929
rect 8807 13873 8833 13879
rect 7345 13847 7351 13873
rect 7377 13847 7383 13873
rect 8409 13847 8415 13873
rect 8441 13847 8447 13873
rect 8807 13841 8833 13847
rect 9143 13873 9169 13879
rect 12727 13873 12753 13879
rect 9641 13847 9647 13873
rect 9673 13847 9679 13873
rect 9143 13841 9169 13847
rect 12727 13841 12753 13847
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 10207 13649 10233 13655
rect 10207 13617 10233 13623
rect 13623 13649 13649 13655
rect 13623 13617 13649 13623
rect 8415 13593 8441 13599
rect 10711 13593 10737 13599
rect 20007 13593 20033 13599
rect 8185 13567 8191 13593
rect 8217 13567 8223 13593
rect 10033 13567 10039 13593
rect 10065 13567 10071 13593
rect 12329 13567 12335 13593
rect 12361 13567 12367 13593
rect 8415 13561 8441 13567
rect 10711 13561 10737 13567
rect 20007 13561 20033 13567
rect 12503 13537 12529 13543
rect 6729 13511 6735 13537
rect 6761 13511 6767 13537
rect 8633 13511 8639 13537
rect 8665 13511 8671 13537
rect 10929 13511 10935 13537
rect 10961 13511 10967 13537
rect 12503 13505 12529 13511
rect 13119 13537 13145 13543
rect 13119 13505 13145 13511
rect 13399 13537 13425 13543
rect 13399 13505 13425 13511
rect 13567 13537 13593 13543
rect 18825 13511 18831 13537
rect 18857 13511 18863 13537
rect 13567 13505 13593 13511
rect 10263 13481 10289 13487
rect 12951 13481 12977 13487
rect 7121 13455 7127 13481
rect 7153 13455 7159 13481
rect 8969 13455 8975 13481
rect 9001 13455 9007 13481
rect 11265 13455 11271 13481
rect 11297 13455 11303 13481
rect 12665 13455 12671 13481
rect 12697 13455 12703 13481
rect 10263 13449 10289 13455
rect 12951 13449 12977 13455
rect 13063 13481 13089 13487
rect 13063 13449 13089 13455
rect 13343 13481 13369 13487
rect 13343 13449 13369 13455
rect 13623 13481 13649 13487
rect 13623 13449 13649 13455
rect 13231 13425 13257 13431
rect 13231 13393 13257 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 7687 13257 7713 13263
rect 7687 13225 7713 13231
rect 8247 13257 8273 13263
rect 8247 13225 8273 13231
rect 8751 13257 8777 13263
rect 9367 13257 9393 13263
rect 9025 13231 9031 13257
rect 9057 13231 9063 13257
rect 8751 13225 8777 13231
rect 9367 13225 9393 13231
rect 9927 13257 9953 13263
rect 9927 13225 9953 13231
rect 9983 13257 10009 13263
rect 9983 13225 10009 13231
rect 10767 13257 10793 13263
rect 10767 13225 10793 13231
rect 11271 13257 11297 13263
rect 11271 13225 11297 13231
rect 11663 13257 11689 13263
rect 11663 13225 11689 13231
rect 7799 13201 7825 13207
rect 7799 13169 7825 13175
rect 7855 13201 7881 13207
rect 7855 13169 7881 13175
rect 8639 13201 8665 13207
rect 8639 13169 8665 13175
rect 8807 13201 8833 13207
rect 8807 13169 8833 13175
rect 10879 13201 10905 13207
rect 10879 13169 10905 13175
rect 11551 13201 11577 13207
rect 11551 13169 11577 13175
rect 11775 13201 11801 13207
rect 11775 13169 11801 13175
rect 7519 13145 7545 13151
rect 7519 13113 7545 13119
rect 7575 13145 7601 13151
rect 8135 13145 8161 13151
rect 8017 13119 8023 13145
rect 8049 13119 8055 13145
rect 7575 13113 7601 13119
rect 8135 13113 8161 13119
rect 8191 13145 8217 13151
rect 10039 13145 10065 13151
rect 11215 13145 11241 13151
rect 14295 13145 14321 13151
rect 8353 13119 8359 13145
rect 8385 13119 8391 13145
rect 9137 13119 9143 13145
rect 9169 13119 9175 13145
rect 9809 13119 9815 13145
rect 9841 13119 9847 13145
rect 10145 13119 10151 13145
rect 10177 13119 10183 13145
rect 10649 13119 10655 13145
rect 10681 13119 10687 13145
rect 10985 13119 10991 13145
rect 11017 13119 11023 13145
rect 11433 13119 11439 13145
rect 11465 13119 11471 13145
rect 12665 13119 12671 13145
rect 12697 13119 12703 13145
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 8191 13113 8217 13119
rect 10039 13113 10065 13119
rect 11215 13113 11241 13119
rect 14295 13113 14321 13119
rect 9423 13089 9449 13095
rect 10761 13063 10767 13089
rect 10793 13063 10799 13089
rect 11489 13063 11495 13089
rect 11521 13063 11527 13089
rect 13001 13063 13007 13089
rect 13033 13063 13039 13089
rect 14065 13063 14071 13089
rect 14097 13063 14103 13089
rect 9423 13057 9449 13063
rect 20007 13033 20033 13039
rect 20007 13001 20033 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 14631 12809 14657 12815
rect 13225 12783 13231 12809
rect 13257 12783 13263 12809
rect 14289 12783 14295 12809
rect 14321 12783 14327 12809
rect 14631 12777 14657 12783
rect 8415 12753 8441 12759
rect 8415 12721 8441 12727
rect 8583 12753 8609 12759
rect 12889 12727 12895 12753
rect 12921 12727 12927 12753
rect 8583 12721 8609 12727
rect 8527 12697 8553 12703
rect 8527 12665 8553 12671
rect 12503 12697 12529 12703
rect 12503 12665 12529 12671
rect 12559 12697 12585 12703
rect 12559 12665 12585 12671
rect 12671 12641 12697 12647
rect 12671 12609 12697 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 7687 12473 7713 12479
rect 7687 12441 7713 12447
rect 11383 12473 11409 12479
rect 11383 12441 11409 12447
rect 11047 12417 11073 12423
rect 11047 12385 11073 12391
rect 11215 12417 11241 12423
rect 11215 12385 11241 12391
rect 11271 12417 11297 12423
rect 11271 12385 11297 12391
rect 10711 12361 10737 12367
rect 6057 12335 6063 12361
rect 6089 12335 6095 12361
rect 10711 12329 10737 12335
rect 10935 12361 10961 12367
rect 10935 12329 10961 12335
rect 7967 12305 7993 12311
rect 6393 12279 6399 12305
rect 6425 12279 6431 12305
rect 7457 12279 7463 12305
rect 7489 12279 7495 12305
rect 7967 12273 7993 12279
rect 10823 12305 10849 12311
rect 10823 12273 10849 12279
rect 8023 12249 8049 12255
rect 8023 12217 8049 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 7799 12025 7825 12031
rect 12105 11999 12111 12025
rect 12137 11999 12143 12025
rect 13617 11999 13623 12025
rect 13649 11999 13655 12025
rect 7799 11993 7825 11999
rect 7855 11969 7881 11975
rect 7855 11937 7881 11943
rect 8079 11969 8105 11975
rect 8079 11937 8105 11943
rect 8359 11969 8385 11975
rect 10375 11969 10401 11975
rect 8633 11943 8639 11969
rect 8665 11943 8671 11969
rect 8857 11943 8863 11969
rect 8889 11943 8895 11969
rect 10649 11943 10655 11969
rect 10681 11943 10687 11969
rect 13337 11943 13343 11969
rect 13369 11943 13375 11969
rect 8359 11937 8385 11943
rect 10375 11937 10401 11943
rect 7519 11913 7545 11919
rect 8185 11887 8191 11913
rect 8217 11887 8223 11913
rect 11041 11887 11047 11913
rect 11073 11887 11079 11913
rect 7519 11881 7545 11887
rect 7575 11857 7601 11863
rect 7575 11825 7601 11831
rect 7743 11857 7769 11863
rect 7743 11825 7769 11831
rect 8583 11857 8609 11863
rect 12335 11857 12361 11863
rect 10201 11831 10207 11857
rect 10233 11831 10239 11857
rect 8583 11825 8609 11831
rect 12335 11825 12361 11831
rect 13455 11857 13481 11863
rect 13455 11825 13481 11831
rect 13567 11857 13593 11863
rect 13567 11825 13593 11831
rect 13623 11857 13649 11863
rect 13623 11825 13649 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 7575 11689 7601 11695
rect 7575 11657 7601 11663
rect 7911 11689 7937 11695
rect 8303 11689 8329 11695
rect 10319 11689 10345 11695
rect 8073 11663 8079 11689
rect 8105 11663 8111 11689
rect 10089 11663 10095 11689
rect 10121 11663 10127 11689
rect 7911 11657 7937 11663
rect 8303 11657 8329 11663
rect 10319 11657 10345 11663
rect 10991 11689 11017 11695
rect 10991 11657 11017 11663
rect 10599 11633 10625 11639
rect 7401 11607 7407 11633
rect 7433 11607 7439 11633
rect 7737 11607 7743 11633
rect 7769 11607 7775 11633
rect 10705 11607 10711 11633
rect 10737 11607 10743 11633
rect 13673 11607 13679 11633
rect 13705 11607 13711 11633
rect 10599 11601 10625 11607
rect 9927 11577 9953 11583
rect 10823 11577 10849 11583
rect 14967 11577 14993 11583
rect 5497 11551 5503 11577
rect 5529 11551 5535 11577
rect 7289 11551 7295 11577
rect 7321 11551 7327 11577
rect 10425 11551 10431 11577
rect 10457 11551 10463 11577
rect 10873 11551 10879 11577
rect 10905 11551 10911 11577
rect 13281 11551 13287 11577
rect 13313 11551 13319 11577
rect 18825 11551 18831 11577
rect 18857 11551 18863 11577
rect 9927 11545 9953 11551
rect 10823 11545 10849 11551
rect 14967 11545 14993 11551
rect 5833 11495 5839 11521
rect 5865 11495 5871 11521
rect 6897 11495 6903 11521
rect 6929 11495 6935 11521
rect 14737 11495 14743 11521
rect 14769 11495 14775 11521
rect 8247 11465 8273 11471
rect 8247 11433 8273 11439
rect 8415 11465 8441 11471
rect 8415 11433 8441 11439
rect 10263 11465 10289 11471
rect 10263 11433 10289 11439
rect 20007 11465 20033 11471
rect 20007 11433 20033 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 7519 11297 7545 11303
rect 7519 11265 7545 11271
rect 11103 11297 11129 11303
rect 11103 11265 11129 11271
rect 7015 11241 7041 11247
rect 10319 11241 10345 11247
rect 14911 11241 14937 11247
rect 8409 11215 8415 11241
rect 8441 11215 8447 11241
rect 10089 11215 10095 11241
rect 10121 11215 10127 11241
rect 14289 11215 14295 11241
rect 14321 11215 14327 11241
rect 7015 11209 7041 11215
rect 10319 11209 10345 11215
rect 14911 11209 14937 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 7855 11185 7881 11191
rect 11215 11185 11241 11191
rect 7345 11159 7351 11185
rect 7377 11159 7383 11185
rect 8577 11159 8583 11185
rect 8609 11159 8615 11185
rect 9921 11159 9927 11185
rect 9953 11159 9959 11185
rect 10985 11159 10991 11185
rect 11017 11159 11023 11185
rect 7855 11153 7881 11159
rect 11215 11153 11241 11159
rect 11887 11185 11913 11191
rect 11887 11153 11913 11159
rect 12111 11185 12137 11191
rect 14743 11185 14769 11191
rect 12889 11159 12895 11185
rect 12921 11159 12927 11185
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 12111 11153 12137 11159
rect 14743 11153 14769 11159
rect 10655 11129 10681 11135
rect 11271 11129 11297 11135
rect 7681 11103 7687 11129
rect 7713 11103 7719 11129
rect 8857 11103 8863 11129
rect 8889 11103 8895 11129
rect 10817 11103 10823 11129
rect 10849 11103 10855 11129
rect 10655 11097 10681 11103
rect 11271 11097 11297 11103
rect 12391 11129 12417 11135
rect 14575 11129 14601 11135
rect 13225 11103 13231 11129
rect 13257 11103 13263 11129
rect 12391 11097 12417 11103
rect 14575 11097 14601 11103
rect 14631 11129 14657 11135
rect 14631 11097 14657 11103
rect 7463 11073 7489 11079
rect 7463 11041 7489 11047
rect 8023 11073 8049 11079
rect 9031 11073 9057 11079
rect 8185 11047 8191 11073
rect 8217 11047 8223 11073
rect 8023 11041 8049 11047
rect 9031 11041 9057 11047
rect 9311 11073 9337 11079
rect 12167 11073 12193 11079
rect 9473 11047 9479 11073
rect 9505 11047 9511 11073
rect 9311 11041 9337 11047
rect 12167 11041 12193 11047
rect 12223 11073 12249 11079
rect 12553 11047 12559 11073
rect 12585 11047 12591 11073
rect 12223 11041 12249 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 9031 10905 9057 10911
rect 9031 10873 9057 10879
rect 9535 10905 9561 10911
rect 9535 10873 9561 10879
rect 12671 10905 12697 10911
rect 12671 10873 12697 10879
rect 13287 10905 13313 10911
rect 13287 10873 13313 10879
rect 14015 10905 14041 10911
rect 14015 10873 14041 10879
rect 7463 10849 7489 10855
rect 7463 10817 7489 10823
rect 7575 10849 7601 10855
rect 7575 10817 7601 10823
rect 13119 10849 13145 10855
rect 13119 10817 13145 10823
rect 7351 10793 7377 10799
rect 7351 10761 7377 10767
rect 7687 10793 7713 10799
rect 7687 10761 7713 10767
rect 7855 10793 7881 10799
rect 12727 10793 12753 10799
rect 9697 10767 9703 10793
rect 9729 10767 9735 10793
rect 7855 10761 7881 10767
rect 12727 10761 12753 10767
rect 13231 10793 13257 10799
rect 13231 10761 13257 10767
rect 13343 10793 13369 10799
rect 13903 10793 13929 10799
rect 13449 10767 13455 10793
rect 13481 10767 13487 10793
rect 13343 10761 13369 10767
rect 13903 10761 13929 10767
rect 14071 10793 14097 10799
rect 14071 10761 14097 10767
rect 8073 10711 8079 10737
rect 8105 10711 8111 10737
rect 9249 10711 9255 10737
rect 9281 10711 9287 10737
rect 11545 10711 11551 10737
rect 11577 10711 11583 10737
rect 12671 10681 12697 10687
rect 12671 10649 12697 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 967 10457 993 10463
rect 6791 10457 6817 10463
rect 4993 10431 4999 10457
rect 5025 10431 5031 10457
rect 7849 10431 7855 10457
rect 7881 10431 7887 10457
rect 10929 10431 10935 10457
rect 10961 10431 10967 10457
rect 967 10425 993 10431
rect 6791 10425 6817 10431
rect 10991 10401 11017 10407
rect 2137 10375 2143 10401
rect 2169 10375 2175 10401
rect 6393 10375 6399 10401
rect 6425 10375 6431 10401
rect 7513 10375 7519 10401
rect 7545 10375 7551 10401
rect 10033 10375 10039 10401
rect 10065 10375 10071 10401
rect 11097 10375 11103 10401
rect 11129 10375 11135 10401
rect 11545 10375 11551 10401
rect 11577 10375 11583 10401
rect 10991 10369 11017 10375
rect 6057 10319 6063 10345
rect 6089 10319 6095 10345
rect 13057 10319 13063 10345
rect 13089 10319 13095 10345
rect 7407 10289 7433 10295
rect 7407 10257 7433 10263
rect 11439 10289 11465 10295
rect 11439 10257 11465 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 7127 10121 7153 10127
rect 9983 10121 10009 10127
rect 8745 10095 8751 10121
rect 8777 10095 8783 10121
rect 7127 10089 7153 10095
rect 9983 10089 10009 10095
rect 12279 10121 12305 10127
rect 12279 10089 12305 10095
rect 13287 10121 13313 10127
rect 13287 10089 13313 10095
rect 6903 10065 6929 10071
rect 6903 10033 6929 10039
rect 6959 10065 6985 10071
rect 6959 10033 6985 10039
rect 7799 10065 7825 10071
rect 9927 10065 9953 10071
rect 9249 10039 9255 10065
rect 9281 10039 9287 10065
rect 7799 10033 7825 10039
rect 9927 10033 9953 10039
rect 10207 10065 10233 10071
rect 10207 10033 10233 10039
rect 10319 10065 10345 10071
rect 11047 10065 11073 10071
rect 12167 10065 12193 10071
rect 10649 10039 10655 10065
rect 10681 10039 10687 10065
rect 11321 10039 11327 10065
rect 11353 10039 11359 10065
rect 11657 10039 11663 10065
rect 11689 10039 11695 10065
rect 10319 10033 10345 10039
rect 11047 10033 11073 10039
rect 12167 10033 12193 10039
rect 12335 10065 12361 10071
rect 12335 10033 12361 10039
rect 12615 10065 12641 10071
rect 12615 10033 12641 10039
rect 12839 10065 12865 10071
rect 13449 10039 13455 10065
rect 13481 10039 13487 10065
rect 14177 10039 14183 10065
rect 14209 10039 14215 10065
rect 12839 10033 12865 10039
rect 7519 10009 7545 10015
rect 2137 9983 2143 10009
rect 2169 9983 2175 10009
rect 7233 9983 7239 10009
rect 7265 9983 7271 10009
rect 7401 9983 7407 10009
rect 7433 9983 7439 10009
rect 7519 9977 7545 9983
rect 7687 10009 7713 10015
rect 7687 9977 7713 9983
rect 8023 10009 8049 10015
rect 10095 10009 10121 10015
rect 8801 9983 8807 10009
rect 8833 9983 8839 10009
rect 9137 9983 9143 10009
rect 9169 9983 9175 10009
rect 9697 9983 9703 10009
rect 9729 9983 9735 10009
rect 8023 9977 8049 9983
rect 10095 9977 10121 9983
rect 10375 10009 10401 10015
rect 10375 9977 10401 9983
rect 10823 10009 10849 10015
rect 10823 9977 10849 9983
rect 10935 10009 10961 10015
rect 10935 9977 10961 9983
rect 11103 10009 11129 10015
rect 12783 10009 12809 10015
rect 11265 9983 11271 10009
rect 11297 9983 11303 10009
rect 11881 9983 11887 10009
rect 11913 9983 11919 10009
rect 11993 9983 11999 10009
rect 12025 9983 12031 10009
rect 11103 9977 11129 9983
rect 12783 9977 12809 9983
rect 12895 10009 12921 10015
rect 13785 9983 13791 10009
rect 13817 9983 13823 10009
rect 18825 9983 18831 10009
rect 18857 9983 18863 10009
rect 12895 9977 12921 9983
rect 7295 9953 7321 9959
rect 7295 9921 7321 9927
rect 7743 9953 7769 9959
rect 13119 9953 13145 9959
rect 9921 9927 9927 9953
rect 9953 9927 9959 9953
rect 15241 9927 15247 9953
rect 15273 9927 15279 9953
rect 7743 9921 7769 9927
rect 13119 9921 13145 9927
rect 967 9897 993 9903
rect 967 9865 993 9871
rect 6903 9897 6929 9903
rect 6903 9865 6929 9871
rect 20007 9897 20033 9903
rect 20007 9865 20033 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 9473 9703 9479 9729
rect 9505 9703 9511 9729
rect 11657 9703 11663 9729
rect 11689 9703 11695 9729
rect 8807 9673 8833 9679
rect 13735 9673 13761 9679
rect 4993 9647 4999 9673
rect 5025 9647 5031 9673
rect 7177 9647 7183 9673
rect 7209 9647 7215 9673
rect 10873 9647 10879 9673
rect 10905 9647 10911 9673
rect 8807 9641 8833 9647
rect 13735 9641 13761 9647
rect 7239 9617 7265 9623
rect 6057 9591 6063 9617
rect 6089 9591 6095 9617
rect 6393 9591 6399 9617
rect 6425 9591 6431 9617
rect 7239 9585 7265 9591
rect 7351 9617 7377 9623
rect 8695 9617 8721 9623
rect 9871 9617 9897 9623
rect 7457 9591 7463 9617
rect 7489 9591 7495 9617
rect 9305 9591 9311 9617
rect 9337 9591 9343 9617
rect 9473 9591 9479 9617
rect 9505 9591 9511 9617
rect 9697 9591 9703 9617
rect 9729 9591 9735 9617
rect 7351 9585 7377 9591
rect 8695 9585 8721 9591
rect 9871 9585 9897 9591
rect 9983 9617 10009 9623
rect 9983 9585 10009 9591
rect 10263 9617 10289 9623
rect 10263 9585 10289 9591
rect 10431 9617 10457 9623
rect 11495 9617 11521 9623
rect 12391 9617 12417 9623
rect 10929 9591 10935 9617
rect 10961 9591 10967 9617
rect 11097 9591 11103 9617
rect 11129 9591 11135 9617
rect 11601 9591 11607 9617
rect 11633 9591 11639 9617
rect 12105 9591 12111 9617
rect 12137 9591 12143 9617
rect 12217 9591 12223 9617
rect 12249 9591 12255 9617
rect 10431 9585 10457 9591
rect 11495 9585 11521 9591
rect 12391 9585 12417 9591
rect 12615 9617 12641 9623
rect 12615 9585 12641 9591
rect 13119 9617 13145 9623
rect 13119 9585 13145 9591
rect 13343 9617 13369 9623
rect 14575 9617 14601 9623
rect 13897 9591 13903 9617
rect 13929 9591 13935 9617
rect 13343 9585 13369 9591
rect 14575 9585 14601 9591
rect 14743 9617 14769 9623
rect 14743 9585 14769 9591
rect 12335 9561 12361 9567
rect 8409 9535 8415 9561
rect 8441 9535 8447 9561
rect 12335 9529 12361 9535
rect 12671 9561 12697 9567
rect 12671 9529 12697 9535
rect 13567 9561 13593 9567
rect 13567 9529 13593 9535
rect 14631 9561 14657 9567
rect 14631 9529 14657 9535
rect 6791 9505 6817 9511
rect 6791 9473 6817 9479
rect 7183 9505 7209 9511
rect 7183 9473 7209 9479
rect 8583 9505 8609 9511
rect 8583 9473 8609 9479
rect 8863 9505 8889 9511
rect 8863 9473 8889 9479
rect 8975 9505 9001 9511
rect 8975 9473 9001 9479
rect 9927 9505 9953 9511
rect 9927 9473 9953 9479
rect 10319 9505 10345 9511
rect 10319 9473 10345 9479
rect 12783 9505 12809 9511
rect 12783 9473 12809 9479
rect 13175 9505 13201 9511
rect 13175 9473 13201 9479
rect 13231 9505 13257 9511
rect 13231 9473 13257 9479
rect 13287 9505 13313 9511
rect 13287 9473 13313 9479
rect 13679 9505 13705 9511
rect 13679 9473 13705 9479
rect 13791 9505 13817 9511
rect 13791 9473 13817 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 7799 9337 7825 9343
rect 7799 9305 7825 9311
rect 10319 9337 10345 9343
rect 10991 9337 11017 9343
rect 10705 9311 10711 9337
rect 10737 9311 10743 9337
rect 11601 9311 11607 9337
rect 11633 9311 11639 9337
rect 10319 9305 10345 9311
rect 10991 9305 11017 9311
rect 10151 9281 10177 9287
rect 10151 9249 10177 9255
rect 10207 9281 10233 9287
rect 11377 9255 11383 9281
rect 11409 9255 11415 9281
rect 10207 9249 10233 9255
rect 7183 9225 7209 9231
rect 7743 9225 7769 9231
rect 7569 9199 7575 9225
rect 7601 9199 7607 9225
rect 7183 9193 7209 9199
rect 7743 9193 7769 9199
rect 7799 9225 7825 9231
rect 7799 9193 7825 9199
rect 8023 9225 8049 9231
rect 8023 9193 8049 9199
rect 9703 9225 9729 9231
rect 9703 9193 9729 9199
rect 9815 9225 9841 9231
rect 10431 9225 10457 9231
rect 9977 9199 9983 9225
rect 10009 9199 10015 9225
rect 9815 9193 9841 9199
rect 10431 9193 10457 9199
rect 10823 9225 10849 9231
rect 10823 9193 10849 9199
rect 10991 9225 11017 9231
rect 10991 9193 11017 9199
rect 11159 9225 11185 9231
rect 13063 9225 13089 9231
rect 11321 9199 11327 9225
rect 11353 9199 11359 9225
rect 11825 9199 11831 9225
rect 11857 9199 11863 9225
rect 12945 9199 12951 9225
rect 12977 9199 12983 9225
rect 11159 9193 11185 9199
rect 13063 9193 13089 9199
rect 13175 9225 13201 9231
rect 13281 9199 13287 9225
rect 13313 9199 13319 9225
rect 13729 9199 13735 9225
rect 13761 9199 13767 9225
rect 14121 9199 14127 9225
rect 14153 9199 14159 9225
rect 18825 9199 18831 9225
rect 18857 9199 18863 9225
rect 13175 9193 13201 9199
rect 7071 9169 7097 9175
rect 7071 9137 7097 9143
rect 7351 9169 7377 9175
rect 7351 9137 7377 9143
rect 7911 9169 7937 9175
rect 7911 9137 7937 9143
rect 9759 9169 9785 9175
rect 9759 9137 9785 9143
rect 11719 9169 11745 9175
rect 11719 9137 11745 9143
rect 13119 9169 13145 9175
rect 13119 9137 13145 9143
rect 13567 9169 13593 9175
rect 15185 9143 15191 9169
rect 15217 9143 15223 9169
rect 13567 9137 13593 9143
rect 10543 9113 10569 9119
rect 10543 9081 10569 9087
rect 20007 9113 20033 9119
rect 20007 9081 20033 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 6791 8945 6817 8951
rect 10039 8945 10065 8951
rect 9529 8919 9535 8945
rect 9561 8919 9567 8945
rect 6791 8913 6817 8919
rect 10039 8913 10065 8919
rect 14071 8945 14097 8951
rect 14071 8913 14097 8919
rect 967 8889 993 8895
rect 6735 8889 6761 8895
rect 4937 8863 4943 8889
rect 4969 8863 4975 8889
rect 6001 8863 6007 8889
rect 6033 8863 6039 8889
rect 967 8857 993 8863
rect 6735 8857 6761 8863
rect 9815 8889 9841 8895
rect 10767 8889 10793 8895
rect 20007 8889 20033 8895
rect 10257 8863 10263 8889
rect 10289 8863 10295 8889
rect 11265 8863 11271 8889
rect 11297 8863 11303 8889
rect 9815 8857 9841 8863
rect 10767 8857 10793 8863
rect 20007 8857 20033 8863
rect 8191 8833 8217 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 6393 8807 6399 8833
rect 6425 8807 6431 8833
rect 8191 8801 8217 8807
rect 8359 8833 8385 8839
rect 9703 8833 9729 8839
rect 9249 8807 9255 8833
rect 9281 8807 9287 8833
rect 8359 8801 8385 8807
rect 9703 8801 9729 8807
rect 9983 8833 10009 8839
rect 10375 8833 10401 8839
rect 10823 8833 10849 8839
rect 12055 8833 12081 8839
rect 10201 8807 10207 8833
rect 10233 8807 10239 8833
rect 10649 8807 10655 8833
rect 10681 8807 10687 8833
rect 10985 8807 10991 8833
rect 11017 8807 11023 8833
rect 11545 8807 11551 8833
rect 11577 8807 11583 8833
rect 11769 8807 11775 8833
rect 11801 8807 11807 8833
rect 9983 8801 10009 8807
rect 10375 8801 10401 8807
rect 10823 8801 10849 8807
rect 12055 8801 12081 8807
rect 13567 8833 13593 8839
rect 13567 8801 13593 8807
rect 13735 8833 13761 8839
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 13735 8801 13761 8807
rect 7911 8777 7937 8783
rect 7911 8745 7937 8751
rect 8247 8777 8273 8783
rect 13847 8777 13873 8783
rect 9361 8751 9367 8777
rect 9393 8751 9399 8777
rect 11153 8751 11159 8777
rect 11185 8751 11191 8777
rect 11881 8751 11887 8777
rect 11913 8751 11919 8777
rect 8247 8745 8273 8751
rect 13847 8745 13873 8751
rect 14015 8777 14041 8783
rect 14015 8745 14041 8751
rect 14071 8777 14097 8783
rect 14071 8745 14097 8751
rect 7015 8721 7041 8727
rect 7015 8689 7041 8695
rect 7743 8721 7769 8727
rect 7743 8689 7769 8695
rect 8303 8721 8329 8727
rect 8303 8689 8329 8695
rect 8415 8721 8441 8727
rect 8415 8689 8441 8695
rect 12223 8721 12249 8727
rect 12223 8689 12249 8695
rect 13735 8721 13761 8727
rect 13735 8689 13761 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 7799 8553 7825 8559
rect 7799 8521 7825 8527
rect 8751 8553 8777 8559
rect 8751 8521 8777 8527
rect 8807 8553 8833 8559
rect 8807 8521 8833 8527
rect 8919 8553 8945 8559
rect 13455 8553 13481 8559
rect 10481 8527 10487 8553
rect 10513 8527 10519 8553
rect 8919 8521 8945 8527
rect 13455 8521 13481 8527
rect 13847 8553 13873 8559
rect 13847 8521 13873 8527
rect 13959 8553 13985 8559
rect 13959 8521 13985 8527
rect 7407 8497 7433 8503
rect 7407 8465 7433 8471
rect 7967 8497 7993 8503
rect 7967 8465 7993 8471
rect 9871 8497 9897 8503
rect 9871 8465 9897 8471
rect 13567 8497 13593 8503
rect 13567 8465 13593 8471
rect 13623 8497 13649 8503
rect 13623 8465 13649 8471
rect 14015 8497 14041 8503
rect 14015 8465 14041 8471
rect 7575 8441 7601 8447
rect 8023 8441 8049 8447
rect 2137 8415 2143 8441
rect 2169 8415 2175 8441
rect 7737 8415 7743 8441
rect 7769 8415 7775 8441
rect 7575 8409 7601 8415
rect 8023 8409 8049 8415
rect 8135 8441 8161 8447
rect 8975 8441 9001 8447
rect 8241 8415 8247 8441
rect 8273 8415 8279 8441
rect 8135 8409 8161 8415
rect 8975 8409 9001 8415
rect 10039 8441 10065 8447
rect 10039 8409 10065 8415
rect 10319 8441 10345 8447
rect 18825 8415 18831 8441
rect 18857 8415 18863 8441
rect 10319 8409 10345 8415
rect 967 8385 993 8391
rect 967 8353 993 8359
rect 7631 8385 7657 8391
rect 7631 8353 7657 8359
rect 8863 8385 8889 8391
rect 19945 8359 19951 8385
rect 19977 8359 19983 8385
rect 8863 8353 8889 8359
rect 8241 8303 8247 8329
rect 8273 8303 8279 8329
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 10711 8161 10737 8167
rect 10711 8129 10737 8135
rect 11943 8161 11969 8167
rect 11943 8129 11969 8135
rect 20007 8105 20033 8111
rect 6729 8079 6735 8105
rect 6761 8079 6767 8105
rect 7793 8079 7799 8105
rect 7825 8079 7831 8105
rect 10201 8079 10207 8105
rect 10233 8079 10239 8105
rect 13225 8079 13231 8105
rect 13257 8079 13263 8105
rect 14289 8079 14295 8105
rect 14321 8079 14327 8105
rect 20007 8073 20033 8079
rect 9983 8049 10009 8055
rect 8129 8023 8135 8049
rect 8161 8023 8167 8049
rect 9983 8017 10009 8023
rect 10655 8049 10681 8055
rect 12167 8049 12193 8055
rect 14631 8049 14657 8055
rect 11769 8023 11775 8049
rect 11801 8023 11807 8049
rect 12889 8023 12895 8049
rect 12921 8023 12927 8049
rect 18825 8023 18831 8049
rect 18857 8023 18863 8049
rect 10655 8017 10681 8023
rect 12167 8017 12193 8023
rect 14631 8017 14657 8023
rect 12049 7967 12055 7993
rect 12081 7967 12087 7993
rect 8415 7937 8441 7943
rect 8415 7905 8441 7911
rect 11775 7937 11801 7943
rect 11775 7905 11801 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 8191 7769 8217 7775
rect 8191 7737 8217 7743
rect 10543 7769 10569 7775
rect 10543 7737 10569 7743
rect 12615 7769 12641 7775
rect 12615 7737 12641 7743
rect 14855 7769 14881 7775
rect 14855 7737 14881 7743
rect 6953 7687 6959 7713
rect 6985 7687 6991 7713
rect 8353 7687 8359 7713
rect 8385 7687 8391 7713
rect 13225 7687 13231 7713
rect 13257 7687 13263 7713
rect 14625 7687 14631 7713
rect 14657 7687 14663 7713
rect 10711 7657 10737 7663
rect 6561 7631 6567 7657
rect 6593 7631 6599 7657
rect 9361 7631 9367 7657
rect 9393 7631 9399 7657
rect 10711 7625 10737 7631
rect 10879 7657 10905 7663
rect 10879 7625 10905 7631
rect 11159 7657 11185 7663
rect 12889 7631 12895 7657
rect 12921 7631 12927 7657
rect 14513 7631 14519 7657
rect 14545 7631 14551 7657
rect 11159 7625 11185 7631
rect 9031 7601 9057 7607
rect 12671 7601 12697 7607
rect 8017 7575 8023 7601
rect 8049 7575 8055 7601
rect 9417 7575 9423 7601
rect 9449 7575 9455 7601
rect 14289 7575 14295 7601
rect 14321 7575 14327 7601
rect 9031 7569 9057 7575
rect 12671 7569 12697 7575
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 10145 7295 10151 7321
rect 10177 7295 10183 7321
rect 11713 7295 11719 7321
rect 11745 7295 11751 7321
rect 12777 7295 12783 7321
rect 12809 7295 12815 7321
rect 13063 7265 13089 7271
rect 8745 7239 8751 7265
rect 8777 7239 8783 7265
rect 11377 7239 11383 7265
rect 11409 7239 11415 7265
rect 13063 7233 13089 7239
rect 8135 7209 8161 7215
rect 9081 7183 9087 7209
rect 9113 7183 9119 7209
rect 8135 7177 8161 7183
rect 10375 7153 10401 7159
rect 10375 7121 10401 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 8919 6985 8945 6991
rect 8919 6953 8945 6959
rect 9087 6985 9113 6991
rect 9087 6953 9113 6959
rect 9809 6903 9815 6929
rect 9841 6903 9847 6929
rect 9193 6847 9199 6873
rect 9225 6847 9231 6873
rect 9473 6847 9479 6873
rect 9505 6847 9511 6873
rect 10873 6791 10879 6817
rect 10905 6791 10911 6817
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 8689 2143 8695 2169
rect 8721 2143 8727 2169
rect 9249 2087 9255 2113
rect 9281 2087 9287 2113
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 13063 1833 13089 1839
rect 13063 1801 13089 1807
rect 8521 1751 8527 1777
rect 8553 1751 8559 1777
rect 12609 1751 12615 1777
rect 12641 1751 12647 1777
rect 9031 1665 9057 1671
rect 9031 1633 9057 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9311 19111 9337 19137
rect 11215 19111 11241 19137
rect 12783 19111 12809 19137
rect 8807 18999 8833 19025
rect 10879 18999 10905 19025
rect 12279 18999 12305 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 11383 18719 11409 18745
rect 13119 18719 13145 18745
rect 10487 18607 10513 18633
rect 10935 18607 10961 18633
rect 12671 18607 12697 18633
rect 10039 18551 10065 18577
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 8695 18327 8721 18353
rect 11159 18327 11185 18353
rect 13063 18327 13089 18353
rect 8191 18215 8217 18241
rect 10655 18215 10681 18241
rect 12559 18215 12585 18241
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 20119 17319 20145 17345
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 10655 14295 10681 14321
rect 11103 14295 11129 14321
rect 10823 14239 10849 14265
rect 10991 14239 11017 14265
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 10767 14015 10793 14041
rect 7015 13903 7041 13929
rect 9311 13903 9337 13929
rect 7351 13847 7377 13873
rect 8415 13847 8441 13873
rect 8807 13847 8833 13873
rect 9143 13847 9169 13873
rect 9647 13847 9673 13873
rect 12727 13847 12753 13873
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 10207 13623 10233 13649
rect 13623 13623 13649 13649
rect 8191 13567 8217 13593
rect 8415 13567 8441 13593
rect 10039 13567 10065 13593
rect 10711 13567 10737 13593
rect 12335 13567 12361 13593
rect 20007 13567 20033 13593
rect 6735 13511 6761 13537
rect 8639 13511 8665 13537
rect 10935 13511 10961 13537
rect 12503 13511 12529 13537
rect 13119 13511 13145 13537
rect 13399 13511 13425 13537
rect 13567 13511 13593 13537
rect 18831 13511 18857 13537
rect 7127 13455 7153 13481
rect 8975 13455 9001 13481
rect 10263 13455 10289 13481
rect 11271 13455 11297 13481
rect 12671 13455 12697 13481
rect 12951 13455 12977 13481
rect 13063 13455 13089 13481
rect 13343 13455 13369 13481
rect 13623 13455 13649 13481
rect 13231 13399 13257 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 7687 13231 7713 13257
rect 8247 13231 8273 13257
rect 8751 13231 8777 13257
rect 9031 13231 9057 13257
rect 9367 13231 9393 13257
rect 9927 13231 9953 13257
rect 9983 13231 10009 13257
rect 10767 13231 10793 13257
rect 11271 13231 11297 13257
rect 11663 13231 11689 13257
rect 7799 13175 7825 13201
rect 7855 13175 7881 13201
rect 8639 13175 8665 13201
rect 8807 13175 8833 13201
rect 10879 13175 10905 13201
rect 11551 13175 11577 13201
rect 11775 13175 11801 13201
rect 7519 13119 7545 13145
rect 7575 13119 7601 13145
rect 8023 13119 8049 13145
rect 8135 13119 8161 13145
rect 8191 13119 8217 13145
rect 8359 13119 8385 13145
rect 9143 13119 9169 13145
rect 9815 13119 9841 13145
rect 10039 13119 10065 13145
rect 10151 13119 10177 13145
rect 10655 13119 10681 13145
rect 10991 13119 11017 13145
rect 11215 13119 11241 13145
rect 11439 13119 11465 13145
rect 12671 13119 12697 13145
rect 14295 13119 14321 13145
rect 18831 13119 18857 13145
rect 9423 13063 9449 13089
rect 10767 13063 10793 13089
rect 11495 13063 11521 13089
rect 13007 13063 13033 13089
rect 14071 13063 14097 13089
rect 20007 13007 20033 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 13231 12783 13257 12809
rect 14295 12783 14321 12809
rect 14631 12783 14657 12809
rect 8415 12727 8441 12753
rect 8583 12727 8609 12753
rect 12895 12727 12921 12753
rect 8527 12671 8553 12697
rect 12503 12671 12529 12697
rect 12559 12671 12585 12697
rect 12671 12615 12697 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 7687 12447 7713 12473
rect 11383 12447 11409 12473
rect 11047 12391 11073 12417
rect 11215 12391 11241 12417
rect 11271 12391 11297 12417
rect 6063 12335 6089 12361
rect 10711 12335 10737 12361
rect 10935 12335 10961 12361
rect 6399 12279 6425 12305
rect 7463 12279 7489 12305
rect 7967 12279 7993 12305
rect 10823 12279 10849 12305
rect 8023 12223 8049 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 7799 11999 7825 12025
rect 12111 11999 12137 12025
rect 13623 11999 13649 12025
rect 7855 11943 7881 11969
rect 8079 11943 8105 11969
rect 8359 11943 8385 11969
rect 8639 11943 8665 11969
rect 8863 11943 8889 11969
rect 10375 11943 10401 11969
rect 10655 11943 10681 11969
rect 13343 11943 13369 11969
rect 7519 11887 7545 11913
rect 8191 11887 8217 11913
rect 11047 11887 11073 11913
rect 7575 11831 7601 11857
rect 7743 11831 7769 11857
rect 8583 11831 8609 11857
rect 10207 11831 10233 11857
rect 12335 11831 12361 11857
rect 13455 11831 13481 11857
rect 13567 11831 13593 11857
rect 13623 11831 13649 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 7575 11663 7601 11689
rect 7911 11663 7937 11689
rect 8079 11663 8105 11689
rect 8303 11663 8329 11689
rect 10095 11663 10121 11689
rect 10319 11663 10345 11689
rect 10991 11663 11017 11689
rect 7407 11607 7433 11633
rect 7743 11607 7769 11633
rect 10599 11607 10625 11633
rect 10711 11607 10737 11633
rect 13679 11607 13705 11633
rect 5503 11551 5529 11577
rect 7295 11551 7321 11577
rect 9927 11551 9953 11577
rect 10431 11551 10457 11577
rect 10823 11551 10849 11577
rect 10879 11551 10905 11577
rect 13287 11551 13313 11577
rect 14967 11551 14993 11577
rect 18831 11551 18857 11577
rect 5839 11495 5865 11521
rect 6903 11495 6929 11521
rect 14743 11495 14769 11521
rect 8247 11439 8273 11465
rect 8415 11439 8441 11465
rect 10263 11439 10289 11465
rect 20007 11439 20033 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 7519 11271 7545 11297
rect 11103 11271 11129 11297
rect 7015 11215 7041 11241
rect 8415 11215 8441 11241
rect 10095 11215 10121 11241
rect 10319 11215 10345 11241
rect 14295 11215 14321 11241
rect 14911 11215 14937 11241
rect 20007 11215 20033 11241
rect 7351 11159 7377 11185
rect 7855 11159 7881 11185
rect 8583 11159 8609 11185
rect 9927 11159 9953 11185
rect 10991 11159 11017 11185
rect 11215 11159 11241 11185
rect 11887 11159 11913 11185
rect 12111 11159 12137 11185
rect 12895 11159 12921 11185
rect 14743 11159 14769 11185
rect 18831 11159 18857 11185
rect 7687 11103 7713 11129
rect 8863 11103 8889 11129
rect 10655 11103 10681 11129
rect 10823 11103 10849 11129
rect 11271 11103 11297 11129
rect 12391 11103 12417 11129
rect 13231 11103 13257 11129
rect 14575 11103 14601 11129
rect 14631 11103 14657 11129
rect 7463 11047 7489 11073
rect 8023 11047 8049 11073
rect 8191 11047 8217 11073
rect 9031 11047 9057 11073
rect 9311 11047 9337 11073
rect 9479 11047 9505 11073
rect 12167 11047 12193 11073
rect 12223 11047 12249 11073
rect 12559 11047 12585 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 9031 10879 9057 10905
rect 9535 10879 9561 10905
rect 12671 10879 12697 10905
rect 13287 10879 13313 10905
rect 14015 10879 14041 10905
rect 7463 10823 7489 10849
rect 7575 10823 7601 10849
rect 13119 10823 13145 10849
rect 7351 10767 7377 10793
rect 7687 10767 7713 10793
rect 7855 10767 7881 10793
rect 9703 10767 9729 10793
rect 12727 10767 12753 10793
rect 13231 10767 13257 10793
rect 13343 10767 13369 10793
rect 13455 10767 13481 10793
rect 13903 10767 13929 10793
rect 14071 10767 14097 10793
rect 8079 10711 8105 10737
rect 9255 10711 9281 10737
rect 11551 10711 11577 10737
rect 12671 10655 12697 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 967 10431 993 10457
rect 4999 10431 5025 10457
rect 6791 10431 6817 10457
rect 7855 10431 7881 10457
rect 10935 10431 10961 10457
rect 2143 10375 2169 10401
rect 6399 10375 6425 10401
rect 7519 10375 7545 10401
rect 10039 10375 10065 10401
rect 10991 10375 11017 10401
rect 11103 10375 11129 10401
rect 11551 10375 11577 10401
rect 6063 10319 6089 10345
rect 13063 10319 13089 10345
rect 7407 10263 7433 10289
rect 11439 10263 11465 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 7127 10095 7153 10121
rect 8751 10095 8777 10121
rect 9983 10095 10009 10121
rect 12279 10095 12305 10121
rect 13287 10095 13313 10121
rect 6903 10039 6929 10065
rect 6959 10039 6985 10065
rect 7799 10039 7825 10065
rect 9255 10039 9281 10065
rect 9927 10039 9953 10065
rect 10207 10039 10233 10065
rect 10319 10039 10345 10065
rect 10655 10039 10681 10065
rect 11047 10039 11073 10065
rect 11327 10039 11353 10065
rect 11663 10039 11689 10065
rect 12167 10039 12193 10065
rect 12335 10039 12361 10065
rect 12615 10039 12641 10065
rect 12839 10039 12865 10065
rect 13455 10039 13481 10065
rect 14183 10039 14209 10065
rect 2143 9983 2169 10009
rect 7239 9983 7265 10009
rect 7407 9983 7433 10009
rect 7519 9983 7545 10009
rect 7687 9983 7713 10009
rect 8023 9983 8049 10009
rect 8807 9983 8833 10009
rect 9143 9983 9169 10009
rect 9703 9983 9729 10009
rect 10095 9983 10121 10009
rect 10375 9983 10401 10009
rect 10823 9983 10849 10009
rect 10935 9983 10961 10009
rect 11103 9983 11129 10009
rect 11271 9983 11297 10009
rect 11887 9983 11913 10009
rect 11999 9983 12025 10009
rect 12783 9983 12809 10009
rect 12895 9983 12921 10009
rect 13791 9983 13817 10009
rect 18831 9983 18857 10009
rect 7295 9927 7321 9953
rect 7743 9927 7769 9953
rect 9927 9927 9953 9953
rect 13119 9927 13145 9953
rect 15247 9927 15273 9953
rect 967 9871 993 9897
rect 6903 9871 6929 9897
rect 20007 9871 20033 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 9479 9703 9505 9729
rect 11663 9703 11689 9729
rect 4999 9647 5025 9673
rect 7183 9647 7209 9673
rect 8807 9647 8833 9673
rect 10879 9647 10905 9673
rect 13735 9647 13761 9673
rect 6063 9591 6089 9617
rect 6399 9591 6425 9617
rect 7239 9591 7265 9617
rect 7351 9591 7377 9617
rect 7463 9591 7489 9617
rect 8695 9591 8721 9617
rect 9311 9591 9337 9617
rect 9479 9591 9505 9617
rect 9703 9591 9729 9617
rect 9871 9591 9897 9617
rect 9983 9591 10009 9617
rect 10263 9591 10289 9617
rect 10431 9591 10457 9617
rect 10935 9591 10961 9617
rect 11103 9591 11129 9617
rect 11495 9591 11521 9617
rect 11607 9591 11633 9617
rect 12111 9591 12137 9617
rect 12223 9591 12249 9617
rect 12391 9591 12417 9617
rect 12615 9591 12641 9617
rect 13119 9591 13145 9617
rect 13343 9591 13369 9617
rect 13903 9591 13929 9617
rect 14575 9591 14601 9617
rect 14743 9591 14769 9617
rect 8415 9535 8441 9561
rect 12335 9535 12361 9561
rect 12671 9535 12697 9561
rect 13567 9535 13593 9561
rect 14631 9535 14657 9561
rect 6791 9479 6817 9505
rect 7183 9479 7209 9505
rect 8583 9479 8609 9505
rect 8863 9479 8889 9505
rect 8975 9479 9001 9505
rect 9927 9479 9953 9505
rect 10319 9479 10345 9505
rect 12783 9479 12809 9505
rect 13175 9479 13201 9505
rect 13231 9479 13257 9505
rect 13287 9479 13313 9505
rect 13679 9479 13705 9505
rect 13791 9479 13817 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 7799 9311 7825 9337
rect 10319 9311 10345 9337
rect 10711 9311 10737 9337
rect 10991 9311 11017 9337
rect 11607 9311 11633 9337
rect 10151 9255 10177 9281
rect 10207 9255 10233 9281
rect 11383 9255 11409 9281
rect 7183 9199 7209 9225
rect 7575 9199 7601 9225
rect 7743 9199 7769 9225
rect 7799 9199 7825 9225
rect 8023 9199 8049 9225
rect 9703 9199 9729 9225
rect 9815 9199 9841 9225
rect 9983 9199 10009 9225
rect 10431 9199 10457 9225
rect 10823 9199 10849 9225
rect 10991 9199 11017 9225
rect 11159 9199 11185 9225
rect 11327 9199 11353 9225
rect 11831 9199 11857 9225
rect 12951 9199 12977 9225
rect 13063 9199 13089 9225
rect 13175 9199 13201 9225
rect 13287 9199 13313 9225
rect 13735 9199 13761 9225
rect 14127 9199 14153 9225
rect 18831 9199 18857 9225
rect 7071 9143 7097 9169
rect 7351 9143 7377 9169
rect 7911 9143 7937 9169
rect 9759 9143 9785 9169
rect 11719 9143 11745 9169
rect 13119 9143 13145 9169
rect 13567 9143 13593 9169
rect 15191 9143 15217 9169
rect 10543 9087 10569 9113
rect 20007 9087 20033 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 6791 8919 6817 8945
rect 9535 8919 9561 8945
rect 10039 8919 10065 8945
rect 14071 8919 14097 8945
rect 967 8863 993 8889
rect 4943 8863 4969 8889
rect 6007 8863 6033 8889
rect 6735 8863 6761 8889
rect 9815 8863 9841 8889
rect 10263 8863 10289 8889
rect 10767 8863 10793 8889
rect 11271 8863 11297 8889
rect 20007 8863 20033 8889
rect 2143 8807 2169 8833
rect 6399 8807 6425 8833
rect 8191 8807 8217 8833
rect 8359 8807 8385 8833
rect 9255 8807 9281 8833
rect 9703 8807 9729 8833
rect 9983 8807 10009 8833
rect 10207 8807 10233 8833
rect 10375 8807 10401 8833
rect 10655 8807 10681 8833
rect 10823 8807 10849 8833
rect 10991 8807 11017 8833
rect 11551 8807 11577 8833
rect 11775 8807 11801 8833
rect 12055 8807 12081 8833
rect 13567 8807 13593 8833
rect 13735 8807 13761 8833
rect 18831 8807 18857 8833
rect 7911 8751 7937 8777
rect 8247 8751 8273 8777
rect 9367 8751 9393 8777
rect 11159 8751 11185 8777
rect 11887 8751 11913 8777
rect 13847 8751 13873 8777
rect 14015 8751 14041 8777
rect 14071 8751 14097 8777
rect 7015 8695 7041 8721
rect 7743 8695 7769 8721
rect 8303 8695 8329 8721
rect 8415 8695 8441 8721
rect 12223 8695 12249 8721
rect 13735 8695 13761 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7799 8527 7825 8553
rect 8751 8527 8777 8553
rect 8807 8527 8833 8553
rect 8919 8527 8945 8553
rect 10487 8527 10513 8553
rect 13455 8527 13481 8553
rect 13847 8527 13873 8553
rect 13959 8527 13985 8553
rect 7407 8471 7433 8497
rect 7967 8471 7993 8497
rect 9871 8471 9897 8497
rect 13567 8471 13593 8497
rect 13623 8471 13649 8497
rect 14015 8471 14041 8497
rect 2143 8415 2169 8441
rect 7575 8415 7601 8441
rect 7743 8415 7769 8441
rect 8023 8415 8049 8441
rect 8135 8415 8161 8441
rect 8247 8415 8273 8441
rect 8975 8415 9001 8441
rect 10039 8415 10065 8441
rect 10319 8415 10345 8441
rect 18831 8415 18857 8441
rect 967 8359 993 8385
rect 7631 8359 7657 8385
rect 8863 8359 8889 8385
rect 19951 8359 19977 8385
rect 8247 8303 8273 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 10711 8135 10737 8161
rect 11943 8135 11969 8161
rect 6735 8079 6761 8105
rect 7799 8079 7825 8105
rect 10207 8079 10233 8105
rect 13231 8079 13257 8105
rect 14295 8079 14321 8105
rect 20007 8079 20033 8105
rect 8135 8023 8161 8049
rect 9983 8023 10009 8049
rect 10655 8023 10681 8049
rect 11775 8023 11801 8049
rect 12167 8023 12193 8049
rect 12895 8023 12921 8049
rect 14631 8023 14657 8049
rect 18831 8023 18857 8049
rect 12055 7967 12081 7993
rect 8415 7911 8441 7937
rect 11775 7911 11801 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 8191 7743 8217 7769
rect 10543 7743 10569 7769
rect 12615 7743 12641 7769
rect 14855 7743 14881 7769
rect 6959 7687 6985 7713
rect 8359 7687 8385 7713
rect 13231 7687 13257 7713
rect 14631 7687 14657 7713
rect 6567 7631 6593 7657
rect 9367 7631 9393 7657
rect 10711 7631 10737 7657
rect 10879 7631 10905 7657
rect 11159 7631 11185 7657
rect 12895 7631 12921 7657
rect 14519 7631 14545 7657
rect 8023 7575 8049 7601
rect 9031 7575 9057 7601
rect 9423 7575 9449 7601
rect 12671 7575 12697 7601
rect 14295 7575 14321 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 10151 7295 10177 7321
rect 11719 7295 11745 7321
rect 12783 7295 12809 7321
rect 8751 7239 8777 7265
rect 11383 7239 11409 7265
rect 13063 7239 13089 7265
rect 8135 7183 8161 7209
rect 9087 7183 9113 7209
rect 10375 7127 10401 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 8919 6959 8945 6985
rect 9087 6959 9113 6985
rect 9815 6903 9841 6929
rect 9199 6847 9225 6873
rect 9479 6847 9505 6873
rect 10879 6791 10905 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 8695 2143 8721 2169
rect 9255 2087 9281 2113
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 13063 1807 13089 1833
rect 8527 1751 8553 1777
rect 12615 1751 12641 1777
rect 9031 1639 9057 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8064 20600 8120 21000
rect 8736 20600 8792 21000
rect 10080 20600 10136 21000
rect 10416 20600 10472 21000
rect 10752 20600 10808 21000
rect 11088 20600 11144 21000
rect 11760 20600 11816 21000
rect 12096 20600 12152 21000
rect 12432 20600 12488 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 8078 18354 8106 20600
rect 8750 19138 8778 20600
rect 8750 19105 8778 19110
rect 9310 19138 9338 19143
rect 9310 19091 9338 19110
rect 8806 19025 8834 19031
rect 8806 18999 8807 19025
rect 8833 18999 8834 19025
rect 8078 18321 8106 18326
rect 8694 18354 8722 18359
rect 8694 18307 8722 18326
rect 8190 18241 8218 18247
rect 8190 18215 8191 18241
rect 8217 18215 8218 18241
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 7014 13929 7042 13935
rect 7014 13903 7015 13929
rect 7041 13903 7042 13929
rect 5782 13818 5810 13823
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 5502 11746 5530 11751
rect 5502 11577 5530 11718
rect 5502 11551 5503 11577
rect 5529 11551 5530 11577
rect 5502 11545 5530 11551
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 5782 10906 5810 13790
rect 6734 13594 6762 13599
rect 6734 13537 6762 13566
rect 6734 13511 6735 13537
rect 6761 13511 6762 13537
rect 6734 13505 6762 13511
rect 7014 13594 7042 13903
rect 7350 13874 7378 13879
rect 7350 13873 7546 13874
rect 7350 13847 7351 13873
rect 7377 13847 7546 13873
rect 7350 13846 7546 13847
rect 7350 13841 7378 13846
rect 6174 12474 6202 12479
rect 6062 12446 6174 12474
rect 6062 12361 6090 12446
rect 6174 12441 6202 12446
rect 6846 12474 6874 12479
rect 6062 12335 6063 12361
rect 6089 12335 6090 12361
rect 6062 11746 6090 12335
rect 6398 12306 6426 12311
rect 6398 12259 6426 12278
rect 6062 11713 6090 11718
rect 5782 10873 5810 10878
rect 5838 11521 5866 11527
rect 5838 11495 5839 11521
rect 5865 11495 5866 11521
rect 5838 10850 5866 11495
rect 6846 11410 6874 12446
rect 7014 12474 7042 13566
rect 7126 13482 7154 13487
rect 7126 13481 7266 13482
rect 7126 13455 7127 13481
rect 7153 13455 7266 13481
rect 7126 13454 7266 13455
rect 7126 13449 7154 13454
rect 7238 13202 7266 13454
rect 7518 13426 7546 13846
rect 8190 13594 8218 18215
rect 8806 15974 8834 18999
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 10038 18578 10066 18583
rect 10094 18578 10122 20600
rect 10038 18577 10122 18578
rect 10038 18551 10039 18577
rect 10065 18551 10122 18577
rect 10038 18550 10122 18551
rect 10038 18545 10066 18550
rect 10430 18354 10458 20600
rect 10766 18746 10794 20600
rect 11102 19138 11130 20600
rect 11214 19138 11242 19143
rect 11102 19137 11242 19138
rect 11102 19111 11215 19137
rect 11241 19111 11242 19137
rect 11102 19110 11242 19111
rect 11214 19105 11242 19110
rect 11774 19138 11802 20600
rect 11774 19105 11802 19110
rect 10878 19026 10906 19031
rect 10878 19025 11018 19026
rect 10878 18999 10879 19025
rect 10905 18999 11018 19025
rect 10878 18998 11018 18999
rect 10878 18993 10906 18998
rect 10766 18713 10794 18718
rect 10430 18321 10458 18326
rect 10486 18633 10514 18639
rect 10486 18607 10487 18633
rect 10513 18607 10514 18633
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 8414 15946 8834 15974
rect 8414 13874 8442 15946
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 10038 14042 10066 14047
rect 9310 13929 9338 13935
rect 9310 13903 9311 13929
rect 9337 13903 9338 13929
rect 8806 13874 8834 13879
rect 8414 13873 8610 13874
rect 8414 13847 8415 13873
rect 8441 13847 8610 13873
rect 8414 13846 8610 13847
rect 8414 13841 8442 13846
rect 8582 13818 8610 13846
rect 8582 13790 8778 13818
rect 8414 13594 8442 13599
rect 8190 13593 8274 13594
rect 8190 13567 8191 13593
rect 8217 13567 8274 13593
rect 8190 13566 8274 13567
rect 8190 13561 8218 13566
rect 7518 13398 7714 13426
rect 7686 13257 7714 13398
rect 7686 13231 7687 13257
rect 7713 13231 7714 13257
rect 7686 13225 7714 13231
rect 8246 13257 8274 13566
rect 8414 13547 8442 13566
rect 8638 13594 8666 13599
rect 8638 13537 8666 13566
rect 8638 13511 8639 13537
rect 8665 13511 8666 13537
rect 8638 13505 8666 13511
rect 8246 13231 8247 13257
rect 8273 13231 8274 13257
rect 8246 13225 8274 13231
rect 8750 13257 8778 13790
rect 8806 13594 8834 13846
rect 9142 13874 9170 13879
rect 9310 13874 9338 13903
rect 9142 13873 9310 13874
rect 9142 13847 9143 13873
rect 9169 13847 9310 13873
rect 9142 13846 9310 13847
rect 9142 13841 9170 13846
rect 9310 13841 9338 13846
rect 9646 13873 9674 13879
rect 9646 13847 9647 13873
rect 9673 13847 9674 13873
rect 9646 13650 9674 13847
rect 9646 13617 9674 13622
rect 9814 13818 9842 13823
rect 8806 13561 8834 13566
rect 8974 13481 9002 13487
rect 8974 13455 8975 13481
rect 9001 13455 9002 13481
rect 8750 13231 8751 13257
rect 8777 13231 8778 13257
rect 8750 13225 8778 13231
rect 8806 13426 8834 13431
rect 7238 13174 7322 13202
rect 7294 13146 7322 13174
rect 7798 13201 7826 13207
rect 7798 13175 7799 13201
rect 7825 13175 7826 13201
rect 7518 13146 7546 13151
rect 7294 13145 7546 13146
rect 7294 13119 7519 13145
rect 7545 13119 7546 13145
rect 7294 13118 7546 13119
rect 7518 13113 7546 13118
rect 7574 13146 7602 13151
rect 7574 13099 7602 13118
rect 7798 12866 7826 13175
rect 7854 13202 7882 13207
rect 7854 13155 7882 13174
rect 8638 13202 8666 13207
rect 8638 13155 8666 13174
rect 8806 13201 8834 13398
rect 8974 13258 9002 13455
rect 8974 13225 9002 13230
rect 9030 13426 9058 13431
rect 9030 13257 9058 13398
rect 9030 13231 9031 13257
rect 9057 13231 9058 13257
rect 9030 13225 9058 13231
rect 9366 13258 9394 13263
rect 9814 13258 9842 13790
rect 10038 13593 10066 14014
rect 10486 14042 10514 18607
rect 10934 18633 10962 18639
rect 10934 18607 10935 18633
rect 10961 18607 10962 18633
rect 10654 18241 10682 18247
rect 10654 18215 10655 18241
rect 10681 18215 10682 18241
rect 10654 14322 10682 18215
rect 10934 15106 10962 18607
rect 10822 15078 10962 15106
rect 10766 14322 10794 14327
rect 10654 14321 10766 14322
rect 10654 14295 10655 14321
rect 10681 14295 10766 14321
rect 10654 14294 10766 14295
rect 10654 14289 10682 14294
rect 10486 14009 10514 14014
rect 10710 14042 10738 14047
rect 10598 13874 10626 13879
rect 10626 13846 10682 13874
rect 10598 13841 10626 13846
rect 10206 13650 10234 13655
rect 10206 13603 10234 13622
rect 10038 13567 10039 13593
rect 10065 13567 10066 13593
rect 10038 13561 10066 13567
rect 10654 13594 10682 13846
rect 10710 13706 10738 14014
rect 10766 14041 10794 14294
rect 10822 14265 10850 15078
rect 10822 14239 10823 14265
rect 10849 14239 10850 14265
rect 10822 14233 10850 14239
rect 10990 14265 11018 18998
rect 11382 18746 11410 18751
rect 11382 18699 11410 18718
rect 12110 18746 12138 20600
rect 12110 18713 12138 18718
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 11158 18354 11186 18359
rect 11158 18307 11186 18326
rect 12278 15974 12306 18999
rect 12446 18354 12474 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 13118 18746 13146 18751
rect 13118 18699 13146 18718
rect 12446 18321 12474 18326
rect 12670 18633 12698 18639
rect 12670 18607 12671 18633
rect 12697 18607 12698 18633
rect 12558 18241 12586 18247
rect 12558 18215 12559 18241
rect 12585 18215 12586 18241
rect 12558 15974 12586 18215
rect 12110 15946 12306 15974
rect 12502 15946 12586 15974
rect 11102 14322 11130 14327
rect 11102 14275 11130 14294
rect 10990 14239 10991 14265
rect 11017 14239 11018 14265
rect 10990 14233 11018 14239
rect 10766 14015 10767 14041
rect 10793 14015 10794 14041
rect 10766 13818 10794 14015
rect 10766 13785 10794 13790
rect 10710 13678 10794 13706
rect 10710 13594 10738 13599
rect 10654 13593 10738 13594
rect 10654 13567 10711 13593
rect 10737 13567 10738 13593
rect 10654 13566 10738 13567
rect 10710 13561 10738 13566
rect 10262 13482 10290 13487
rect 10094 13481 10290 13482
rect 10094 13455 10263 13481
rect 10289 13455 10290 13481
rect 10094 13454 10290 13455
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9926 13258 9954 13263
rect 9814 13257 9954 13258
rect 9814 13231 9927 13257
rect 9953 13231 9954 13257
rect 9814 13230 9954 13231
rect 9366 13211 9394 13230
rect 9926 13225 9954 13230
rect 9982 13258 10010 13263
rect 10094 13258 10122 13454
rect 10262 13449 10290 13454
rect 9982 13257 10122 13258
rect 9982 13231 9983 13257
rect 10009 13231 10122 13257
rect 9982 13230 10122 13231
rect 10766 13257 10794 13678
rect 10766 13231 10767 13257
rect 10793 13231 10794 13257
rect 9982 13225 10010 13230
rect 10766 13225 10794 13231
rect 10934 13537 10962 13543
rect 10934 13511 10935 13537
rect 10961 13511 10962 13537
rect 8806 13175 8807 13201
rect 8833 13175 8834 13201
rect 8806 13169 8834 13175
rect 10654 13202 10682 13207
rect 10878 13202 10906 13207
rect 8022 13146 8050 13151
rect 7798 12833 7826 12838
rect 7910 13145 8050 13146
rect 7910 13119 8023 13145
rect 8049 13119 8050 13145
rect 7910 13118 8050 13119
rect 7910 12586 7938 13118
rect 8022 13113 8050 13118
rect 8134 13145 8162 13151
rect 8134 13119 8135 13145
rect 8161 13119 8162 13145
rect 7014 12441 7042 12446
rect 7630 12558 7938 12586
rect 8078 12866 8106 12871
rect 7462 12305 7490 12311
rect 7462 12279 7463 12305
rect 7489 12279 7490 12305
rect 7462 12250 7490 12279
rect 7462 12217 7490 12222
rect 7518 11914 7546 11919
rect 7294 11913 7546 11914
rect 7294 11887 7519 11913
rect 7545 11887 7546 11913
rect 7294 11886 7546 11887
rect 7294 11634 7322 11886
rect 7518 11881 7546 11886
rect 7574 11857 7602 11863
rect 7574 11831 7575 11857
rect 7601 11831 7602 11857
rect 7574 11690 7602 11831
rect 7518 11689 7602 11690
rect 7518 11663 7575 11689
rect 7601 11663 7602 11689
rect 7518 11662 7602 11663
rect 6902 11606 7322 11634
rect 6902 11521 6930 11606
rect 7294 11577 7322 11606
rect 7294 11551 7295 11577
rect 7321 11551 7322 11577
rect 7294 11545 7322 11551
rect 7350 11634 7378 11639
rect 6902 11495 6903 11521
rect 6929 11495 6930 11521
rect 6902 11489 6930 11495
rect 5838 10817 5866 10822
rect 6790 11382 7042 11410
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 966 10457 994 10463
rect 966 10431 967 10457
rect 993 10431 994 10457
rect 966 10122 994 10431
rect 4998 10457 5026 10463
rect 4998 10431 4999 10457
rect 5025 10431 5026 10457
rect 2142 10402 2170 10407
rect 2142 10355 2170 10374
rect 4998 10346 5026 10431
rect 6790 10458 6818 11382
rect 7014 11241 7042 11382
rect 7014 11215 7015 11241
rect 7041 11215 7042 11241
rect 7014 11209 7042 11215
rect 7350 11185 7378 11606
rect 7406 11633 7434 11639
rect 7406 11607 7407 11633
rect 7433 11607 7434 11633
rect 7406 11466 7434 11607
rect 7406 11433 7434 11438
rect 7518 11297 7546 11662
rect 7574 11643 7602 11662
rect 7518 11271 7519 11297
rect 7545 11271 7546 11297
rect 7518 11265 7546 11271
rect 7350 11159 7351 11185
rect 7377 11159 7378 11185
rect 7350 11153 7378 11159
rect 7462 11074 7490 11079
rect 7630 11074 7658 12558
rect 7686 12474 7714 12479
rect 7686 12427 7714 12446
rect 7798 12306 7826 12311
rect 7966 12306 7994 12311
rect 7798 12025 7826 12278
rect 7910 12305 7994 12306
rect 7910 12279 7967 12305
rect 7993 12279 7994 12305
rect 7910 12278 7994 12279
rect 7910 12250 7938 12278
rect 7966 12273 7994 12278
rect 7798 11999 7799 12025
rect 7825 11999 7826 12025
rect 7798 11993 7826 11999
rect 7854 12026 7882 12031
rect 7854 11969 7882 11998
rect 7854 11943 7855 11969
rect 7881 11943 7882 11969
rect 7854 11937 7882 11943
rect 7742 11858 7770 11863
rect 7462 11073 7546 11074
rect 7462 11047 7463 11073
rect 7489 11047 7546 11073
rect 7462 11046 7546 11047
rect 7462 11041 7490 11046
rect 6398 10401 6426 10407
rect 6398 10375 6399 10401
rect 6425 10375 6426 10401
rect 4998 10313 5026 10318
rect 6062 10345 6090 10351
rect 6062 10319 6063 10345
rect 6089 10319 6090 10345
rect 966 10089 994 10094
rect 6062 10122 6090 10319
rect 6062 10089 6090 10094
rect 4998 10066 5026 10071
rect 2142 10010 2170 10015
rect 2142 9963 2170 9982
rect 966 9898 994 9903
rect 966 9851 994 9870
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 4998 9673 5026 10038
rect 4998 9647 4999 9673
rect 5025 9647 5026 9673
rect 4998 9641 5026 9647
rect 6062 9618 6090 9623
rect 6062 9571 6090 9590
rect 6398 9617 6426 10375
rect 6398 9591 6399 9617
rect 6425 9591 6426 9617
rect 6398 9506 6426 9591
rect 6790 9506 6818 10430
rect 7350 10962 7378 10967
rect 7350 10793 7378 10934
rect 7462 10850 7490 10855
rect 7462 10803 7490 10822
rect 7350 10767 7351 10793
rect 7377 10767 7378 10793
rect 7126 10122 7154 10141
rect 7126 10089 7154 10094
rect 6902 10066 6930 10071
rect 6902 10019 6930 10038
rect 6958 10065 6986 10071
rect 6958 10039 6959 10065
rect 6985 10039 6986 10065
rect 6958 10010 6986 10039
rect 6958 9977 6986 9982
rect 7238 10066 7266 10071
rect 7238 10009 7266 10038
rect 7238 9983 7239 10009
rect 7265 9983 7266 10009
rect 6902 9898 6930 9903
rect 6902 9851 6930 9870
rect 7238 9786 7266 9983
rect 7350 10010 7378 10767
rect 7518 10794 7546 11046
rect 7630 11041 7658 11046
rect 7686 11857 7770 11858
rect 7686 11831 7743 11857
rect 7769 11831 7770 11857
rect 7686 11830 7770 11831
rect 7686 11129 7714 11830
rect 7742 11825 7770 11830
rect 7910 11689 7938 12222
rect 8022 12249 8050 12255
rect 8022 12223 8023 12249
rect 8049 12223 8050 12249
rect 8022 11970 8050 12223
rect 8022 11937 8050 11942
rect 8078 11969 8106 12838
rect 8078 11943 8079 11969
rect 8105 11943 8106 11969
rect 8078 11937 8106 11943
rect 8134 12698 8162 13119
rect 8190 13146 8218 13151
rect 8190 13099 8218 13118
rect 8358 13146 8386 13151
rect 8358 12978 8386 13118
rect 9142 13146 9170 13151
rect 9142 13099 9170 13118
rect 9814 13146 9842 13151
rect 9814 13099 9842 13118
rect 10038 13145 10066 13151
rect 10038 13119 10039 13145
rect 10065 13119 10066 13145
rect 9422 13090 9450 13095
rect 9422 13043 9450 13062
rect 8358 12950 8498 12978
rect 8414 12866 8442 12871
rect 8414 12753 8442 12838
rect 8414 12727 8415 12753
rect 8441 12727 8442 12753
rect 8414 12721 8442 12727
rect 7910 11663 7911 11689
rect 7937 11663 7938 11689
rect 7910 11657 7938 11663
rect 8078 11690 8106 11695
rect 8078 11643 8106 11662
rect 7742 11634 7770 11639
rect 7742 11587 7770 11606
rect 8134 11242 8162 12670
rect 8190 12026 8218 12031
rect 8190 11914 8218 11998
rect 8358 11970 8386 11975
rect 8302 11942 8358 11970
rect 8190 11913 8274 11914
rect 8190 11887 8191 11913
rect 8217 11887 8274 11913
rect 8190 11886 8274 11887
rect 8190 11881 8218 11886
rect 8246 11578 8274 11886
rect 8302 11689 8330 11942
rect 8358 11923 8386 11942
rect 8470 11858 8498 12950
rect 8582 12754 8610 12759
rect 8582 12707 8610 12726
rect 10038 12754 10066 13119
rect 10150 13146 10178 13151
rect 10150 13099 10178 13118
rect 10654 13145 10682 13174
rect 10654 13119 10655 13145
rect 10681 13119 10682 13145
rect 10654 13113 10682 13119
rect 10822 13201 10906 13202
rect 10822 13175 10879 13201
rect 10905 13175 10906 13201
rect 10822 13174 10906 13175
rect 10822 13146 10850 13174
rect 10878 13169 10906 13174
rect 10766 13090 10794 13095
rect 10766 13043 10794 13062
rect 8526 12698 8554 12703
rect 8526 12651 8554 12670
rect 10038 12642 10066 12726
rect 10038 12614 10178 12642
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 10094 12474 10122 12479
rect 8638 11970 8666 11975
rect 8638 11923 8666 11942
rect 8862 11970 8890 11975
rect 8862 11969 8946 11970
rect 8862 11943 8863 11969
rect 8889 11943 8946 11969
rect 8862 11942 8946 11943
rect 8862 11937 8890 11942
rect 8582 11858 8610 11863
rect 8470 11857 8610 11858
rect 8470 11831 8583 11857
rect 8609 11831 8610 11857
rect 8470 11830 8610 11831
rect 8582 11825 8610 11830
rect 8302 11663 8303 11689
rect 8329 11663 8330 11689
rect 8302 11657 8330 11663
rect 8806 11690 8834 11695
rect 8246 11550 8330 11578
rect 7854 11214 8162 11242
rect 8246 11465 8274 11471
rect 8246 11439 8247 11465
rect 8273 11439 8274 11465
rect 7854 11185 7882 11214
rect 7854 11159 7855 11185
rect 7881 11159 7882 11185
rect 7854 11153 7882 11159
rect 7686 11103 7687 11129
rect 7713 11103 7714 11129
rect 7686 10962 7714 11103
rect 7686 10929 7714 10934
rect 7574 10850 7602 10855
rect 7574 10803 7602 10822
rect 7462 10626 7490 10631
rect 7406 10289 7434 10295
rect 7406 10263 7407 10289
rect 7433 10263 7434 10289
rect 7406 10094 7434 10263
rect 7406 10061 7434 10066
rect 7406 10010 7434 10015
rect 7350 10009 7434 10010
rect 7350 9983 7407 10009
rect 7433 9983 7434 10009
rect 7350 9982 7434 9983
rect 7294 9954 7322 9959
rect 7294 9907 7322 9926
rect 6398 9505 6818 9506
rect 6398 9479 6791 9505
rect 6817 9479 6818 9505
rect 6398 9478 6818 9479
rect 6006 9338 6034 9343
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 966 8890 994 8895
rect 966 8843 994 8862
rect 4942 8890 4970 8895
rect 4942 8843 4970 8862
rect 6006 8889 6034 9310
rect 6006 8863 6007 8889
rect 6033 8863 6034 8889
rect 6006 8857 6034 8863
rect 2142 8834 2170 8839
rect 2142 8787 2170 8806
rect 6398 8833 6426 9478
rect 6790 9473 6818 9478
rect 7126 9758 7266 9786
rect 7070 9170 7098 9175
rect 6790 9169 7098 9170
rect 6790 9143 7071 9169
rect 7097 9143 7098 9169
rect 6790 9142 7098 9143
rect 6790 8945 6818 9142
rect 7070 9137 7098 9142
rect 6790 8919 6791 8945
rect 6817 8919 6818 8945
rect 6790 8913 6818 8919
rect 6734 8890 6762 8895
rect 6734 8843 6762 8862
rect 6398 8807 6399 8833
rect 6425 8807 6426 8833
rect 966 8442 994 8447
rect 966 8385 994 8414
rect 2142 8442 2170 8447
rect 6398 8442 6426 8807
rect 7014 8721 7042 8727
rect 7014 8695 7015 8721
rect 7041 8695 7042 8721
rect 7014 8442 7042 8695
rect 7126 8554 7154 9758
rect 7182 9673 7210 9679
rect 7182 9647 7183 9673
rect 7209 9647 7210 9673
rect 7182 9618 7210 9647
rect 7182 9585 7210 9590
rect 7238 9617 7266 9758
rect 7238 9591 7239 9617
rect 7265 9591 7266 9617
rect 7238 9585 7266 9591
rect 7350 9898 7378 9903
rect 7350 9617 7378 9870
rect 7350 9591 7351 9617
rect 7377 9591 7378 9617
rect 7350 9585 7378 9591
rect 7182 9505 7210 9511
rect 7182 9479 7183 9505
rect 7209 9479 7210 9505
rect 7182 9450 7210 9479
rect 7406 9450 7434 9982
rect 7462 9617 7490 10598
rect 7518 10401 7546 10766
rect 7518 10375 7519 10401
rect 7545 10375 7546 10401
rect 7518 10369 7546 10375
rect 7686 10793 7714 10799
rect 7686 10767 7687 10793
rect 7713 10767 7714 10793
rect 7686 10122 7714 10767
rect 7854 10794 7882 10799
rect 7854 10747 7882 10766
rect 7854 10458 7882 10463
rect 7854 10411 7882 10430
rect 7462 9591 7463 9617
rect 7489 9591 7490 9617
rect 7462 9585 7490 9591
rect 7518 10009 7546 10015
rect 7518 9983 7519 10009
rect 7545 9983 7546 10009
rect 7182 9422 7434 9450
rect 7518 9338 7546 9983
rect 7686 10009 7714 10094
rect 7798 10346 7826 10351
rect 7798 10065 7826 10318
rect 7798 10039 7799 10065
rect 7825 10039 7826 10065
rect 7798 10033 7826 10039
rect 7686 9983 7687 10009
rect 7713 9983 7714 10009
rect 7518 9310 7658 9338
rect 7182 9282 7210 9287
rect 7182 9225 7210 9254
rect 7182 9199 7183 9225
rect 7209 9199 7210 9225
rect 7182 9193 7210 9199
rect 7574 9225 7602 9231
rect 7574 9199 7575 9225
rect 7601 9199 7602 9225
rect 7350 9170 7378 9175
rect 7574 9170 7602 9199
rect 7350 9169 7602 9170
rect 7350 9143 7351 9169
rect 7377 9143 7602 9169
rect 7350 9142 7602 9143
rect 7350 9137 7378 9142
rect 7630 8946 7658 9310
rect 7686 9282 7714 9983
rect 7742 9954 7770 9959
rect 7742 9907 7770 9926
rect 7686 9249 7714 9254
rect 7742 9674 7770 9679
rect 7742 9225 7770 9646
rect 7910 9562 7938 11214
rect 8246 11186 8274 11439
rect 8134 11158 8274 11186
rect 8022 11074 8050 11079
rect 8134 11074 8162 11158
rect 7910 9529 7938 9534
rect 7966 11073 8162 11074
rect 7966 11047 8023 11073
rect 8049 11047 8162 11073
rect 7966 11046 8162 11047
rect 8190 11074 8218 11079
rect 7798 9338 7826 9343
rect 7798 9291 7826 9310
rect 7742 9199 7743 9225
rect 7769 9199 7770 9225
rect 7742 9193 7770 9199
rect 7798 9226 7826 9231
rect 7798 9179 7826 9198
rect 7910 9170 7938 9175
rect 7126 8521 7154 8526
rect 7406 8918 7658 8946
rect 7406 8497 7434 8918
rect 7630 8722 7658 8918
rect 7854 9169 7938 9170
rect 7854 9143 7911 9169
rect 7937 9143 7938 9169
rect 7854 9142 7938 9143
rect 7742 8722 7770 8727
rect 7854 8722 7882 9142
rect 7910 9137 7938 9142
rect 7630 8721 7882 8722
rect 7630 8695 7743 8721
rect 7769 8695 7882 8721
rect 7630 8694 7882 8695
rect 7742 8689 7770 8694
rect 7406 8471 7407 8497
rect 7433 8471 7434 8497
rect 7406 8465 7434 8471
rect 7574 8666 7602 8671
rect 7126 8442 7154 8447
rect 6398 8414 7042 8442
rect 7070 8414 7126 8442
rect 2142 8395 2170 8414
rect 966 8359 967 8385
rect 993 8359 994 8385
rect 966 8353 994 8359
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 6566 7658 6594 7663
rect 6678 7658 6706 8414
rect 6734 8330 6762 8335
rect 6734 8105 6762 8302
rect 6734 8079 6735 8105
rect 6761 8079 6762 8105
rect 6734 8073 6762 8079
rect 7070 8050 7098 8414
rect 7126 8409 7154 8414
rect 7574 8441 7602 8638
rect 7630 8610 7658 8615
rect 7630 8498 7658 8582
rect 7798 8553 7826 8559
rect 7798 8527 7799 8553
rect 7825 8527 7826 8553
rect 7630 8465 7658 8470
rect 7742 8498 7770 8503
rect 7574 8415 7575 8441
rect 7601 8415 7602 8441
rect 7574 8409 7602 8415
rect 7742 8441 7770 8470
rect 7742 8415 7743 8441
rect 7769 8415 7770 8441
rect 7742 8409 7770 8415
rect 7630 8386 7658 8391
rect 7630 8339 7658 8358
rect 7798 8105 7826 8527
rect 7854 8498 7882 8694
rect 7910 8778 7938 8783
rect 7966 8778 7994 11046
rect 8022 11041 8050 11046
rect 8190 11027 8218 11046
rect 8078 10737 8106 10743
rect 8078 10711 8079 10737
rect 8105 10711 8106 10737
rect 8022 10009 8050 10015
rect 8022 9983 8023 10009
rect 8049 9983 8050 10009
rect 8022 9954 8050 9983
rect 8022 9921 8050 9926
rect 8022 9562 8050 9567
rect 8022 9225 8050 9534
rect 8022 9199 8023 9225
rect 8049 9199 8050 9225
rect 8022 9193 8050 9199
rect 8078 9226 8106 10711
rect 8302 9618 8330 11550
rect 8414 11466 8442 11471
rect 8442 11438 8610 11466
rect 8414 11419 8442 11438
rect 8414 11241 8442 11247
rect 8414 11215 8415 11241
rect 8441 11215 8442 11241
rect 8414 10850 8442 11215
rect 8582 11242 8610 11438
rect 8582 11185 8610 11214
rect 8582 11159 8583 11185
rect 8609 11159 8610 11185
rect 8582 11153 8610 11159
rect 8806 11186 8834 11662
rect 8918 11634 8946 11942
rect 10094 11802 10122 12446
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 10094 11689 10122 11774
rect 10094 11663 10095 11689
rect 10121 11663 10122 11689
rect 10094 11657 10122 11663
rect 10150 11858 10178 12614
rect 10822 12474 10850 13118
rect 10934 12978 10962 13511
rect 11270 13481 11298 13487
rect 11270 13455 11271 13481
rect 11297 13455 11298 13481
rect 11270 13257 11298 13455
rect 11662 13426 11690 13431
rect 11270 13231 11271 13257
rect 11297 13231 11298 13257
rect 11270 13225 11298 13231
rect 11326 13230 11522 13258
rect 10822 12441 10850 12446
rect 10878 12950 10962 12978
rect 10990 13145 11018 13151
rect 10990 13119 10991 13145
rect 11017 13119 11018 13145
rect 10990 12978 11018 13119
rect 11214 13146 11242 13151
rect 11326 13146 11354 13230
rect 11214 13145 11354 13146
rect 11214 13119 11215 13145
rect 11241 13119 11354 13145
rect 11214 13118 11354 13119
rect 11438 13145 11466 13151
rect 11438 13119 11439 13145
rect 11465 13119 11466 13145
rect 11214 13113 11242 13118
rect 11438 12978 11466 13119
rect 11494 13089 11522 13230
rect 11662 13257 11690 13398
rect 11662 13231 11663 13257
rect 11689 13231 11690 13257
rect 11662 13225 11690 13231
rect 11550 13202 11578 13207
rect 11774 13202 11802 13207
rect 11550 13201 11634 13202
rect 11550 13175 11551 13201
rect 11577 13175 11634 13201
rect 11550 13174 11634 13175
rect 11550 13169 11578 13174
rect 11606 13146 11634 13174
rect 11774 13155 11802 13174
rect 11606 13118 11690 13146
rect 11494 13063 11495 13089
rect 11521 13063 11522 13089
rect 11494 13057 11522 13063
rect 10990 12950 11466 12978
rect 10710 12362 10738 12367
rect 10374 12361 10738 12362
rect 10374 12335 10711 12361
rect 10737 12335 10738 12361
rect 10374 12334 10738 12335
rect 10374 11970 10402 12334
rect 10710 12329 10738 12334
rect 10822 12305 10850 12311
rect 10822 12279 10823 12305
rect 10849 12279 10850 12305
rect 10318 11969 10402 11970
rect 10318 11943 10375 11969
rect 10401 11943 10402 11969
rect 10318 11942 10402 11943
rect 10206 11858 10234 11863
rect 10150 11857 10234 11858
rect 10150 11831 10207 11857
rect 10233 11831 10234 11857
rect 10150 11830 10234 11831
rect 8414 10346 8442 10822
rect 8414 10313 8442 10318
rect 8470 11130 8498 11135
rect 8302 9585 8330 9590
rect 8414 9562 8442 9567
rect 8414 9515 8442 9534
rect 8078 9002 8106 9198
rect 8078 8969 8106 8974
rect 7910 8777 7994 8778
rect 7910 8751 7911 8777
rect 7937 8751 7994 8777
rect 7910 8750 7994 8751
rect 8190 8833 8218 8839
rect 8190 8807 8191 8833
rect 8217 8807 8218 8833
rect 7910 8722 7938 8750
rect 7910 8689 7938 8694
rect 8134 8666 8162 8671
rect 7966 8498 7994 8503
rect 7854 8497 7994 8498
rect 7854 8471 7967 8497
rect 7993 8471 7994 8497
rect 7854 8470 7994 8471
rect 7966 8465 7994 8470
rect 8022 8442 8050 8447
rect 8022 8395 8050 8414
rect 8134 8442 8162 8638
rect 8134 8395 8162 8414
rect 7798 8079 7799 8105
rect 7825 8079 7826 8105
rect 7798 8073 7826 8079
rect 6958 8022 7098 8050
rect 8134 8049 8162 8055
rect 8134 8023 8135 8049
rect 8161 8023 8162 8049
rect 6958 7713 6986 8022
rect 6958 7687 6959 7713
rect 6985 7687 6986 7713
rect 6958 7681 6986 7687
rect 6566 7657 6678 7658
rect 6566 7631 6567 7657
rect 6593 7631 6678 7657
rect 6566 7630 6678 7631
rect 6566 7625 6594 7630
rect 6678 7625 6706 7630
rect 8134 7658 8162 8023
rect 8134 7625 8162 7630
rect 8190 7769 8218 8807
rect 8358 8834 8386 8839
rect 8470 8834 8498 11102
rect 8694 11074 8722 11079
rect 8694 9617 8722 11046
rect 8806 10962 8834 11158
rect 8862 11298 8890 11303
rect 8862 11130 8890 11270
rect 8862 11083 8890 11102
rect 8918 11074 8946 11606
rect 10150 11634 10178 11830
rect 10206 11825 10234 11830
rect 10318 11689 10346 11942
rect 10374 11937 10402 11942
rect 10654 11969 10682 11975
rect 10654 11943 10655 11969
rect 10681 11943 10682 11969
rect 10654 11858 10682 11943
rect 10654 11825 10682 11830
rect 10318 11663 10319 11689
rect 10345 11663 10346 11689
rect 10318 11657 10346 11663
rect 10598 11802 10626 11807
rect 9926 11578 9954 11583
rect 9814 11577 9954 11578
rect 9814 11551 9927 11577
rect 9953 11551 9954 11577
rect 9814 11550 9954 11551
rect 9030 11074 9058 11079
rect 9310 11074 9338 11079
rect 8918 11073 9338 11074
rect 8918 11047 9031 11073
rect 9057 11047 9311 11073
rect 9337 11047 9338 11073
rect 8918 11046 9338 11047
rect 9030 11041 9058 11046
rect 8806 10934 9058 10962
rect 9030 10905 9058 10934
rect 9030 10879 9031 10905
rect 9057 10879 9058 10905
rect 9030 10873 9058 10879
rect 9254 10737 9282 10743
rect 9254 10711 9255 10737
rect 9281 10711 9282 10737
rect 8806 10346 8834 10351
rect 8750 10122 8778 10127
rect 8750 10075 8778 10094
rect 8806 10009 8834 10318
rect 9254 10122 9282 10711
rect 9254 10065 9282 10094
rect 9254 10039 9255 10065
rect 9281 10039 9282 10065
rect 9254 10033 9282 10039
rect 8806 9983 8807 10009
rect 8833 9983 8834 10009
rect 8806 9977 8834 9983
rect 9142 10009 9170 10015
rect 9142 9983 9143 10009
rect 9169 9983 9170 10009
rect 8806 9674 8834 9679
rect 8806 9627 8834 9646
rect 8694 9591 8695 9617
rect 8721 9591 8722 9617
rect 8582 9505 8610 9511
rect 8582 9479 8583 9505
rect 8609 9479 8610 9505
rect 8582 9226 8610 9479
rect 8582 9193 8610 9198
rect 8694 9058 8722 9591
rect 8694 9025 8722 9030
rect 8862 9505 8890 9511
rect 8862 9479 8863 9505
rect 8889 9479 8890 9505
rect 8358 8833 8498 8834
rect 8358 8807 8359 8833
rect 8385 8807 8498 8833
rect 8358 8806 8498 8807
rect 8862 8834 8890 9479
rect 8974 9506 9002 9511
rect 8974 9459 9002 9478
rect 8358 8801 8386 8806
rect 8862 8801 8890 8806
rect 8918 9394 8946 9399
rect 8246 8778 8274 8783
rect 8246 8731 8274 8750
rect 8918 8778 8946 9366
rect 9142 9226 9170 9983
rect 9310 9617 9338 11046
rect 9478 11073 9506 11079
rect 9478 11047 9479 11073
rect 9505 11047 9506 11073
rect 9422 10458 9450 10463
rect 9422 10010 9450 10430
rect 9478 10122 9506 11047
rect 9534 10906 9562 10911
rect 9562 10878 9730 10906
rect 9534 10859 9562 10878
rect 9702 10793 9730 10878
rect 9702 10767 9703 10793
rect 9729 10767 9730 10793
rect 9702 10761 9730 10767
rect 9478 10094 9730 10122
rect 9478 10010 9506 10015
rect 9422 9982 9478 10010
rect 9478 9729 9506 9982
rect 9478 9703 9479 9729
rect 9505 9703 9506 9729
rect 9478 9697 9506 9703
rect 9702 10009 9730 10094
rect 9702 9983 9703 10009
rect 9729 9983 9730 10009
rect 9702 9730 9730 9983
rect 9814 9786 9842 11550
rect 9926 11545 9954 11550
rect 10094 11242 10122 11247
rect 10094 11195 10122 11214
rect 9926 11186 9954 11191
rect 9926 11139 9954 11158
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 10038 10402 10066 10407
rect 10038 10355 10066 10374
rect 10094 10290 10122 10295
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9982 10122 10010 10127
rect 9926 10066 9954 10085
rect 9982 10075 10010 10094
rect 9926 10033 9954 10038
rect 10094 10009 10122 10262
rect 10094 9983 10095 10009
rect 10121 9983 10122 10009
rect 9926 9954 9954 9959
rect 9926 9907 9954 9926
rect 9814 9758 10010 9786
rect 9310 9591 9311 9617
rect 9337 9591 9338 9617
rect 9310 9585 9338 9591
rect 9478 9617 9506 9623
rect 9478 9591 9479 9617
rect 9505 9591 9506 9617
rect 9478 9562 9506 9591
rect 9702 9617 9730 9702
rect 9702 9591 9703 9617
rect 9729 9591 9730 9617
rect 9702 9585 9730 9591
rect 9870 9618 9898 9637
rect 9870 9585 9898 9590
rect 9982 9617 10010 9758
rect 9982 9591 9983 9617
rect 10009 9591 10010 9617
rect 9478 9529 9506 9534
rect 9702 9506 9730 9511
rect 9926 9506 9954 9511
rect 9702 9338 9730 9478
rect 9814 9505 9954 9506
rect 9814 9479 9927 9505
rect 9953 9479 9954 9505
rect 9814 9478 9954 9479
rect 9982 9506 10010 9591
rect 10094 9618 10122 9983
rect 10150 9954 10178 11606
rect 10598 11633 10626 11774
rect 10598 11607 10599 11633
rect 10625 11607 10626 11633
rect 10598 11601 10626 11607
rect 10710 11634 10738 11639
rect 10710 11587 10738 11606
rect 10430 11578 10458 11583
rect 10430 11531 10458 11550
rect 10766 11578 10794 11583
rect 10262 11465 10290 11471
rect 10262 11439 10263 11465
rect 10289 11439 10290 11465
rect 10262 11242 10290 11439
rect 10262 11209 10290 11214
rect 10318 11241 10346 11247
rect 10318 11215 10319 11241
rect 10345 11215 10346 11241
rect 10318 11186 10346 11215
rect 10262 10962 10290 10967
rect 10206 10934 10262 10962
rect 10206 10065 10234 10934
rect 10262 10929 10290 10934
rect 10206 10039 10207 10065
rect 10233 10039 10234 10065
rect 10206 10033 10234 10039
rect 10262 10066 10290 10071
rect 10150 9926 10234 9954
rect 10094 9585 10122 9590
rect 10150 9786 10178 9791
rect 9982 9478 10122 9506
rect 9814 9394 9842 9478
rect 9926 9473 9954 9478
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9814 9361 9842 9366
rect 9702 9310 9786 9338
rect 9758 9282 9786 9310
rect 10038 9282 10066 9287
rect 9758 9254 9842 9282
rect 9702 9226 9730 9231
rect 9142 8946 9170 9198
rect 9142 8913 9170 8918
rect 9366 9225 9730 9226
rect 9366 9199 9703 9225
rect 9729 9199 9730 9225
rect 9366 9198 9730 9199
rect 8302 8721 8330 8727
rect 8302 8695 8303 8721
rect 8329 8695 8330 8721
rect 8246 8498 8274 8503
rect 8246 8441 8274 8470
rect 8246 8415 8247 8441
rect 8273 8415 8274 8441
rect 8246 8409 8274 8415
rect 8246 8330 8274 8335
rect 8302 8330 8330 8695
rect 8414 8721 8442 8727
rect 8414 8695 8415 8721
rect 8441 8695 8442 8721
rect 8414 8554 8442 8695
rect 8750 8722 8778 8727
rect 8470 8554 8498 8559
rect 8414 8526 8470 8554
rect 8470 8521 8498 8526
rect 8750 8553 8778 8694
rect 8750 8527 8751 8553
rect 8777 8527 8778 8553
rect 8750 8521 8778 8527
rect 8806 8554 8834 8559
rect 8806 8507 8834 8526
rect 8918 8553 8946 8750
rect 9254 8834 9282 8839
rect 8918 8527 8919 8553
rect 8945 8527 8946 8553
rect 8918 8521 8946 8527
rect 8974 8610 9002 8615
rect 8974 8441 9002 8582
rect 9254 8498 9282 8806
rect 9366 8778 9394 9198
rect 9702 9193 9730 9198
rect 9814 9225 9842 9254
rect 9814 9199 9815 9225
rect 9841 9199 9842 9225
rect 9814 9193 9842 9199
rect 9982 9226 10010 9231
rect 9982 9179 10010 9198
rect 9758 9170 9786 9175
rect 9758 9123 9786 9142
rect 9534 8946 9562 8951
rect 9534 8899 9562 8918
rect 10038 8945 10066 9254
rect 10094 9114 10122 9478
rect 10150 9338 10178 9758
rect 10206 9394 10234 9926
rect 10206 9361 10234 9366
rect 10262 9617 10290 10038
rect 10318 10065 10346 11158
rect 10654 11130 10682 11135
rect 10766 11130 10794 11550
rect 10822 11577 10850 12279
rect 10878 11858 10906 12950
rect 11214 12474 11242 12479
rect 11046 12418 11074 12423
rect 11046 12371 11074 12390
rect 11214 12417 11242 12446
rect 11382 12474 11410 12479
rect 11382 12427 11410 12446
rect 11214 12391 11215 12417
rect 11241 12391 11242 12417
rect 11214 12385 11242 12391
rect 11270 12418 11298 12423
rect 11270 12417 11354 12418
rect 11270 12391 11271 12417
rect 11297 12391 11354 12417
rect 11270 12390 11354 12391
rect 11270 12385 11298 12390
rect 10878 11825 10906 11830
rect 10934 12361 10962 12367
rect 10934 12335 10935 12361
rect 10961 12335 10962 12361
rect 10822 11551 10823 11577
rect 10849 11551 10850 11577
rect 10822 11545 10850 11551
rect 10878 11577 10906 11583
rect 10878 11551 10879 11577
rect 10905 11551 10906 11577
rect 10822 11130 10850 11135
rect 10766 11102 10822 11130
rect 10654 11083 10682 11102
rect 10822 11083 10850 11102
rect 10878 10962 10906 11551
rect 10878 10929 10906 10934
rect 10934 11298 10962 12335
rect 11046 11914 11074 11919
rect 10990 11913 11074 11914
rect 10990 11887 11047 11913
rect 11073 11887 11074 11913
rect 10990 11886 11074 11887
rect 10990 11689 11018 11886
rect 11046 11881 11074 11886
rect 10990 11663 10991 11689
rect 11017 11663 11018 11689
rect 10990 11657 11018 11663
rect 11102 11298 11130 11303
rect 10934 11297 11130 11298
rect 10934 11271 11103 11297
rect 11129 11271 11130 11297
rect 10934 11270 11130 11271
rect 10934 10458 10962 11270
rect 11102 11265 11130 11270
rect 10990 11186 11018 11191
rect 10990 11139 11018 11158
rect 11214 11185 11242 11191
rect 11214 11159 11215 11185
rect 11241 11159 11242 11185
rect 11214 10626 11242 11159
rect 10654 10457 10962 10458
rect 10654 10431 10935 10457
rect 10961 10431 10962 10457
rect 10654 10430 10962 10431
rect 10654 10178 10682 10430
rect 10934 10425 10962 10430
rect 11046 10598 11242 10626
rect 11270 11129 11298 11135
rect 11270 11103 11271 11129
rect 11297 11103 11298 11129
rect 10990 10402 11018 10407
rect 11046 10402 11074 10598
rect 11270 10570 11298 11103
rect 11326 11074 11354 12390
rect 11438 12362 11466 12950
rect 11326 11041 11354 11046
rect 11382 12334 11466 12362
rect 11270 10537 11298 10542
rect 10990 10401 11074 10402
rect 10990 10375 10991 10401
rect 11017 10375 11074 10401
rect 10990 10374 11074 10375
rect 11102 10402 11130 10407
rect 11102 10401 11186 10402
rect 11102 10375 11103 10401
rect 11129 10375 11186 10401
rect 11102 10374 11186 10375
rect 10934 10290 10962 10295
rect 10990 10290 11018 10374
rect 11102 10369 11130 10374
rect 10962 10262 11018 10290
rect 10934 10257 10962 10262
rect 11158 10234 11186 10374
rect 11158 10201 11186 10206
rect 10318 10039 10319 10065
rect 10345 10039 10346 10065
rect 10318 9674 10346 10039
rect 10430 10122 10458 10127
rect 10374 10010 10402 10015
rect 10374 9963 10402 9982
rect 10318 9641 10346 9646
rect 10262 9591 10263 9617
rect 10289 9591 10290 9617
rect 10262 9338 10290 9591
rect 10374 9618 10402 9623
rect 10318 9505 10346 9511
rect 10318 9479 10319 9505
rect 10345 9479 10346 9505
rect 10318 9450 10346 9479
rect 10318 9417 10346 9422
rect 10318 9338 10346 9343
rect 10262 9337 10346 9338
rect 10262 9311 10319 9337
rect 10345 9311 10346 9337
rect 10262 9310 10346 9311
rect 10150 9281 10178 9310
rect 10318 9305 10346 9310
rect 10150 9255 10151 9281
rect 10177 9255 10178 9281
rect 10150 9249 10178 9255
rect 10206 9281 10234 9287
rect 10206 9255 10207 9281
rect 10233 9255 10234 9281
rect 10206 9226 10234 9255
rect 10374 9226 10402 9590
rect 10430 9617 10458 10094
rect 10654 10065 10682 10150
rect 10654 10039 10655 10065
rect 10681 10039 10682 10065
rect 10654 10033 10682 10039
rect 11046 10065 11074 10071
rect 11046 10039 11047 10065
rect 11073 10039 11074 10065
rect 10822 10009 10850 10015
rect 10822 9983 10823 10009
rect 10849 9983 10850 10009
rect 10822 9786 10850 9983
rect 10934 10010 10962 10015
rect 10934 9963 10962 9982
rect 10822 9758 10962 9786
rect 10878 9674 10906 9679
rect 10878 9627 10906 9646
rect 10430 9591 10431 9617
rect 10457 9591 10458 9617
rect 10430 9585 10458 9591
rect 10934 9617 10962 9758
rect 10934 9591 10935 9617
rect 10961 9591 10962 9617
rect 10654 9506 10682 9511
rect 10206 9193 10234 9198
rect 10318 9198 10402 9226
rect 10430 9226 10458 9231
rect 10262 9170 10290 9175
rect 10262 9114 10290 9142
rect 10094 9086 10290 9114
rect 10038 8919 10039 8945
rect 10065 8919 10066 8945
rect 10038 8913 10066 8919
rect 9814 8890 9842 8895
rect 9702 8834 9730 8839
rect 9702 8787 9730 8806
rect 9366 8777 9450 8778
rect 9366 8751 9367 8777
rect 9393 8751 9450 8777
rect 9366 8750 9450 8751
rect 9366 8745 9394 8750
rect 9254 8465 9282 8470
rect 8974 8415 8975 8441
rect 9001 8415 9002 8441
rect 8974 8409 9002 8415
rect 9422 8442 9450 8750
rect 8862 8386 8890 8391
rect 8862 8339 8890 8358
rect 8246 8329 8330 8330
rect 8246 8303 8247 8329
rect 8273 8303 8330 8329
rect 8246 8302 8330 8303
rect 8246 8297 8274 8302
rect 8190 7743 8191 7769
rect 8217 7743 8218 7769
rect 8022 7601 8050 7607
rect 8022 7575 8023 7601
rect 8049 7575 8050 7601
rect 8022 7574 8050 7575
rect 8190 7602 8218 7743
rect 8414 7937 8442 7943
rect 8414 7911 8415 7937
rect 8441 7911 8442 7937
rect 8022 7546 8218 7574
rect 8358 7713 8386 7719
rect 8358 7687 8359 7713
rect 8385 7687 8386 7713
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 8134 7209 8162 7215
rect 8134 7183 8135 7209
rect 8161 7183 8162 7209
rect 8134 7154 8162 7183
rect 8190 7154 8218 7159
rect 8134 7126 8190 7154
rect 8190 7121 8218 7126
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 8078 2114 8106 2119
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8078 400 8106 2086
rect 8358 1778 8386 7687
rect 8414 7658 8442 7911
rect 8414 7154 8442 7630
rect 9366 7658 9394 7663
rect 9366 7611 9394 7630
rect 8414 7121 8442 7126
rect 8694 7602 8722 7607
rect 8694 2169 8722 7574
rect 9030 7601 9058 7607
rect 9030 7575 9031 7601
rect 9057 7575 9058 7601
rect 9030 7574 9058 7575
rect 9422 7601 9450 8414
rect 9814 8050 9842 8862
rect 10206 8890 10234 8895
rect 9982 8834 10010 8839
rect 10010 8806 10122 8834
rect 9982 8787 10010 8806
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9870 8498 9898 8503
rect 9870 8451 9898 8470
rect 10038 8442 10066 8447
rect 10094 8442 10122 8806
rect 10206 8833 10234 8862
rect 10262 8889 10290 9086
rect 10262 8863 10263 8889
rect 10289 8863 10290 8889
rect 10262 8857 10290 8863
rect 10206 8807 10207 8833
rect 10233 8807 10234 8833
rect 10206 8801 10234 8807
rect 10318 8722 10346 9198
rect 10430 9179 10458 9198
rect 10542 9114 10570 9119
rect 10486 9113 10570 9114
rect 10486 9087 10543 9113
rect 10569 9087 10570 9113
rect 10486 9086 10570 9087
rect 10374 8834 10402 8839
rect 10486 8834 10514 9086
rect 10542 9081 10570 9086
rect 10402 8806 10514 8834
rect 10374 8787 10402 8806
rect 10318 8694 10402 8722
rect 10318 8442 10346 8447
rect 10038 8441 10346 8442
rect 10038 8415 10039 8441
rect 10065 8415 10319 8441
rect 10345 8415 10346 8441
rect 10038 8414 10346 8415
rect 10038 8409 10066 8414
rect 9982 8050 10010 8055
rect 9814 8022 9982 8050
rect 9982 8003 10010 8022
rect 9422 7575 9423 7601
rect 9449 7575 9450 7601
rect 9030 7546 9226 7574
rect 9422 7569 9450 7575
rect 9814 7938 9842 7943
rect 8750 7265 8778 7271
rect 8750 7239 8751 7265
rect 8777 7239 8778 7265
rect 8750 7154 8778 7239
rect 9086 7209 9114 7215
rect 9086 7183 9087 7209
rect 9113 7183 9114 7209
rect 8918 7154 8946 7159
rect 8750 7126 8918 7154
rect 8918 6985 8946 7126
rect 8918 6959 8919 6985
rect 8945 6959 8946 6985
rect 8918 6953 8946 6959
rect 9086 6985 9114 7183
rect 9086 6959 9087 6985
rect 9113 6959 9114 6985
rect 9086 6953 9114 6959
rect 9198 6873 9226 7546
rect 9198 6847 9199 6873
rect 9225 6847 9226 6873
rect 9198 6841 9226 6847
rect 9478 7154 9506 7159
rect 9478 6873 9506 7126
rect 9814 6929 9842 7910
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 10094 7574 10122 8414
rect 10318 8409 10346 8414
rect 10206 8106 10234 8111
rect 10374 8106 10402 8694
rect 10486 8553 10514 8806
rect 10486 8527 10487 8553
rect 10513 8527 10514 8553
rect 10486 8521 10514 8527
rect 10654 8833 10682 9478
rect 10710 9338 10738 9343
rect 10710 9291 10738 9310
rect 10934 9282 10962 9591
rect 10990 9506 11018 9511
rect 10990 9337 11018 9478
rect 11046 9450 11074 10039
rect 11326 10066 11354 10071
rect 11326 10019 11354 10038
rect 11102 10009 11130 10015
rect 11270 10010 11298 10015
rect 11102 9983 11103 10009
rect 11129 9983 11130 10009
rect 11102 9786 11130 9983
rect 11102 9753 11130 9758
rect 11214 10009 11298 10010
rect 11214 9983 11271 10009
rect 11297 9983 11298 10009
rect 11214 9982 11298 9983
rect 11046 9417 11074 9422
rect 11102 9617 11130 9623
rect 11102 9591 11103 9617
rect 11129 9591 11130 9617
rect 10990 9311 10991 9337
rect 11017 9311 11018 9337
rect 10990 9305 11018 9311
rect 10934 9249 10962 9254
rect 10822 9225 10850 9231
rect 10822 9199 10823 9225
rect 10849 9199 10850 9225
rect 10822 9170 10850 9199
rect 10822 9137 10850 9142
rect 10990 9225 11018 9231
rect 10990 9199 10991 9225
rect 11017 9199 11018 9225
rect 10990 9058 11018 9199
rect 10990 9025 11018 9030
rect 11102 9226 11130 9591
rect 11214 9618 11242 9982
rect 11270 9977 11298 9982
rect 11382 9954 11410 12334
rect 11662 11802 11690 13118
rect 12110 12418 12138 15946
rect 12334 13594 12362 13599
rect 12502 13594 12530 15946
rect 12334 13593 12530 13594
rect 12334 13567 12335 13593
rect 12361 13567 12530 13593
rect 12334 13566 12530 13567
rect 12334 13454 12362 13566
rect 12502 13537 12530 13566
rect 12502 13511 12503 13537
rect 12529 13511 12530 13537
rect 12502 13505 12530 13511
rect 12278 13426 12362 13454
rect 12558 13482 12586 13487
rect 12278 13202 12306 13426
rect 12278 13169 12306 13174
rect 12110 12025 12138 12390
rect 12110 11999 12111 12025
rect 12137 11999 12138 12025
rect 12110 11993 12138 11999
rect 12502 12697 12530 12703
rect 12502 12671 12503 12697
rect 12529 12671 12530 12697
rect 12334 11858 12362 11863
rect 12502 11858 12530 12671
rect 12558 12697 12586 13454
rect 12670 13481 12698 18607
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 13062 18354 13090 18359
rect 13062 18307 13090 18326
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 20118 17345 20146 17351
rect 20118 17319 20119 17345
rect 20145 17319 20146 17345
rect 20118 17178 20146 17319
rect 20118 17145 20146 17150
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 12670 13455 12671 13481
rect 12697 13455 12698 13481
rect 12670 13449 12698 13455
rect 12726 13873 12754 13879
rect 12726 13847 12727 13873
rect 12753 13847 12754 13873
rect 12670 13146 12698 13151
rect 12726 13146 12754 13847
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 13622 13650 13650 13655
rect 13398 13649 13650 13650
rect 13398 13623 13623 13649
rect 13649 13623 13650 13649
rect 13398 13622 13650 13623
rect 13118 13538 13146 13543
rect 13118 13491 13146 13510
rect 13398 13537 13426 13622
rect 13622 13617 13650 13622
rect 20006 13593 20034 13599
rect 20006 13567 20007 13593
rect 20033 13567 20034 13593
rect 13398 13511 13399 13537
rect 13425 13511 13426 13537
rect 13398 13505 13426 13511
rect 13454 13538 13482 13543
rect 13566 13538 13594 13543
rect 13482 13537 13594 13538
rect 13482 13511 13567 13537
rect 13593 13511 13594 13537
rect 13482 13510 13594 13511
rect 13454 13505 13482 13510
rect 13566 13505 13594 13510
rect 13622 13538 13650 13543
rect 14406 13538 14434 13543
rect 12950 13482 12978 13487
rect 12950 13435 12978 13454
rect 13062 13482 13090 13487
rect 13062 13435 13090 13454
rect 13342 13481 13370 13487
rect 13342 13455 13343 13481
rect 13369 13455 13370 13481
rect 12698 13118 12754 13146
rect 13230 13425 13258 13431
rect 13230 13399 13231 13425
rect 13257 13399 13258 13425
rect 12670 12754 12698 13118
rect 13006 13089 13034 13095
rect 13006 13063 13007 13089
rect 13033 13063 13034 13089
rect 12894 12754 12922 12759
rect 12670 12753 12922 12754
rect 12670 12727 12895 12753
rect 12921 12727 12922 12753
rect 12670 12726 12922 12727
rect 12558 12671 12559 12697
rect 12585 12671 12586 12697
rect 12558 12665 12586 12671
rect 12670 12642 12698 12647
rect 12670 12595 12698 12614
rect 12894 11858 12922 12726
rect 13006 12642 13034 13063
rect 13230 12809 13258 13399
rect 13230 12783 13231 12809
rect 13257 12783 13258 12809
rect 13230 12777 13258 12783
rect 13006 12609 13034 12614
rect 13342 12474 13370 13455
rect 13622 13481 13650 13510
rect 14350 13510 14406 13538
rect 13622 13455 13623 13481
rect 13649 13455 13650 13481
rect 13622 13449 13650 13455
rect 14070 13482 14098 13487
rect 14070 13089 14098 13454
rect 14294 13146 14322 13151
rect 14294 13099 14322 13118
rect 14070 13063 14071 13089
rect 14097 13063 14098 13089
rect 14070 13034 14098 13063
rect 14070 13001 14098 13006
rect 14294 12810 14322 12815
rect 14350 12810 14378 13510
rect 14406 13505 14434 13510
rect 18830 13538 18858 13543
rect 18830 13491 18858 13510
rect 14294 12809 14378 12810
rect 14294 12783 14295 12809
rect 14321 12783 14378 12809
rect 14294 12782 14378 12783
rect 14630 13146 14658 13151
rect 14630 12809 14658 13118
rect 18830 13146 18858 13151
rect 18830 13099 18858 13118
rect 20006 13146 20034 13567
rect 20006 13113 20034 13118
rect 20006 13033 20034 13039
rect 20006 13007 20007 13033
rect 20033 13007 20034 13033
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 14630 12783 14631 12809
rect 14657 12783 14658 12809
rect 14294 12777 14322 12782
rect 14630 12777 14658 12783
rect 20006 12810 20034 13007
rect 20006 12777 20034 12782
rect 13342 11969 13370 12446
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 13622 12026 13650 12031
rect 13622 12025 13706 12026
rect 13622 11999 13623 12025
rect 13649 11999 13706 12025
rect 13622 11998 13706 11999
rect 13622 11993 13650 11998
rect 13342 11943 13343 11969
rect 13369 11943 13370 11969
rect 13342 11937 13370 11943
rect 12502 11830 12642 11858
rect 12334 11811 12362 11830
rect 11886 11802 11914 11807
rect 11662 11769 11690 11774
rect 11830 11774 11886 11802
rect 11550 10737 11578 10743
rect 11550 10711 11551 10737
rect 11577 10711 11578 10737
rect 11550 10402 11578 10711
rect 11550 10355 11578 10374
rect 11438 10290 11466 10295
rect 11438 10243 11466 10262
rect 11662 10066 11690 10071
rect 11662 10065 11746 10066
rect 11662 10039 11663 10065
rect 11689 10039 11746 10065
rect 11662 10038 11746 10039
rect 11662 10033 11690 10038
rect 11214 9338 11242 9590
rect 11326 9926 11410 9954
rect 11214 9305 11242 9310
rect 11270 9562 11298 9567
rect 10766 8890 10794 8895
rect 10766 8843 10794 8862
rect 10654 8807 10655 8833
rect 10681 8807 10682 8833
rect 10654 8162 10682 8807
rect 10822 8834 10850 8839
rect 10990 8834 11018 8839
rect 10850 8833 11018 8834
rect 10850 8807 10991 8833
rect 11017 8807 11018 8833
rect 10850 8806 11018 8807
rect 10822 8787 10850 8806
rect 10990 8801 11018 8806
rect 11102 8778 11130 9198
rect 11158 9225 11186 9231
rect 11158 9199 11159 9225
rect 11185 9199 11186 9225
rect 11158 9170 11186 9199
rect 11158 9137 11186 9142
rect 11270 8889 11298 9534
rect 11326 9225 11354 9926
rect 11494 9730 11522 9735
rect 11494 9617 11522 9702
rect 11662 9729 11690 9735
rect 11662 9703 11663 9729
rect 11689 9703 11690 9729
rect 11494 9591 11495 9617
rect 11521 9591 11522 9617
rect 11494 9585 11522 9591
rect 11606 9617 11634 9623
rect 11606 9591 11607 9617
rect 11633 9591 11634 9617
rect 11606 9562 11634 9591
rect 11606 9529 11634 9534
rect 11606 9338 11634 9343
rect 11606 9291 11634 9310
rect 11326 9199 11327 9225
rect 11353 9199 11354 9225
rect 11326 9002 11354 9199
rect 11326 8969 11354 8974
rect 11382 9281 11410 9287
rect 11382 9255 11383 9281
rect 11409 9255 11410 9281
rect 11270 8863 11271 8889
rect 11297 8863 11298 8889
rect 11158 8778 11186 8783
rect 11102 8777 11186 8778
rect 11102 8751 11159 8777
rect 11185 8751 11186 8777
rect 11102 8750 11186 8751
rect 10710 8162 10738 8167
rect 10654 8161 10738 8162
rect 10654 8135 10711 8161
rect 10737 8135 10738 8161
rect 10654 8134 10738 8135
rect 10206 8105 10402 8106
rect 10206 8079 10207 8105
rect 10233 8079 10402 8105
rect 10206 8078 10402 8079
rect 10206 7658 10234 8078
rect 10654 8050 10682 8055
rect 10542 8022 10654 8050
rect 10542 7769 10570 8022
rect 10654 8003 10682 8022
rect 10710 7938 10738 8134
rect 10710 7905 10738 7910
rect 10542 7743 10543 7769
rect 10569 7743 10570 7769
rect 10542 7737 10570 7743
rect 10206 7625 10234 7630
rect 10710 7658 10738 7663
rect 10878 7658 10906 7663
rect 10710 7657 10906 7658
rect 10710 7631 10711 7657
rect 10737 7631 10879 7657
rect 10905 7631 10906 7657
rect 10710 7630 10906 7631
rect 10710 7625 10738 7630
rect 10094 7546 10178 7574
rect 10150 7321 10178 7546
rect 10150 7295 10151 7321
rect 10177 7295 10178 7321
rect 10150 7289 10178 7295
rect 10374 7154 10402 7159
rect 10374 7107 10402 7126
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9814 6903 9815 6929
rect 9841 6903 9842 6929
rect 9814 6897 9842 6903
rect 9478 6847 9479 6873
rect 9505 6847 9506 6873
rect 9478 6841 9506 6847
rect 10878 6817 10906 7630
rect 11158 7657 11186 8750
rect 11270 8050 11298 8863
rect 11382 8890 11410 9255
rect 11662 9282 11690 9703
rect 11718 9338 11746 10038
rect 11830 9898 11858 11774
rect 11886 11769 11914 11774
rect 12110 11802 12138 11807
rect 11886 11298 11914 11303
rect 11886 11186 11914 11270
rect 11886 11185 11970 11186
rect 11886 11159 11887 11185
rect 11913 11159 11970 11185
rect 11886 11158 11970 11159
rect 11886 11153 11914 11158
rect 11942 10906 11970 11158
rect 12110 11185 12138 11774
rect 12110 11159 12111 11185
rect 12137 11159 12138 11185
rect 12110 11153 12138 11159
rect 11886 10346 11914 10351
rect 11886 10178 11914 10318
rect 11886 10009 11914 10150
rect 11886 9983 11887 10009
rect 11913 9983 11914 10009
rect 11886 9977 11914 9983
rect 11830 9870 11914 9898
rect 11718 9310 11802 9338
rect 11662 9254 11746 9282
rect 11718 9170 11746 9254
rect 11774 9226 11802 9310
rect 11830 9226 11858 9231
rect 11774 9225 11858 9226
rect 11774 9199 11831 9225
rect 11857 9199 11858 9225
rect 11774 9198 11858 9199
rect 11830 9193 11858 9198
rect 11718 9123 11746 9142
rect 11382 8857 11410 8862
rect 11718 8890 11746 8895
rect 11746 8862 11802 8890
rect 11718 8857 11746 8862
rect 11550 8834 11578 8839
rect 11550 8787 11578 8806
rect 11774 8833 11802 8862
rect 11774 8807 11775 8833
rect 11801 8807 11802 8833
rect 11774 8801 11802 8807
rect 11886 8777 11914 9870
rect 11886 8751 11887 8777
rect 11913 8751 11914 8777
rect 11886 8554 11914 8751
rect 11886 8521 11914 8526
rect 11942 8161 11970 10878
rect 12054 11130 12082 11135
rect 11998 10234 12026 10239
rect 11998 10009 12026 10206
rect 11998 9983 11999 10009
rect 12025 9983 12026 10009
rect 11998 9977 12026 9983
rect 12054 8834 12082 11102
rect 12390 11130 12418 11135
rect 12390 11083 12418 11102
rect 12166 11073 12194 11079
rect 12166 11047 12167 11073
rect 12193 11047 12194 11073
rect 12166 10850 12194 11047
rect 12166 10817 12194 10822
rect 12222 11073 12250 11079
rect 12222 11047 12223 11073
rect 12249 11047 12250 11073
rect 12222 10794 12250 11047
rect 12166 10626 12194 10631
rect 12166 10065 12194 10598
rect 12222 10290 12250 10766
rect 12558 11073 12586 11079
rect 12558 11047 12559 11073
rect 12585 11047 12586 11073
rect 12558 10738 12586 11047
rect 12334 10290 12362 10295
rect 12222 10262 12334 10290
rect 12278 10178 12306 10183
rect 12278 10121 12306 10150
rect 12278 10095 12279 10121
rect 12305 10095 12306 10121
rect 12278 10089 12306 10095
rect 12166 10039 12167 10065
rect 12193 10039 12194 10065
rect 12110 9618 12138 9623
rect 12110 9571 12138 9590
rect 12166 9338 12194 10039
rect 12334 10065 12362 10262
rect 12334 10039 12335 10065
rect 12361 10039 12362 10065
rect 12334 10033 12362 10039
rect 12558 9954 12586 10710
rect 12614 10682 12642 11830
rect 12894 11578 12922 11830
rect 13454 11857 13482 11863
rect 13454 11831 13455 11857
rect 13481 11831 13482 11857
rect 12894 11185 12922 11550
rect 13286 11578 13314 11583
rect 13286 11531 13314 11550
rect 12894 11159 12895 11185
rect 12921 11159 12922 11185
rect 12670 10906 12698 10911
rect 12670 10859 12698 10878
rect 12726 10794 12754 10799
rect 12726 10747 12754 10766
rect 12670 10682 12698 10687
rect 12614 10681 12698 10682
rect 12614 10655 12671 10681
rect 12697 10655 12698 10681
rect 12614 10654 12698 10655
rect 12670 10649 12698 10654
rect 12614 10570 12642 10575
rect 12614 10065 12642 10542
rect 12894 10346 12922 11159
rect 13230 11129 13258 11135
rect 13230 11103 13231 11129
rect 13257 11103 13258 11129
rect 13230 10906 13258 11103
rect 13342 10962 13370 10967
rect 13286 10906 13314 10911
rect 13230 10905 13314 10906
rect 13230 10879 13287 10905
rect 13313 10879 13314 10905
rect 13230 10878 13314 10879
rect 13286 10873 13314 10878
rect 13118 10850 13146 10855
rect 13146 10822 13202 10850
rect 13118 10803 13146 10822
rect 13062 10346 13090 10351
rect 12894 10345 13090 10346
rect 12894 10319 13063 10345
rect 13089 10319 13090 10345
rect 12894 10318 13090 10319
rect 12614 10039 12615 10065
rect 12641 10039 12642 10065
rect 12614 10033 12642 10039
rect 12782 10122 12810 10127
rect 12782 10010 12810 10094
rect 12838 10066 12866 10071
rect 12838 10019 12866 10038
rect 12334 9926 12586 9954
rect 12670 10009 12810 10010
rect 12670 9983 12783 10009
rect 12809 9983 12810 10009
rect 12670 9982 12810 9983
rect 12222 9730 12250 9735
rect 12222 9617 12250 9702
rect 12222 9591 12223 9617
rect 12249 9591 12250 9617
rect 12222 9585 12250 9591
rect 12334 9561 12362 9926
rect 12390 9618 12418 9623
rect 12390 9571 12418 9590
rect 12614 9618 12642 9623
rect 12614 9571 12642 9590
rect 12334 9535 12335 9561
rect 12361 9535 12362 9561
rect 12334 9529 12362 9535
rect 12670 9561 12698 9982
rect 12782 9977 12810 9982
rect 12894 10009 12922 10015
rect 12894 9983 12895 10009
rect 12921 9983 12922 10009
rect 12894 9618 12922 9983
rect 12894 9585 12922 9590
rect 13062 9954 13090 10318
rect 13118 9954 13146 9959
rect 13062 9953 13146 9954
rect 13062 9927 13119 9953
rect 13145 9927 13146 9953
rect 13062 9926 13146 9927
rect 12670 9535 12671 9561
rect 12697 9535 12698 9561
rect 12670 9529 12698 9535
rect 12782 9506 12810 9511
rect 12782 9505 12978 9506
rect 12782 9479 12783 9505
rect 12809 9479 12978 9505
rect 12782 9478 12978 9479
rect 12782 9473 12810 9478
rect 12166 9305 12194 9310
rect 12950 9225 12978 9478
rect 13006 9338 13034 9343
rect 13062 9338 13090 9926
rect 13118 9921 13146 9926
rect 13118 9618 13146 9623
rect 13174 9618 13202 10822
rect 13230 10793 13258 10799
rect 13230 10767 13231 10793
rect 13257 10767 13258 10793
rect 13230 10066 13258 10767
rect 13342 10793 13370 10934
rect 13454 10906 13482 11831
rect 13566 11857 13594 11863
rect 13566 11831 13567 11857
rect 13593 11831 13594 11857
rect 13566 10962 13594 11831
rect 13622 11857 13650 11863
rect 13622 11831 13623 11857
rect 13649 11831 13650 11857
rect 13622 11298 13650 11831
rect 13678 11633 13706 11998
rect 13678 11607 13679 11633
rect 13705 11607 13706 11633
rect 13678 11601 13706 11607
rect 14910 11578 14938 11583
rect 14966 11578 14994 11583
rect 14938 11577 14994 11578
rect 14938 11551 14967 11577
rect 14993 11551 14994 11577
rect 14938 11550 14994 11551
rect 14742 11522 14770 11527
rect 13622 11265 13650 11270
rect 14630 11494 14742 11522
rect 13566 10929 13594 10934
rect 14014 11242 14042 11247
rect 13342 10767 13343 10793
rect 13369 10767 13370 10793
rect 13286 10458 13314 10463
rect 13342 10458 13370 10767
rect 13398 10878 13482 10906
rect 14014 10905 14042 11214
rect 14294 11242 14322 11247
rect 14294 11195 14322 11214
rect 14014 10879 14015 10905
rect 14041 10879 14042 10905
rect 13398 10682 13426 10878
rect 14014 10873 14042 10879
rect 14574 11129 14602 11135
rect 14574 11103 14575 11129
rect 14601 11103 14602 11129
rect 13454 10794 13482 10799
rect 13902 10794 13930 10799
rect 13454 10793 13930 10794
rect 13454 10767 13455 10793
rect 13481 10767 13903 10793
rect 13929 10767 13930 10793
rect 13454 10766 13930 10767
rect 13454 10761 13482 10766
rect 13902 10761 13930 10766
rect 14070 10794 14098 10799
rect 14070 10747 14098 10766
rect 14574 10794 14602 11103
rect 14630 11129 14658 11494
rect 14742 11475 14770 11494
rect 14686 11298 14714 11303
rect 14686 11186 14714 11270
rect 14910 11241 14938 11550
rect 14966 11545 14994 11550
rect 18830 11578 18858 11583
rect 18830 11531 18858 11550
rect 20006 11466 20034 11471
rect 20006 11419 20034 11438
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 14910 11215 14911 11241
rect 14937 11215 14938 11241
rect 14910 11209 14938 11215
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 14742 11186 14770 11191
rect 14686 11185 14770 11186
rect 14686 11159 14743 11185
rect 14769 11159 14770 11185
rect 14686 11158 14770 11159
rect 14742 11153 14770 11158
rect 18830 11186 18858 11191
rect 18830 11139 18858 11158
rect 14630 11103 14631 11129
rect 14657 11103 14658 11129
rect 14630 11097 14658 11103
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 13398 10654 13650 10682
rect 13314 10430 13370 10458
rect 13286 10121 13314 10430
rect 13286 10095 13287 10121
rect 13313 10095 13314 10121
rect 13286 10089 13314 10095
rect 13454 10066 13482 10071
rect 13230 10033 13258 10038
rect 13342 10065 13482 10066
rect 13342 10039 13455 10065
rect 13481 10039 13482 10065
rect 13342 10038 13482 10039
rect 13118 9617 13202 9618
rect 13118 9591 13119 9617
rect 13145 9591 13202 9617
rect 13118 9590 13202 9591
rect 13342 9617 13370 10038
rect 13454 10033 13482 10038
rect 13622 9674 13650 10654
rect 13342 9591 13343 9617
rect 13369 9591 13370 9617
rect 13118 9585 13146 9590
rect 13174 9506 13202 9511
rect 13174 9459 13202 9478
rect 13230 9505 13258 9511
rect 13230 9479 13231 9505
rect 13257 9479 13258 9505
rect 13118 9338 13146 9343
rect 13062 9310 13118 9338
rect 13006 9282 13034 9310
rect 13118 9305 13146 9310
rect 13006 9254 13090 9282
rect 12950 9199 12951 9225
rect 12977 9199 12978 9225
rect 12950 9193 12978 9199
rect 13062 9225 13090 9254
rect 13062 9199 13063 9225
rect 13089 9199 13090 9225
rect 13062 9193 13090 9199
rect 13174 9225 13202 9231
rect 13174 9199 13175 9225
rect 13201 9199 13202 9225
rect 12054 8787 12082 8806
rect 13118 9169 13146 9175
rect 13118 9143 13119 9169
rect 13145 9143 13146 9169
rect 12222 8721 12250 8727
rect 12222 8695 12223 8721
rect 12249 8695 12250 8721
rect 12222 8498 12250 8695
rect 11942 8135 11943 8161
rect 11969 8135 11970 8161
rect 11942 8129 11970 8135
rect 12166 8470 12222 8498
rect 11270 8017 11298 8022
rect 11774 8050 11802 8069
rect 11774 8017 11802 8022
rect 12166 8049 12194 8470
rect 12222 8465 12250 8470
rect 12166 8023 12167 8049
rect 12193 8023 12194 8049
rect 12166 8017 12194 8023
rect 12894 8050 12922 8055
rect 12054 7994 12082 7999
rect 12054 7947 12082 7966
rect 12614 7994 12642 7999
rect 11158 7631 11159 7657
rect 11185 7631 11186 7657
rect 11158 7625 11186 7631
rect 11774 7937 11802 7943
rect 11774 7911 11775 7937
rect 11801 7911 11802 7937
rect 11774 7574 11802 7911
rect 12614 7769 12642 7966
rect 12614 7743 12615 7769
rect 12641 7743 12642 7769
rect 12614 7737 12642 7743
rect 12894 7657 12922 8022
rect 13118 7994 13146 9143
rect 13174 8554 13202 9199
rect 13230 9226 13258 9479
rect 13286 9505 13314 9511
rect 13286 9479 13287 9505
rect 13313 9479 13314 9505
rect 13286 9394 13314 9479
rect 13286 9361 13314 9366
rect 13230 9193 13258 9198
rect 13286 9226 13314 9231
rect 13342 9226 13370 9591
rect 13286 9225 13370 9226
rect 13286 9199 13287 9225
rect 13313 9199 13370 9225
rect 13286 9198 13370 9199
rect 13454 9646 13650 9674
rect 13734 10066 14210 10094
rect 13734 9673 13762 10066
rect 14182 10065 14210 10066
rect 14182 10039 14183 10065
rect 14209 10039 14210 10065
rect 14182 10033 14210 10039
rect 13734 9647 13735 9673
rect 13761 9647 13762 9673
rect 13454 9282 13482 9646
rect 13734 9641 13762 9647
rect 13790 10009 13818 10015
rect 13790 9983 13791 10009
rect 13817 9983 13818 10009
rect 13790 9618 13818 9983
rect 13902 9618 13930 9623
rect 13790 9590 13874 9618
rect 13566 9561 13594 9567
rect 13566 9535 13567 9561
rect 13593 9535 13594 9561
rect 13566 9282 13594 9535
rect 13678 9506 13706 9511
rect 13678 9459 13706 9478
rect 13790 9505 13818 9511
rect 13790 9479 13791 9505
rect 13817 9479 13818 9505
rect 13286 9058 13314 9198
rect 13454 9058 13482 9254
rect 13510 9254 13594 9282
rect 13734 9282 13762 9287
rect 13510 9170 13538 9254
rect 13734 9225 13762 9254
rect 13734 9199 13735 9225
rect 13761 9199 13762 9225
rect 13510 9137 13538 9142
rect 13566 9170 13594 9175
rect 13734 9170 13762 9199
rect 13566 9169 13762 9170
rect 13566 9143 13567 9169
rect 13593 9143 13762 9169
rect 13566 9142 13762 9143
rect 13566 9137 13594 9142
rect 13454 9030 13594 9058
rect 13286 9025 13314 9030
rect 13566 8833 13594 9030
rect 13566 8807 13567 8833
rect 13593 8807 13594 8833
rect 13566 8801 13594 8807
rect 13174 8521 13202 8526
rect 13230 8722 13258 8727
rect 13230 8105 13258 8694
rect 13622 8610 13650 9142
rect 13790 9058 13818 9479
rect 13846 9338 13874 9590
rect 13902 9571 13930 9590
rect 14574 9617 14602 10766
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 18830 10010 18858 10015
rect 18830 9963 18858 9982
rect 14574 9591 14575 9617
rect 14601 9591 14602 9617
rect 14574 9585 14602 9591
rect 14630 9954 14658 9959
rect 14630 9561 14658 9926
rect 15246 9954 15274 9959
rect 15246 9907 15274 9926
rect 20006 9897 20034 9903
rect 20006 9871 20007 9897
rect 20033 9871 20034 9897
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 20006 9786 20034 9871
rect 20006 9753 20034 9758
rect 14742 9618 14770 9623
rect 14742 9571 14770 9590
rect 14630 9535 14631 9561
rect 14657 9535 14658 9561
rect 14630 9529 14658 9535
rect 13846 9305 13874 9310
rect 14014 9394 14042 9399
rect 13734 8834 13762 8839
rect 13790 8834 13818 9030
rect 14014 8946 14042 9366
rect 14126 9226 14154 9231
rect 14126 9179 14154 9198
rect 18830 9226 18858 9231
rect 18830 9179 18858 9198
rect 15190 9170 15218 9175
rect 14070 8946 14098 8951
rect 14014 8945 14098 8946
rect 14014 8919 14071 8945
rect 14097 8919 14098 8945
rect 14014 8918 14098 8919
rect 14070 8913 14098 8918
rect 13734 8833 13818 8834
rect 13734 8807 13735 8833
rect 13761 8807 13818 8833
rect 13734 8806 13818 8807
rect 13958 8834 13986 8839
rect 13734 8801 13762 8806
rect 13846 8777 13874 8783
rect 13846 8751 13847 8777
rect 13873 8751 13874 8777
rect 13734 8722 13762 8727
rect 13734 8675 13762 8694
rect 13510 8582 13650 8610
rect 13454 8554 13482 8559
rect 13454 8507 13482 8526
rect 13510 8442 13538 8582
rect 13846 8553 13874 8751
rect 13846 8527 13847 8553
rect 13873 8527 13874 8553
rect 13846 8521 13874 8527
rect 13958 8553 13986 8806
rect 14294 8834 14322 8839
rect 13958 8527 13959 8553
rect 13985 8527 13986 8553
rect 13958 8521 13986 8527
rect 14014 8777 14042 8783
rect 14014 8751 14015 8777
rect 14041 8751 14042 8777
rect 13230 8079 13231 8105
rect 13257 8079 13258 8105
rect 13230 8073 13258 8079
rect 13398 8414 13538 8442
rect 13566 8497 13594 8503
rect 13566 8471 13567 8497
rect 13593 8471 13594 8497
rect 13566 8442 13594 8471
rect 13622 8498 13650 8503
rect 13622 8451 13650 8470
rect 14014 8498 14042 8751
rect 14070 8778 14098 8783
rect 14070 8731 14098 8750
rect 14014 8451 14042 8470
rect 13398 8050 13426 8414
rect 13566 8409 13594 8414
rect 14294 8105 14322 8806
rect 15190 8778 15218 9142
rect 20006 9114 20034 9119
rect 20006 9067 20034 9086
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 15190 8745 15218 8750
rect 14294 8079 14295 8105
rect 14321 8079 14322 8105
rect 14294 8073 14322 8079
rect 14518 8442 14546 8447
rect 13398 8017 13426 8022
rect 13118 7966 13202 7994
rect 13174 7714 13202 7966
rect 13230 7714 13258 7719
rect 13174 7713 13258 7714
rect 13174 7687 13231 7713
rect 13257 7687 13258 7713
rect 13174 7686 13258 7687
rect 13230 7681 13258 7686
rect 14518 7658 14546 8414
rect 18830 8442 18858 8447
rect 18830 8395 18858 8414
rect 20006 8442 20034 8863
rect 20006 8409 20034 8414
rect 19950 8385 19978 8391
rect 19950 8359 19951 8385
rect 19977 8359 19978 8385
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 19950 8106 19978 8359
rect 19950 8073 19978 8078
rect 20006 8105 20034 8111
rect 20006 8079 20007 8105
rect 20033 8079 20034 8105
rect 14630 8050 14658 8055
rect 14630 8003 14658 8022
rect 14854 8050 14882 8055
rect 14854 7769 14882 8022
rect 14854 7743 14855 7769
rect 14881 7743 14882 7769
rect 14854 7737 14882 7743
rect 18830 8049 18858 8055
rect 18830 8023 18831 8049
rect 18857 8023 18858 8049
rect 14630 7714 14658 7719
rect 14630 7667 14658 7686
rect 18830 7714 18858 8023
rect 20006 7770 20034 8079
rect 20006 7737 20034 7742
rect 18830 7681 18858 7686
rect 12894 7631 12895 7657
rect 12921 7631 12922 7657
rect 11718 7546 11802 7574
rect 12670 7601 12698 7607
rect 12670 7575 12671 7601
rect 12697 7575 12698 7601
rect 11718 7321 11746 7546
rect 11718 7295 11719 7321
rect 11745 7295 11746 7321
rect 11718 7289 11746 7295
rect 12670 7322 12698 7575
rect 12782 7322 12810 7327
rect 12670 7321 12810 7322
rect 12670 7295 12783 7321
rect 12809 7295 12810 7321
rect 12670 7294 12810 7295
rect 11382 7266 11410 7271
rect 11382 7219 11410 7238
rect 10878 6791 10879 6817
rect 10905 6791 10906 6817
rect 10878 6785 10906 6791
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 12782 4214 12810 7294
rect 12894 7266 12922 7631
rect 14294 7657 14546 7658
rect 14294 7631 14519 7657
rect 14545 7631 14546 7657
rect 14294 7630 14546 7631
rect 14294 7601 14322 7630
rect 14518 7625 14546 7630
rect 14294 7575 14295 7601
rect 14321 7575 14322 7601
rect 14294 7569 14322 7575
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 12894 7233 12922 7238
rect 13062 7266 13090 7271
rect 13062 7219 13090 7238
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 12614 4186 12810 4214
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 8694 2143 8695 2169
rect 8721 2143 8722 2169
rect 8694 2137 8722 2143
rect 9254 2114 9282 2119
rect 9254 2067 9282 2086
rect 12446 1834 12474 1839
rect 8526 1778 8554 1783
rect 8358 1777 8554 1778
rect 8358 1751 8527 1777
rect 8553 1751 8554 1777
rect 8358 1750 8554 1751
rect 8526 1745 8554 1750
rect 8582 1722 8610 1727
rect 8582 490 8610 1694
rect 9030 1722 9058 1727
rect 9030 1665 9058 1694
rect 9030 1639 9031 1665
rect 9057 1639 9058 1665
rect 9030 1633 9058 1639
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 8414 462 8610 490
rect 8414 400 8442 462
rect 12446 400 12474 1806
rect 12614 1777 12642 4186
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 13062 1834 13090 1839
rect 13062 1787 13090 1806
rect 12614 1751 12615 1777
rect 12641 1751 12642 1777
rect 12614 1745 12642 1751
rect 8064 0 8120 400
rect 8400 0 8456 400
rect 12432 0 12488 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 8750 19110 8778 19138
rect 9310 19137 9338 19138
rect 9310 19111 9311 19137
rect 9311 19111 9337 19137
rect 9337 19111 9338 19137
rect 9310 19110 9338 19111
rect 8078 18326 8106 18354
rect 8694 18353 8722 18354
rect 8694 18327 8695 18353
rect 8695 18327 8721 18353
rect 8721 18327 8722 18353
rect 8694 18326 8722 18327
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 5782 13790 5810 13818
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 5502 11718 5530 11746
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 6734 13566 6762 13594
rect 7014 13566 7042 13594
rect 6174 12446 6202 12474
rect 6846 12446 6874 12474
rect 6398 12305 6426 12306
rect 6398 12279 6399 12305
rect 6399 12279 6425 12305
rect 6425 12279 6426 12305
rect 6398 12278 6426 12279
rect 6062 11718 6090 11746
rect 5782 10878 5810 10906
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 11774 19110 11802 19138
rect 10766 18718 10794 18746
rect 10430 18326 10458 18354
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 10038 14014 10066 14042
rect 8806 13873 8834 13874
rect 8806 13847 8807 13873
rect 8807 13847 8833 13873
rect 8833 13847 8834 13873
rect 8806 13846 8834 13847
rect 8414 13593 8442 13594
rect 8414 13567 8415 13593
rect 8415 13567 8441 13593
rect 8441 13567 8442 13593
rect 8414 13566 8442 13567
rect 8638 13566 8666 13594
rect 9310 13846 9338 13874
rect 9646 13622 9674 13650
rect 9814 13790 9842 13818
rect 8806 13566 8834 13594
rect 8806 13398 8834 13426
rect 7574 13145 7602 13146
rect 7574 13119 7575 13145
rect 7575 13119 7601 13145
rect 7601 13119 7602 13145
rect 7574 13118 7602 13119
rect 7854 13201 7882 13202
rect 7854 13175 7855 13201
rect 7855 13175 7881 13201
rect 7881 13175 7882 13201
rect 7854 13174 7882 13175
rect 8638 13201 8666 13202
rect 8638 13175 8639 13201
rect 8639 13175 8665 13201
rect 8665 13175 8666 13201
rect 8638 13174 8666 13175
rect 8974 13230 9002 13258
rect 9030 13398 9058 13426
rect 9366 13257 9394 13258
rect 9366 13231 9367 13257
rect 9367 13231 9393 13257
rect 9393 13231 9394 13257
rect 9366 13230 9394 13231
rect 10766 14294 10794 14322
rect 10486 14014 10514 14042
rect 10710 14014 10738 14042
rect 10598 13846 10626 13874
rect 10206 13649 10234 13650
rect 10206 13623 10207 13649
rect 10207 13623 10233 13649
rect 10233 13623 10234 13649
rect 10206 13622 10234 13623
rect 11382 18745 11410 18746
rect 11382 18719 11383 18745
rect 11383 18719 11409 18745
rect 11409 18719 11410 18745
rect 11382 18718 11410 18719
rect 12110 18718 12138 18746
rect 11158 18353 11186 18354
rect 11158 18327 11159 18353
rect 11159 18327 11185 18353
rect 11185 18327 11186 18353
rect 11158 18326 11186 18327
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 13118 18745 13146 18746
rect 13118 18719 13119 18745
rect 13119 18719 13145 18745
rect 13145 18719 13146 18745
rect 13118 18718 13146 18719
rect 12446 18326 12474 18354
rect 11102 14321 11130 14322
rect 11102 14295 11103 14321
rect 11103 14295 11129 14321
rect 11129 14295 11130 14321
rect 11102 14294 11130 14295
rect 10766 13790 10794 13818
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 10654 13174 10682 13202
rect 7798 12838 7826 12866
rect 7014 12446 7042 12474
rect 8078 12838 8106 12866
rect 7462 12222 7490 12250
rect 7350 11606 7378 11634
rect 5838 10822 5866 10850
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 2142 10401 2170 10402
rect 2142 10375 2143 10401
rect 2143 10375 2169 10401
rect 2169 10375 2170 10401
rect 2142 10374 2170 10375
rect 7406 11438 7434 11466
rect 7686 12473 7714 12474
rect 7686 12447 7687 12473
rect 7687 12447 7713 12473
rect 7713 12447 7714 12473
rect 7686 12446 7714 12447
rect 7798 12278 7826 12306
rect 7910 12222 7938 12250
rect 7854 11998 7882 12026
rect 6790 10457 6818 10458
rect 6790 10431 6791 10457
rect 6791 10431 6817 10457
rect 6817 10431 6818 10457
rect 6790 10430 6818 10431
rect 4998 10318 5026 10346
rect 966 10094 994 10122
rect 6062 10094 6090 10122
rect 4998 10038 5026 10066
rect 2142 10009 2170 10010
rect 2142 9983 2143 10009
rect 2143 9983 2169 10009
rect 2169 9983 2170 10009
rect 2142 9982 2170 9983
rect 966 9897 994 9898
rect 966 9871 967 9897
rect 967 9871 993 9897
rect 993 9871 994 9897
rect 966 9870 994 9871
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 6062 9617 6090 9618
rect 6062 9591 6063 9617
rect 6063 9591 6089 9617
rect 6089 9591 6090 9617
rect 6062 9590 6090 9591
rect 7350 10934 7378 10962
rect 7462 10849 7490 10850
rect 7462 10823 7463 10849
rect 7463 10823 7489 10849
rect 7489 10823 7490 10849
rect 7462 10822 7490 10823
rect 7126 10121 7154 10122
rect 7126 10095 7127 10121
rect 7127 10095 7153 10121
rect 7153 10095 7154 10121
rect 7126 10094 7154 10095
rect 6902 10065 6930 10066
rect 6902 10039 6903 10065
rect 6903 10039 6929 10065
rect 6929 10039 6930 10065
rect 6902 10038 6930 10039
rect 6958 9982 6986 10010
rect 7238 10038 7266 10066
rect 6902 9897 6930 9898
rect 6902 9871 6903 9897
rect 6903 9871 6929 9897
rect 6929 9871 6930 9897
rect 6902 9870 6930 9871
rect 7630 11046 7658 11074
rect 8022 11942 8050 11970
rect 8190 13145 8218 13146
rect 8190 13119 8191 13145
rect 8191 13119 8217 13145
rect 8217 13119 8218 13145
rect 8190 13118 8218 13119
rect 8358 13145 8386 13146
rect 8358 13119 8359 13145
rect 8359 13119 8385 13145
rect 8385 13119 8386 13145
rect 8358 13118 8386 13119
rect 9142 13145 9170 13146
rect 9142 13119 9143 13145
rect 9143 13119 9169 13145
rect 9169 13119 9170 13145
rect 9142 13118 9170 13119
rect 9814 13145 9842 13146
rect 9814 13119 9815 13145
rect 9815 13119 9841 13145
rect 9841 13119 9842 13145
rect 9814 13118 9842 13119
rect 9422 13089 9450 13090
rect 9422 13063 9423 13089
rect 9423 13063 9449 13089
rect 9449 13063 9450 13089
rect 9422 13062 9450 13063
rect 8414 12838 8442 12866
rect 8134 12670 8162 12698
rect 8078 11689 8106 11690
rect 8078 11663 8079 11689
rect 8079 11663 8105 11689
rect 8105 11663 8106 11689
rect 8078 11662 8106 11663
rect 7742 11633 7770 11634
rect 7742 11607 7743 11633
rect 7743 11607 7769 11633
rect 7769 11607 7770 11633
rect 7742 11606 7770 11607
rect 8190 11998 8218 12026
rect 8358 11969 8386 11970
rect 8358 11943 8359 11969
rect 8359 11943 8385 11969
rect 8385 11943 8386 11969
rect 8358 11942 8386 11943
rect 8582 12753 8610 12754
rect 8582 12727 8583 12753
rect 8583 12727 8609 12753
rect 8609 12727 8610 12753
rect 8582 12726 8610 12727
rect 10150 13145 10178 13146
rect 10150 13119 10151 13145
rect 10151 13119 10177 13145
rect 10177 13119 10178 13145
rect 10150 13118 10178 13119
rect 10822 13118 10850 13146
rect 10766 13089 10794 13090
rect 10766 13063 10767 13089
rect 10767 13063 10793 13089
rect 10793 13063 10794 13089
rect 10766 13062 10794 13063
rect 10038 12726 10066 12754
rect 8526 12697 8554 12698
rect 8526 12671 8527 12697
rect 8527 12671 8553 12697
rect 8553 12671 8554 12697
rect 8526 12670 8554 12671
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 10094 12446 10122 12474
rect 8638 11969 8666 11970
rect 8638 11943 8639 11969
rect 8639 11943 8665 11969
rect 8665 11943 8666 11969
rect 8638 11942 8666 11943
rect 8806 11662 8834 11690
rect 7686 10934 7714 10962
rect 7574 10849 7602 10850
rect 7574 10823 7575 10849
rect 7575 10823 7601 10849
rect 7601 10823 7602 10849
rect 7574 10822 7602 10823
rect 7518 10766 7546 10794
rect 7462 10598 7490 10626
rect 7406 10066 7434 10094
rect 7294 9953 7322 9954
rect 7294 9927 7295 9953
rect 7295 9927 7321 9953
rect 7321 9927 7322 9953
rect 7294 9926 7322 9927
rect 6006 9310 6034 9338
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 966 8889 994 8890
rect 966 8863 967 8889
rect 967 8863 993 8889
rect 993 8863 994 8889
rect 966 8862 994 8863
rect 4942 8889 4970 8890
rect 4942 8863 4943 8889
rect 4943 8863 4969 8889
rect 4969 8863 4970 8889
rect 4942 8862 4970 8863
rect 2142 8833 2170 8834
rect 2142 8807 2143 8833
rect 2143 8807 2169 8833
rect 2169 8807 2170 8833
rect 2142 8806 2170 8807
rect 6734 8889 6762 8890
rect 6734 8863 6735 8889
rect 6735 8863 6761 8889
rect 6761 8863 6762 8889
rect 6734 8862 6762 8863
rect 966 8414 994 8442
rect 2142 8441 2170 8442
rect 2142 8415 2143 8441
rect 2143 8415 2169 8441
rect 2169 8415 2170 8441
rect 2142 8414 2170 8415
rect 7182 9590 7210 9618
rect 7350 9870 7378 9898
rect 7854 10793 7882 10794
rect 7854 10767 7855 10793
rect 7855 10767 7881 10793
rect 7881 10767 7882 10793
rect 7854 10766 7882 10767
rect 7854 10457 7882 10458
rect 7854 10431 7855 10457
rect 7855 10431 7881 10457
rect 7881 10431 7882 10457
rect 7854 10430 7882 10431
rect 7686 10094 7714 10122
rect 7798 10318 7826 10346
rect 7182 9254 7210 9282
rect 7742 9953 7770 9954
rect 7742 9927 7743 9953
rect 7743 9927 7769 9953
rect 7769 9927 7770 9953
rect 7742 9926 7770 9927
rect 7686 9254 7714 9282
rect 7742 9646 7770 9674
rect 7910 9534 7938 9562
rect 8190 11073 8218 11074
rect 8190 11047 8191 11073
rect 8191 11047 8217 11073
rect 8217 11047 8218 11073
rect 8190 11046 8218 11047
rect 7798 9337 7826 9338
rect 7798 9311 7799 9337
rect 7799 9311 7825 9337
rect 7825 9311 7826 9337
rect 7798 9310 7826 9311
rect 7798 9225 7826 9226
rect 7798 9199 7799 9225
rect 7799 9199 7825 9225
rect 7825 9199 7826 9225
rect 7798 9198 7826 9199
rect 7126 8526 7154 8554
rect 7574 8638 7602 8666
rect 7126 8414 7154 8442
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 6734 8302 6762 8330
rect 7630 8582 7658 8610
rect 7630 8470 7658 8498
rect 7742 8470 7770 8498
rect 7630 8385 7658 8386
rect 7630 8359 7631 8385
rect 7631 8359 7657 8385
rect 7657 8359 7658 8385
rect 7630 8358 7658 8359
rect 8022 9926 8050 9954
rect 8022 9534 8050 9562
rect 8414 11465 8442 11466
rect 8414 11439 8415 11465
rect 8415 11439 8441 11465
rect 8441 11439 8442 11465
rect 8414 11438 8442 11439
rect 8582 11214 8610 11242
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 10094 11774 10122 11802
rect 11662 13398 11690 13426
rect 10822 12446 10850 12474
rect 11774 13201 11802 13202
rect 11774 13175 11775 13201
rect 11775 13175 11801 13201
rect 11801 13175 11802 13201
rect 11774 13174 11802 13175
rect 8918 11606 8946 11634
rect 8806 11158 8834 11186
rect 8414 10822 8442 10850
rect 8414 10318 8442 10346
rect 8470 11102 8498 11130
rect 8302 9590 8330 9618
rect 8414 9561 8442 9562
rect 8414 9535 8415 9561
rect 8415 9535 8441 9561
rect 8441 9535 8442 9561
rect 8414 9534 8442 9535
rect 8078 9198 8106 9226
rect 8078 8974 8106 9002
rect 7910 8694 7938 8722
rect 8134 8638 8162 8666
rect 8022 8441 8050 8442
rect 8022 8415 8023 8441
rect 8023 8415 8049 8441
rect 8049 8415 8050 8441
rect 8022 8414 8050 8415
rect 8134 8441 8162 8442
rect 8134 8415 8135 8441
rect 8135 8415 8161 8441
rect 8161 8415 8162 8441
rect 8134 8414 8162 8415
rect 6678 7630 6706 7658
rect 8134 7630 8162 7658
rect 8694 11046 8722 11074
rect 8862 11270 8890 11298
rect 8862 11129 8890 11130
rect 8862 11103 8863 11129
rect 8863 11103 8889 11129
rect 8889 11103 8890 11129
rect 8862 11102 8890 11103
rect 10654 11830 10682 11858
rect 10598 11774 10626 11802
rect 10150 11606 10178 11634
rect 8806 10318 8834 10346
rect 8750 10121 8778 10122
rect 8750 10095 8751 10121
rect 8751 10095 8777 10121
rect 8777 10095 8778 10121
rect 8750 10094 8778 10095
rect 9254 10094 9282 10122
rect 8806 9673 8834 9674
rect 8806 9647 8807 9673
rect 8807 9647 8833 9673
rect 8833 9647 8834 9673
rect 8806 9646 8834 9647
rect 8582 9198 8610 9226
rect 8694 9030 8722 9058
rect 8974 9505 9002 9506
rect 8974 9479 8975 9505
rect 8975 9479 9001 9505
rect 9001 9479 9002 9505
rect 8974 9478 9002 9479
rect 8862 8806 8890 8834
rect 8918 9366 8946 9394
rect 8246 8777 8274 8778
rect 8246 8751 8247 8777
rect 8247 8751 8273 8777
rect 8273 8751 8274 8777
rect 8246 8750 8274 8751
rect 9422 10430 9450 10458
rect 9534 10905 9562 10906
rect 9534 10879 9535 10905
rect 9535 10879 9561 10905
rect 9561 10879 9562 10905
rect 9534 10878 9562 10879
rect 9478 9982 9506 10010
rect 10094 11241 10122 11242
rect 10094 11215 10095 11241
rect 10095 11215 10121 11241
rect 10121 11215 10122 11241
rect 10094 11214 10122 11215
rect 9926 11185 9954 11186
rect 9926 11159 9927 11185
rect 9927 11159 9953 11185
rect 9953 11159 9954 11185
rect 9926 11158 9954 11159
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 10038 10401 10066 10402
rect 10038 10375 10039 10401
rect 10039 10375 10065 10401
rect 10065 10375 10066 10401
rect 10038 10374 10066 10375
rect 10094 10262 10122 10290
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9982 10121 10010 10122
rect 9982 10095 9983 10121
rect 9983 10095 10009 10121
rect 10009 10095 10010 10121
rect 9982 10094 10010 10095
rect 9926 10065 9954 10066
rect 9926 10039 9927 10065
rect 9927 10039 9953 10065
rect 9953 10039 9954 10065
rect 9926 10038 9954 10039
rect 9926 9953 9954 9954
rect 9926 9927 9927 9953
rect 9927 9927 9953 9953
rect 9953 9927 9954 9953
rect 9926 9926 9954 9927
rect 9702 9702 9730 9730
rect 9870 9617 9898 9618
rect 9870 9591 9871 9617
rect 9871 9591 9897 9617
rect 9897 9591 9898 9617
rect 9870 9590 9898 9591
rect 9478 9534 9506 9562
rect 9702 9478 9730 9506
rect 10710 11633 10738 11634
rect 10710 11607 10711 11633
rect 10711 11607 10737 11633
rect 10737 11607 10738 11633
rect 10710 11606 10738 11607
rect 10430 11577 10458 11578
rect 10430 11551 10431 11577
rect 10431 11551 10457 11577
rect 10457 11551 10458 11577
rect 10430 11550 10458 11551
rect 10766 11550 10794 11578
rect 10262 11214 10290 11242
rect 10318 11158 10346 11186
rect 10262 10934 10290 10962
rect 10262 10038 10290 10066
rect 10094 9590 10122 9618
rect 10150 9758 10178 9786
rect 9814 9366 9842 9394
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9142 9198 9170 9226
rect 9142 8918 9170 8946
rect 8918 8750 8946 8778
rect 8246 8470 8274 8498
rect 8750 8694 8778 8722
rect 8470 8526 8498 8554
rect 8806 8553 8834 8554
rect 8806 8527 8807 8553
rect 8807 8527 8833 8553
rect 8833 8527 8834 8553
rect 8806 8526 8834 8527
rect 9254 8833 9282 8834
rect 9254 8807 9255 8833
rect 9255 8807 9281 8833
rect 9281 8807 9282 8833
rect 9254 8806 9282 8807
rect 8974 8582 9002 8610
rect 10038 9254 10066 9282
rect 9982 9225 10010 9226
rect 9982 9199 9983 9225
rect 9983 9199 10009 9225
rect 10009 9199 10010 9225
rect 9982 9198 10010 9199
rect 9758 9169 9786 9170
rect 9758 9143 9759 9169
rect 9759 9143 9785 9169
rect 9785 9143 9786 9169
rect 9758 9142 9786 9143
rect 9534 8945 9562 8946
rect 9534 8919 9535 8945
rect 9535 8919 9561 8945
rect 9561 8919 9562 8945
rect 9534 8918 9562 8919
rect 10206 9366 10234 9394
rect 10654 11129 10682 11130
rect 10654 11103 10655 11129
rect 10655 11103 10681 11129
rect 10681 11103 10682 11129
rect 10654 11102 10682 11103
rect 11214 12446 11242 12474
rect 11046 12417 11074 12418
rect 11046 12391 11047 12417
rect 11047 12391 11073 12417
rect 11073 12391 11074 12417
rect 11046 12390 11074 12391
rect 11382 12473 11410 12474
rect 11382 12447 11383 12473
rect 11383 12447 11409 12473
rect 11409 12447 11410 12473
rect 11382 12446 11410 12447
rect 10878 11830 10906 11858
rect 10822 11129 10850 11130
rect 10822 11103 10823 11129
rect 10823 11103 10849 11129
rect 10849 11103 10850 11129
rect 10822 11102 10850 11103
rect 10878 10934 10906 10962
rect 10990 11185 11018 11186
rect 10990 11159 10991 11185
rect 10991 11159 11017 11185
rect 11017 11159 11018 11185
rect 10990 11158 11018 11159
rect 11326 11046 11354 11074
rect 11270 10542 11298 10570
rect 10934 10262 10962 10290
rect 11158 10206 11186 10234
rect 10654 10150 10682 10178
rect 10430 10094 10458 10122
rect 10374 10009 10402 10010
rect 10374 9983 10375 10009
rect 10375 9983 10401 10009
rect 10401 9983 10402 10009
rect 10374 9982 10402 9983
rect 10318 9646 10346 9674
rect 10150 9310 10178 9338
rect 10374 9590 10402 9618
rect 10318 9422 10346 9450
rect 10934 10009 10962 10010
rect 10934 9983 10935 10009
rect 10935 9983 10961 10009
rect 10961 9983 10962 10009
rect 10934 9982 10962 9983
rect 10878 9673 10906 9674
rect 10878 9647 10879 9673
rect 10879 9647 10905 9673
rect 10905 9647 10906 9673
rect 10878 9646 10906 9647
rect 10654 9478 10682 9506
rect 10206 9198 10234 9226
rect 10430 9225 10458 9226
rect 10430 9199 10431 9225
rect 10431 9199 10457 9225
rect 10457 9199 10458 9225
rect 10430 9198 10458 9199
rect 10262 9142 10290 9170
rect 9814 8889 9842 8890
rect 9814 8863 9815 8889
rect 9815 8863 9841 8889
rect 9841 8863 9842 8889
rect 9814 8862 9842 8863
rect 9702 8833 9730 8834
rect 9702 8807 9703 8833
rect 9703 8807 9729 8833
rect 9729 8807 9730 8833
rect 9702 8806 9730 8807
rect 9254 8470 9282 8498
rect 9422 8414 9450 8442
rect 8862 8385 8890 8386
rect 8862 8359 8863 8385
rect 8863 8359 8889 8385
rect 8889 8359 8890 8385
rect 8862 8358 8890 8359
rect 8190 7574 8218 7602
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 8190 7126 8218 7154
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 8078 2086 8106 2114
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 8414 7630 8442 7658
rect 9366 7657 9394 7658
rect 9366 7631 9367 7657
rect 9367 7631 9393 7657
rect 9393 7631 9394 7657
rect 9366 7630 9394 7631
rect 8414 7126 8442 7154
rect 8694 7574 8722 7602
rect 10206 8862 10234 8890
rect 9982 8833 10010 8834
rect 9982 8807 9983 8833
rect 9983 8807 10009 8833
rect 10009 8807 10010 8833
rect 9982 8806 10010 8807
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 9870 8497 9898 8498
rect 9870 8471 9871 8497
rect 9871 8471 9897 8497
rect 9897 8471 9898 8497
rect 9870 8470 9898 8471
rect 10374 8833 10402 8834
rect 10374 8807 10375 8833
rect 10375 8807 10401 8833
rect 10401 8807 10402 8833
rect 10374 8806 10402 8807
rect 9982 8049 10010 8050
rect 9982 8023 9983 8049
rect 9983 8023 10009 8049
rect 10009 8023 10010 8049
rect 9982 8022 10010 8023
rect 9814 7910 9842 7938
rect 8918 7126 8946 7154
rect 9478 7126 9506 7154
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 10710 9337 10738 9338
rect 10710 9311 10711 9337
rect 10711 9311 10737 9337
rect 10737 9311 10738 9337
rect 10710 9310 10738 9311
rect 10990 9478 11018 9506
rect 11326 10065 11354 10066
rect 11326 10039 11327 10065
rect 11327 10039 11353 10065
rect 11353 10039 11354 10065
rect 11326 10038 11354 10039
rect 11102 9758 11130 9786
rect 11046 9422 11074 9450
rect 10934 9254 10962 9282
rect 10822 9142 10850 9170
rect 10990 9030 11018 9058
rect 12558 13454 12586 13482
rect 12278 13174 12306 13202
rect 12110 12390 12138 12418
rect 12334 11857 12362 11858
rect 12334 11831 12335 11857
rect 12335 11831 12361 11857
rect 12361 11831 12362 11857
rect 12334 11830 12362 11831
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 13062 18353 13090 18354
rect 13062 18327 13063 18353
rect 13063 18327 13089 18353
rect 13089 18327 13090 18353
rect 13062 18326 13090 18327
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 20118 17150 20146 17178
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 13118 13537 13146 13538
rect 13118 13511 13119 13537
rect 13119 13511 13145 13537
rect 13145 13511 13146 13537
rect 13118 13510 13146 13511
rect 13454 13510 13482 13538
rect 13622 13510 13650 13538
rect 12950 13481 12978 13482
rect 12950 13455 12951 13481
rect 12951 13455 12977 13481
rect 12977 13455 12978 13481
rect 12950 13454 12978 13455
rect 13062 13481 13090 13482
rect 13062 13455 13063 13481
rect 13063 13455 13089 13481
rect 13089 13455 13090 13481
rect 13062 13454 13090 13455
rect 12670 13145 12698 13146
rect 12670 13119 12671 13145
rect 12671 13119 12697 13145
rect 12697 13119 12698 13145
rect 12670 13118 12698 13119
rect 12670 12641 12698 12642
rect 12670 12615 12671 12641
rect 12671 12615 12697 12641
rect 12697 12615 12698 12641
rect 12670 12614 12698 12615
rect 13006 12614 13034 12642
rect 14406 13510 14434 13538
rect 14070 13454 14098 13482
rect 14294 13145 14322 13146
rect 14294 13119 14295 13145
rect 14295 13119 14321 13145
rect 14321 13119 14322 13145
rect 14294 13118 14322 13119
rect 14070 13006 14098 13034
rect 18830 13537 18858 13538
rect 18830 13511 18831 13537
rect 18831 13511 18857 13537
rect 18857 13511 18858 13537
rect 18830 13510 18858 13511
rect 14630 13118 14658 13146
rect 18830 13145 18858 13146
rect 18830 13119 18831 13145
rect 18831 13119 18857 13145
rect 18857 13119 18858 13145
rect 18830 13118 18858 13119
rect 20006 13118 20034 13146
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 20006 12782 20034 12810
rect 13342 12446 13370 12474
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 11662 11774 11690 11802
rect 11886 11774 11914 11802
rect 11550 10401 11578 10402
rect 11550 10375 11551 10401
rect 11551 10375 11577 10401
rect 11577 10375 11578 10401
rect 11550 10374 11578 10375
rect 11438 10289 11466 10290
rect 11438 10263 11439 10289
rect 11439 10263 11465 10289
rect 11465 10263 11466 10289
rect 11438 10262 11466 10263
rect 11214 9590 11242 9618
rect 11214 9310 11242 9338
rect 11270 9534 11298 9562
rect 11102 9198 11130 9226
rect 10766 8889 10794 8890
rect 10766 8863 10767 8889
rect 10767 8863 10793 8889
rect 10793 8863 10794 8889
rect 10766 8862 10794 8863
rect 10822 8833 10850 8834
rect 10822 8807 10823 8833
rect 10823 8807 10849 8833
rect 10849 8807 10850 8833
rect 10822 8806 10850 8807
rect 11158 9142 11186 9170
rect 11494 9702 11522 9730
rect 11606 9534 11634 9562
rect 11606 9337 11634 9338
rect 11606 9311 11607 9337
rect 11607 9311 11633 9337
rect 11633 9311 11634 9337
rect 11606 9310 11634 9311
rect 11326 8974 11354 9002
rect 10654 8049 10682 8050
rect 10654 8023 10655 8049
rect 10655 8023 10681 8049
rect 10681 8023 10682 8049
rect 10654 8022 10682 8023
rect 10710 7910 10738 7938
rect 10206 7630 10234 7658
rect 10374 7153 10402 7154
rect 10374 7127 10375 7153
rect 10375 7127 10401 7153
rect 10401 7127 10402 7153
rect 10374 7126 10402 7127
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 12110 11774 12138 11802
rect 11886 11270 11914 11298
rect 11942 10878 11970 10906
rect 11886 10318 11914 10346
rect 11886 10150 11914 10178
rect 11718 9169 11746 9170
rect 11718 9143 11719 9169
rect 11719 9143 11745 9169
rect 11745 9143 11746 9169
rect 11718 9142 11746 9143
rect 11382 8862 11410 8890
rect 11718 8862 11746 8890
rect 11550 8833 11578 8834
rect 11550 8807 11551 8833
rect 11551 8807 11577 8833
rect 11577 8807 11578 8833
rect 11550 8806 11578 8807
rect 11886 8526 11914 8554
rect 12054 11102 12082 11130
rect 11998 10206 12026 10234
rect 12390 11129 12418 11130
rect 12390 11103 12391 11129
rect 12391 11103 12417 11129
rect 12417 11103 12418 11129
rect 12390 11102 12418 11103
rect 12166 10822 12194 10850
rect 12222 10766 12250 10794
rect 12166 10598 12194 10626
rect 12558 10710 12586 10738
rect 12334 10262 12362 10290
rect 12278 10150 12306 10178
rect 12110 9617 12138 9618
rect 12110 9591 12111 9617
rect 12111 9591 12137 9617
rect 12137 9591 12138 9617
rect 12110 9590 12138 9591
rect 12894 11830 12922 11858
rect 12894 11550 12922 11578
rect 13286 11577 13314 11578
rect 13286 11551 13287 11577
rect 13287 11551 13313 11577
rect 13313 11551 13314 11577
rect 13286 11550 13314 11551
rect 12670 10905 12698 10906
rect 12670 10879 12671 10905
rect 12671 10879 12697 10905
rect 12697 10879 12698 10905
rect 12670 10878 12698 10879
rect 12726 10793 12754 10794
rect 12726 10767 12727 10793
rect 12727 10767 12753 10793
rect 12753 10767 12754 10793
rect 12726 10766 12754 10767
rect 12614 10542 12642 10570
rect 13342 10934 13370 10962
rect 13118 10849 13146 10850
rect 13118 10823 13119 10849
rect 13119 10823 13145 10849
rect 13145 10823 13146 10849
rect 13118 10822 13146 10823
rect 12782 10094 12810 10122
rect 12838 10065 12866 10066
rect 12838 10039 12839 10065
rect 12839 10039 12865 10065
rect 12865 10039 12866 10065
rect 12838 10038 12866 10039
rect 12222 9702 12250 9730
rect 12390 9617 12418 9618
rect 12390 9591 12391 9617
rect 12391 9591 12417 9617
rect 12417 9591 12418 9617
rect 12390 9590 12418 9591
rect 12614 9617 12642 9618
rect 12614 9591 12615 9617
rect 12615 9591 12641 9617
rect 12641 9591 12642 9617
rect 12614 9590 12642 9591
rect 12894 9590 12922 9618
rect 12166 9310 12194 9338
rect 13006 9310 13034 9338
rect 14910 11550 14938 11578
rect 13622 11270 13650 11298
rect 14742 11521 14770 11522
rect 14742 11495 14743 11521
rect 14743 11495 14769 11521
rect 14769 11495 14770 11521
rect 14742 11494 14770 11495
rect 13566 10934 13594 10962
rect 14014 11214 14042 11242
rect 14294 11241 14322 11242
rect 14294 11215 14295 11241
rect 14295 11215 14321 11241
rect 14321 11215 14322 11241
rect 14294 11214 14322 11215
rect 14070 10793 14098 10794
rect 14070 10767 14071 10793
rect 14071 10767 14097 10793
rect 14097 10767 14098 10793
rect 14070 10766 14098 10767
rect 14686 11270 14714 11298
rect 18830 11577 18858 11578
rect 18830 11551 18831 11577
rect 18831 11551 18857 11577
rect 18857 11551 18858 11577
rect 18830 11550 18858 11551
rect 20006 11465 20034 11466
rect 20006 11439 20007 11465
rect 20007 11439 20033 11465
rect 20033 11439 20034 11465
rect 20006 11438 20034 11439
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 18830 11185 18858 11186
rect 18830 11159 18831 11185
rect 18831 11159 18857 11185
rect 18857 11159 18858 11185
rect 18830 11158 18858 11159
rect 20006 11102 20034 11130
rect 14574 10766 14602 10794
rect 13286 10430 13314 10458
rect 13230 10038 13258 10066
rect 13174 9505 13202 9506
rect 13174 9479 13175 9505
rect 13175 9479 13201 9505
rect 13201 9479 13202 9505
rect 13174 9478 13202 9479
rect 13118 9310 13146 9338
rect 12054 8833 12082 8834
rect 12054 8807 12055 8833
rect 12055 8807 12081 8833
rect 12081 8807 12082 8833
rect 12054 8806 12082 8807
rect 12222 8470 12250 8498
rect 11270 8022 11298 8050
rect 11774 8049 11802 8050
rect 11774 8023 11775 8049
rect 11775 8023 11801 8049
rect 11801 8023 11802 8049
rect 11774 8022 11802 8023
rect 12894 8049 12922 8050
rect 12894 8023 12895 8049
rect 12895 8023 12921 8049
rect 12921 8023 12922 8049
rect 12894 8022 12922 8023
rect 12054 7993 12082 7994
rect 12054 7967 12055 7993
rect 12055 7967 12081 7993
rect 12081 7967 12082 7993
rect 12054 7966 12082 7967
rect 12614 7966 12642 7994
rect 13286 9366 13314 9394
rect 13230 9198 13258 9226
rect 13678 9505 13706 9506
rect 13678 9479 13679 9505
rect 13679 9479 13705 9505
rect 13705 9479 13706 9505
rect 13678 9478 13706 9479
rect 13454 9254 13482 9282
rect 13286 9030 13314 9058
rect 13734 9254 13762 9282
rect 13510 9142 13538 9170
rect 13174 8526 13202 8554
rect 13230 8694 13258 8722
rect 13902 9617 13930 9618
rect 13902 9591 13903 9617
rect 13903 9591 13929 9617
rect 13929 9591 13930 9617
rect 13902 9590 13930 9591
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 18830 10009 18858 10010
rect 18830 9983 18831 10009
rect 18831 9983 18857 10009
rect 18857 9983 18858 10009
rect 18830 9982 18858 9983
rect 14630 9926 14658 9954
rect 15246 9953 15274 9954
rect 15246 9927 15247 9953
rect 15247 9927 15273 9953
rect 15273 9927 15274 9953
rect 15246 9926 15274 9927
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 20006 9758 20034 9786
rect 14742 9617 14770 9618
rect 14742 9591 14743 9617
rect 14743 9591 14769 9617
rect 14769 9591 14770 9617
rect 14742 9590 14770 9591
rect 13846 9310 13874 9338
rect 14014 9366 14042 9394
rect 13790 9030 13818 9058
rect 14126 9225 14154 9226
rect 14126 9199 14127 9225
rect 14127 9199 14153 9225
rect 14153 9199 14154 9225
rect 14126 9198 14154 9199
rect 18830 9225 18858 9226
rect 18830 9199 18831 9225
rect 18831 9199 18857 9225
rect 18857 9199 18858 9225
rect 18830 9198 18858 9199
rect 15190 9169 15218 9170
rect 15190 9143 15191 9169
rect 15191 9143 15217 9169
rect 15217 9143 15218 9169
rect 15190 9142 15218 9143
rect 13958 8806 13986 8834
rect 13734 8721 13762 8722
rect 13734 8695 13735 8721
rect 13735 8695 13761 8721
rect 13761 8695 13762 8721
rect 13734 8694 13762 8695
rect 13454 8553 13482 8554
rect 13454 8527 13455 8553
rect 13455 8527 13481 8553
rect 13481 8527 13482 8553
rect 13454 8526 13482 8527
rect 14294 8806 14322 8834
rect 13622 8497 13650 8498
rect 13622 8471 13623 8497
rect 13623 8471 13649 8497
rect 13649 8471 13650 8497
rect 13622 8470 13650 8471
rect 14070 8777 14098 8778
rect 14070 8751 14071 8777
rect 14071 8751 14097 8777
rect 14097 8751 14098 8777
rect 14070 8750 14098 8751
rect 14014 8497 14042 8498
rect 14014 8471 14015 8497
rect 14015 8471 14041 8497
rect 14041 8471 14042 8497
rect 14014 8470 14042 8471
rect 13566 8414 13594 8442
rect 20006 9113 20034 9114
rect 20006 9087 20007 9113
rect 20007 9087 20033 9113
rect 20033 9087 20034 9113
rect 20006 9086 20034 9087
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 15190 8750 15218 8778
rect 14518 8414 14546 8442
rect 13398 8022 13426 8050
rect 18830 8441 18858 8442
rect 18830 8415 18831 8441
rect 18831 8415 18857 8441
rect 18857 8415 18858 8441
rect 18830 8414 18858 8415
rect 20006 8414 20034 8442
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 19950 8078 19978 8106
rect 14630 8049 14658 8050
rect 14630 8023 14631 8049
rect 14631 8023 14657 8049
rect 14657 8023 14658 8049
rect 14630 8022 14658 8023
rect 14854 8022 14882 8050
rect 14630 7713 14658 7714
rect 14630 7687 14631 7713
rect 14631 7687 14657 7713
rect 14657 7687 14658 7713
rect 14630 7686 14658 7687
rect 20006 7742 20034 7770
rect 18830 7686 18858 7714
rect 11382 7265 11410 7266
rect 11382 7239 11383 7265
rect 11383 7239 11409 7265
rect 11409 7239 11410 7265
rect 11382 7238 11410 7239
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 12894 7238 12922 7266
rect 13062 7265 13090 7266
rect 13062 7239 13063 7265
rect 13063 7239 13089 7265
rect 13089 7239 13090 7265
rect 13062 7238 13090 7239
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9254 2113 9282 2114
rect 9254 2087 9255 2113
rect 9255 2087 9281 2113
rect 9281 2087 9282 2113
rect 9254 2086 9282 2087
rect 12446 1806 12474 1834
rect 8582 1694 8610 1722
rect 9030 1694 9058 1722
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 13062 1833 13090 1834
rect 13062 1807 13063 1833
rect 13063 1807 13089 1833
rect 13089 1807 13090 1833
rect 13062 1806 13090 1807
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 8745 19110 8750 19138
rect 8778 19110 9310 19138
rect 9338 19110 9343 19138
rect 11769 19110 11774 19138
rect 11802 19110 12782 19138
rect 12810 19110 12815 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 10761 18718 10766 18746
rect 10794 18718 11382 18746
rect 11410 18718 11415 18746
rect 12105 18718 12110 18746
rect 12138 18718 13118 18746
rect 13146 18718 13151 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 8073 18326 8078 18354
rect 8106 18326 8694 18354
rect 8722 18326 8727 18354
rect 10425 18326 10430 18354
rect 10458 18326 11158 18354
rect 11186 18326 11191 18354
rect 12441 18326 12446 18354
rect 12474 18326 13062 18354
rect 13090 18326 13095 18354
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 20600 17178 21000 17192
rect 20113 17150 20118 17178
rect 20146 17150 21000 17178
rect 20600 17136 21000 17150
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 10761 14294 10766 14322
rect 10794 14294 11102 14322
rect 11130 14294 11135 14322
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 10033 14014 10038 14042
rect 10066 14014 10486 14042
rect 10514 14014 10710 14042
rect 10738 14014 10743 14042
rect 8801 13846 8806 13874
rect 8834 13846 9310 13874
rect 9338 13846 10598 13874
rect 10626 13846 10631 13874
rect 0 13818 400 13832
rect 0 13790 5782 13818
rect 5810 13790 5815 13818
rect 9809 13790 9814 13818
rect 9842 13790 10766 13818
rect 10794 13790 10799 13818
rect 0 13776 400 13790
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 9641 13622 9646 13650
rect 9674 13622 10206 13650
rect 10234 13622 10239 13650
rect 6729 13566 6734 13594
rect 6762 13566 7014 13594
rect 7042 13566 8414 13594
rect 8442 13566 8638 13594
rect 8666 13566 8806 13594
rect 8834 13566 8839 13594
rect 11662 13510 13118 13538
rect 13146 13510 13454 13538
rect 13482 13510 13487 13538
rect 13617 13510 13622 13538
rect 13650 13510 14406 13538
rect 14434 13510 18830 13538
rect 18858 13510 18863 13538
rect 11662 13426 11690 13510
rect 12553 13454 12558 13482
rect 12586 13454 12950 13482
rect 12978 13454 12983 13482
rect 13057 13454 13062 13482
rect 13090 13454 14070 13482
rect 14098 13454 14103 13482
rect 8801 13398 8806 13426
rect 8834 13398 9030 13426
rect 9058 13398 11662 13426
rect 11690 13398 11695 13426
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 8969 13230 8974 13258
rect 9002 13230 9366 13258
rect 9394 13230 9399 13258
rect 7849 13174 7854 13202
rect 7882 13174 8638 13202
rect 8666 13174 8671 13202
rect 9814 13174 10654 13202
rect 10682 13174 10687 13202
rect 11769 13174 11774 13202
rect 11802 13174 12278 13202
rect 12306 13174 12311 13202
rect 9814 13146 9842 13174
rect 20600 13146 21000 13160
rect 7569 13118 7574 13146
rect 7602 13118 8190 13146
rect 8218 13118 8223 13146
rect 8353 13118 8358 13146
rect 8386 13118 9142 13146
rect 9170 13118 9814 13146
rect 9842 13118 9847 13146
rect 10145 13118 10150 13146
rect 10178 13118 10822 13146
rect 10850 13118 10855 13146
rect 12665 13118 12670 13146
rect 12698 13118 14294 13146
rect 14322 13118 14630 13146
rect 14658 13118 14663 13146
rect 15946 13118 18830 13146
rect 18858 13118 18863 13146
rect 20001 13118 20006 13146
rect 20034 13118 21000 13146
rect 9417 13062 9422 13090
rect 9450 13062 10766 13090
rect 10794 13062 10799 13090
rect 15946 13034 15974 13118
rect 20600 13104 21000 13118
rect 14065 13006 14070 13034
rect 14098 13006 15974 13034
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 7793 12838 7798 12866
rect 7826 12838 8078 12866
rect 8106 12838 8414 12866
rect 8442 12838 8447 12866
rect 20600 12810 21000 12824
rect 20001 12782 20006 12810
rect 20034 12782 21000 12810
rect 20600 12768 21000 12782
rect 8577 12726 8582 12754
rect 8610 12726 10038 12754
rect 10066 12726 10071 12754
rect 8129 12670 8134 12698
rect 8162 12670 8526 12698
rect 8554 12670 8559 12698
rect 12665 12614 12670 12642
rect 12698 12614 13006 12642
rect 13034 12614 13039 12642
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 6169 12446 6174 12474
rect 6202 12446 6846 12474
rect 6874 12446 7014 12474
rect 7042 12446 7686 12474
rect 7714 12446 7719 12474
rect 10089 12446 10094 12474
rect 10122 12446 10822 12474
rect 10850 12446 11214 12474
rect 11242 12446 11247 12474
rect 11377 12446 11382 12474
rect 11410 12446 13342 12474
rect 13370 12446 13375 12474
rect 11041 12390 11046 12418
rect 11074 12390 12110 12418
rect 12138 12390 12143 12418
rect 6393 12278 6398 12306
rect 6426 12278 7798 12306
rect 7826 12278 7831 12306
rect 7457 12222 7462 12250
rect 7490 12222 7910 12250
rect 7938 12222 7943 12250
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 7849 11998 7854 12026
rect 7882 11998 8190 12026
rect 8218 11998 8223 12026
rect 8017 11942 8022 11970
rect 8050 11942 8358 11970
rect 8386 11942 8638 11970
rect 8666 11942 8671 11970
rect 10649 11830 10654 11858
rect 10682 11830 10878 11858
rect 10906 11830 12334 11858
rect 12362 11830 12894 11858
rect 12922 11830 12927 11858
rect 10089 11774 10094 11802
rect 10122 11774 10598 11802
rect 10626 11774 10631 11802
rect 11657 11774 11662 11802
rect 11690 11774 11886 11802
rect 11914 11774 12110 11802
rect 12138 11774 12143 11802
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 5497 11718 5502 11746
rect 5530 11718 6062 11746
rect 6090 11718 6095 11746
rect 7546 11662 8078 11690
rect 8106 11662 8806 11690
rect 8834 11662 8839 11690
rect 7546 11634 7574 11662
rect 7345 11606 7350 11634
rect 7378 11606 7574 11634
rect 7737 11606 7742 11634
rect 7770 11606 8918 11634
rect 8946 11606 8951 11634
rect 10145 11606 10150 11634
rect 10178 11606 10710 11634
rect 10738 11606 10743 11634
rect 10425 11550 10430 11578
rect 10458 11550 10766 11578
rect 10794 11550 10799 11578
rect 12889 11550 12894 11578
rect 12922 11550 13286 11578
rect 13314 11550 14910 11578
rect 14938 11550 14943 11578
rect 15946 11550 18830 11578
rect 18858 11550 18863 11578
rect 15946 11522 15974 11550
rect 14737 11494 14742 11522
rect 14770 11494 15974 11522
rect 20600 11466 21000 11480
rect 7401 11438 7406 11466
rect 7434 11438 8414 11466
rect 8442 11438 8447 11466
rect 20001 11438 20006 11466
rect 20034 11438 21000 11466
rect 20600 11424 21000 11438
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 8857 11270 8862 11298
rect 8890 11270 11886 11298
rect 11914 11270 11919 11298
rect 13617 11270 13622 11298
rect 13650 11270 14686 11298
rect 14714 11270 14719 11298
rect 8577 11214 8582 11242
rect 8610 11214 10094 11242
rect 10122 11214 10262 11242
rect 10290 11214 10295 11242
rect 14009 11214 14014 11242
rect 14042 11214 14294 11242
rect 14322 11214 15974 11242
rect 15946 11186 15974 11214
rect 8801 11158 8806 11186
rect 8834 11158 9926 11186
rect 9954 11158 9959 11186
rect 10313 11158 10318 11186
rect 10346 11158 10990 11186
rect 11018 11158 11023 11186
rect 15946 11158 18830 11186
rect 18858 11158 18863 11186
rect 9926 11130 9954 11158
rect 20600 11130 21000 11144
rect 8465 11102 8470 11130
rect 8498 11102 8862 11130
rect 8890 11102 8895 11130
rect 9926 11102 10654 11130
rect 10682 11102 10687 11130
rect 10817 11102 10822 11130
rect 10850 11102 12054 11130
rect 12082 11102 12390 11130
rect 12418 11102 12423 11130
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 20600 11088 21000 11102
rect 7625 11046 7630 11074
rect 7658 11046 8190 11074
rect 8218 11046 8694 11074
rect 8722 11046 11326 11074
rect 11354 11046 11359 11074
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 7345 10934 7350 10962
rect 7378 10934 7686 10962
rect 7714 10934 7719 10962
rect 10257 10934 10262 10962
rect 10290 10934 10878 10962
rect 10906 10934 10911 10962
rect 13337 10934 13342 10962
rect 13370 10934 13566 10962
rect 13594 10934 13599 10962
rect 5777 10878 5782 10906
rect 5810 10878 9534 10906
rect 9562 10878 9567 10906
rect 11937 10878 11942 10906
rect 11970 10878 12670 10906
rect 12698 10878 12703 10906
rect 5833 10822 5838 10850
rect 5866 10822 7462 10850
rect 7490 10822 7495 10850
rect 7569 10822 7574 10850
rect 7602 10822 8414 10850
rect 8442 10822 8447 10850
rect 12161 10822 12166 10850
rect 12194 10822 13118 10850
rect 13146 10822 13151 10850
rect 7513 10766 7518 10794
rect 7546 10766 7854 10794
rect 7882 10766 7887 10794
rect 12217 10766 12222 10794
rect 12250 10766 12726 10794
rect 12754 10766 12759 10794
rect 13426 10766 14070 10794
rect 14098 10766 14574 10794
rect 14602 10766 14607 10794
rect 13426 10738 13454 10766
rect 12553 10710 12558 10738
rect 12586 10710 13454 10738
rect 7457 10598 7462 10626
rect 7490 10598 12166 10626
rect 12194 10598 12199 10626
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 11265 10542 11270 10570
rect 11298 10542 12614 10570
rect 12642 10542 12647 10570
rect 6785 10430 6790 10458
rect 6818 10430 7854 10458
rect 7882 10430 7887 10458
rect 9417 10430 9422 10458
rect 9450 10430 13286 10458
rect 13314 10430 13319 10458
rect 2137 10374 2142 10402
rect 2170 10374 4214 10402
rect 10033 10374 10038 10402
rect 10066 10374 11550 10402
rect 11578 10374 11583 10402
rect 4186 10346 4214 10374
rect 4186 10318 4998 10346
rect 5026 10318 7798 10346
rect 7826 10318 7831 10346
rect 8409 10318 8414 10346
rect 8442 10318 8806 10346
rect 8834 10318 11886 10346
rect 11914 10318 11919 10346
rect 10089 10262 10094 10290
rect 10122 10262 10934 10290
rect 10962 10262 10967 10290
rect 11433 10262 11438 10290
rect 11466 10262 12334 10290
rect 12362 10262 12367 10290
rect 10094 10206 11158 10234
rect 11186 10206 11998 10234
rect 12026 10206 12031 10234
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 0 10122 400 10136
rect 10094 10122 10122 10206
rect 0 10094 966 10122
rect 994 10094 999 10122
rect 6057 10094 6062 10122
rect 6090 10094 7126 10122
rect 7154 10094 7159 10122
rect 7681 10094 7686 10122
rect 7714 10094 8750 10122
rect 8778 10094 8783 10122
rect 9249 10094 9254 10122
rect 9282 10094 9982 10122
rect 10010 10094 10122 10122
rect 10150 10150 10654 10178
rect 10682 10150 10687 10178
rect 11881 10150 11886 10178
rect 11914 10150 12278 10178
rect 12306 10150 12311 10178
rect 0 10080 400 10094
rect 7401 10066 7406 10094
rect 7434 10066 7439 10094
rect 10150 10066 10178 10150
rect 10425 10094 10430 10122
rect 10458 10094 12782 10122
rect 12810 10094 12815 10122
rect 4186 10038 4998 10066
rect 5026 10038 6902 10066
rect 6930 10038 6935 10066
rect 7233 10038 7238 10066
rect 7266 10038 7434 10066
rect 9921 10038 9926 10066
rect 9954 10038 10178 10066
rect 10257 10038 10262 10066
rect 10290 10038 11326 10066
rect 11354 10038 11359 10066
rect 12833 10038 12838 10066
rect 12866 10038 13230 10066
rect 13258 10038 13263 10066
rect 4186 10010 4214 10038
rect 2137 9982 2142 10010
rect 2170 9982 4214 10010
rect 6953 9982 6958 10010
rect 6986 9982 9478 10010
rect 9506 9982 9511 10010
rect 10369 9982 10374 10010
rect 10402 9982 10934 10010
rect 10962 9982 10967 10010
rect 15946 9982 18830 10010
rect 18858 9982 18863 10010
rect 15946 9954 15974 9982
rect 7289 9926 7294 9954
rect 7322 9926 7742 9954
rect 7770 9926 7775 9954
rect 8017 9926 8022 9954
rect 8050 9926 9926 9954
rect 9954 9926 9959 9954
rect 14625 9926 14630 9954
rect 14658 9926 15246 9954
rect 15274 9926 15974 9954
rect 961 9870 966 9898
rect 994 9870 999 9898
rect 6897 9870 6902 9898
rect 6930 9870 7350 9898
rect 7378 9870 7383 9898
rect 0 9786 400 9800
rect 966 9786 994 9870
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 20600 9786 21000 9800
rect 0 9758 994 9786
rect 10145 9758 10150 9786
rect 10178 9758 11102 9786
rect 11130 9758 11135 9786
rect 20001 9758 20006 9786
rect 20034 9758 21000 9786
rect 0 9744 400 9758
rect 20600 9744 21000 9758
rect 9697 9702 9702 9730
rect 9730 9702 11494 9730
rect 11522 9702 12222 9730
rect 12250 9702 12255 9730
rect 7737 9646 7742 9674
rect 7770 9646 8806 9674
rect 8834 9646 8839 9674
rect 9870 9646 10150 9674
rect 10178 9646 10183 9674
rect 10313 9646 10318 9674
rect 10346 9646 10878 9674
rect 10906 9646 10911 9674
rect 9870 9618 9898 9646
rect 6057 9590 6062 9618
rect 6090 9590 7182 9618
rect 7210 9590 7215 9618
rect 8297 9590 8302 9618
rect 8330 9590 9870 9618
rect 9898 9590 9903 9618
rect 10089 9590 10094 9618
rect 10122 9590 10374 9618
rect 10402 9590 10407 9618
rect 11209 9590 11214 9618
rect 11242 9590 12110 9618
rect 12138 9590 12143 9618
rect 12385 9590 12390 9618
rect 12418 9590 12614 9618
rect 12642 9590 12894 9618
rect 12922 9590 12927 9618
rect 13897 9590 13902 9618
rect 13930 9590 14742 9618
rect 14770 9590 14775 9618
rect 7905 9534 7910 9562
rect 7938 9534 8022 9562
rect 8050 9534 8414 9562
rect 8442 9534 8447 9562
rect 9473 9534 9478 9562
rect 9506 9534 11270 9562
rect 11298 9534 11606 9562
rect 11634 9534 11639 9562
rect 8969 9478 8974 9506
rect 9002 9478 9702 9506
rect 9730 9478 10654 9506
rect 10682 9478 10687 9506
rect 10985 9478 10990 9506
rect 11018 9478 13174 9506
rect 13202 9478 13678 9506
rect 13706 9478 13711 9506
rect 10145 9422 10150 9450
rect 10178 9422 10318 9450
rect 10346 9422 11046 9450
rect 11074 9422 11079 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 8913 9366 8918 9394
rect 8946 9366 9814 9394
rect 9842 9366 9847 9394
rect 10089 9366 10094 9394
rect 10122 9366 10206 9394
rect 10234 9366 10239 9394
rect 13281 9366 13286 9394
rect 13314 9366 14014 9394
rect 14042 9366 14047 9394
rect 6001 9310 6006 9338
rect 6034 9310 7798 9338
rect 7826 9310 7831 9338
rect 10131 9310 10150 9338
rect 10178 9310 10183 9338
rect 10705 9310 10710 9338
rect 10738 9310 11214 9338
rect 11242 9310 11247 9338
rect 11601 9310 11606 9338
rect 11634 9310 11639 9338
rect 12161 9310 12166 9338
rect 12194 9310 13006 9338
rect 13034 9310 13039 9338
rect 13113 9310 13118 9338
rect 13146 9310 13846 9338
rect 13874 9310 13879 9338
rect 11606 9282 11634 9310
rect 13734 9282 13762 9310
rect 7177 9254 7182 9282
rect 7210 9254 7686 9282
rect 7714 9254 7719 9282
rect 10033 9254 10038 9282
rect 10066 9254 10934 9282
rect 10962 9254 10967 9282
rect 11606 9254 13454 9282
rect 13482 9254 13487 9282
rect 13729 9254 13734 9282
rect 13762 9254 13767 9282
rect 7793 9198 7798 9226
rect 7826 9198 8078 9226
rect 8106 9198 8111 9226
rect 8577 9198 8582 9226
rect 8610 9198 9142 9226
rect 9170 9198 9175 9226
rect 9977 9198 9982 9226
rect 10010 9198 10094 9226
rect 10122 9198 10127 9226
rect 10201 9198 10206 9226
rect 10234 9198 10430 9226
rect 10458 9198 11102 9226
rect 11130 9198 11135 9226
rect 13225 9198 13230 9226
rect 13258 9198 14126 9226
rect 14154 9198 14159 9226
rect 15946 9198 18830 9226
rect 18858 9198 18863 9226
rect 15946 9170 15974 9198
rect 9753 9142 9758 9170
rect 9786 9142 9791 9170
rect 10257 9142 10262 9170
rect 10290 9142 10822 9170
rect 10850 9142 10855 9170
rect 11153 9142 11158 9170
rect 11186 9142 11718 9170
rect 11746 9142 11751 9170
rect 13505 9142 13510 9170
rect 13538 9142 13543 9170
rect 15185 9142 15190 9170
rect 15218 9142 15974 9170
rect 9758 9114 9786 9142
rect 13510 9114 13538 9142
rect 20600 9114 21000 9128
rect 9758 9086 13538 9114
rect 20001 9086 20006 9114
rect 20034 9086 21000 9114
rect 20600 9072 21000 9086
rect 8689 9030 8694 9058
rect 8722 9030 10990 9058
rect 11018 9030 11023 9058
rect 13281 9030 13286 9058
rect 13314 9030 13790 9058
rect 13818 9030 13823 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 8073 8974 8078 9002
rect 8106 8974 11326 9002
rect 11354 8974 11359 9002
rect 9137 8918 9142 8946
rect 9170 8918 9534 8946
rect 9562 8918 9567 8946
rect 961 8862 966 8890
rect 994 8862 999 8890
rect 4186 8862 4942 8890
rect 4970 8862 6734 8890
rect 6762 8862 6767 8890
rect 9809 8862 9814 8890
rect 9842 8862 10206 8890
rect 10234 8862 10239 8890
rect 10761 8862 10766 8890
rect 10794 8862 11382 8890
rect 11410 8862 11718 8890
rect 11746 8862 11751 8890
rect 0 8778 400 8792
rect 966 8778 994 8862
rect 4186 8834 4214 8862
rect 2137 8806 2142 8834
rect 2170 8806 4214 8834
rect 8857 8806 8862 8834
rect 8890 8806 9254 8834
rect 9282 8806 9287 8834
rect 9697 8806 9702 8834
rect 9730 8806 9982 8834
rect 10010 8806 10015 8834
rect 10369 8806 10374 8834
rect 10402 8806 10822 8834
rect 10850 8806 10855 8834
rect 11545 8806 11550 8834
rect 11578 8806 12054 8834
rect 12082 8806 12087 8834
rect 13953 8806 13958 8834
rect 13986 8806 14294 8834
rect 14322 8806 18830 8834
rect 18858 8806 18863 8834
rect 0 8750 994 8778
rect 8241 8750 8246 8778
rect 8274 8750 8918 8778
rect 8946 8750 8951 8778
rect 14065 8750 14070 8778
rect 14098 8750 15190 8778
rect 15218 8750 15223 8778
rect 0 8736 400 8750
rect 7905 8694 7910 8722
rect 7938 8694 8750 8722
rect 8778 8694 8783 8722
rect 13225 8694 13230 8722
rect 13258 8694 13734 8722
rect 13762 8694 13767 8722
rect 7569 8638 7574 8666
rect 7602 8638 8134 8666
rect 8162 8638 8167 8666
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 7625 8582 7630 8610
rect 7658 8582 8974 8610
rect 9002 8582 9007 8610
rect 7121 8526 7126 8554
rect 7154 8526 7770 8554
rect 8465 8526 8470 8554
rect 8498 8526 8806 8554
rect 8834 8526 11886 8554
rect 11914 8526 11919 8554
rect 13169 8526 13174 8554
rect 13202 8526 13454 8554
rect 13482 8526 13487 8554
rect 7742 8498 7770 8526
rect 6734 8470 7630 8498
rect 7658 8470 7663 8498
rect 7737 8470 7742 8498
rect 7770 8470 8246 8498
rect 8274 8470 8279 8498
rect 9249 8470 9254 8498
rect 9282 8470 9870 8498
rect 9898 8470 10150 8498
rect 10178 8470 10183 8498
rect 12217 8470 12222 8498
rect 12250 8470 13622 8498
rect 13650 8470 14014 8498
rect 14042 8470 14047 8498
rect 0 8442 400 8456
rect 6734 8442 6762 8470
rect 20600 8442 21000 8456
rect 0 8414 966 8442
rect 994 8414 999 8442
rect 2137 8414 2142 8442
rect 2170 8414 6762 8442
rect 7121 8414 7126 8442
rect 7154 8414 8022 8442
rect 8050 8414 8055 8442
rect 8129 8414 8134 8442
rect 8162 8414 9422 8442
rect 9450 8414 9455 8442
rect 13561 8414 13566 8442
rect 13594 8414 14518 8442
rect 14546 8414 18830 8442
rect 18858 8414 18863 8442
rect 20001 8414 20006 8442
rect 20034 8414 21000 8442
rect 0 8400 400 8414
rect 6734 8330 6762 8414
rect 20600 8400 21000 8414
rect 7625 8358 7630 8386
rect 7658 8358 8862 8386
rect 8890 8358 8895 8386
rect 6729 8302 6734 8330
rect 6762 8302 6767 8330
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 20600 8106 21000 8120
rect 19945 8078 19950 8106
rect 19978 8078 21000 8106
rect 20600 8064 21000 8078
rect 9977 8022 9982 8050
rect 10010 8022 10654 8050
rect 10682 8022 10687 8050
rect 11265 8022 11270 8050
rect 11298 8022 11774 8050
rect 11802 8022 11807 8050
rect 12889 8022 12894 8050
rect 12922 8022 13398 8050
rect 13426 8022 14630 8050
rect 14658 8022 14854 8050
rect 14882 8022 14887 8050
rect 12049 7966 12054 7994
rect 12082 7966 12614 7994
rect 12642 7966 12647 7994
rect 9809 7910 9814 7938
rect 9842 7910 10710 7938
rect 10738 7910 10743 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 20600 7770 21000 7784
rect 20001 7742 20006 7770
rect 20034 7742 21000 7770
rect 20600 7728 21000 7742
rect 14625 7686 14630 7714
rect 14658 7686 18830 7714
rect 18858 7686 18863 7714
rect 6673 7630 6678 7658
rect 6706 7630 8134 7658
rect 8162 7630 8414 7658
rect 8442 7630 8447 7658
rect 9361 7630 9366 7658
rect 9394 7630 10206 7658
rect 10234 7630 10239 7658
rect 8185 7574 8190 7602
rect 8218 7574 8694 7602
rect 8722 7574 8727 7602
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 11377 7238 11382 7266
rect 11410 7238 12894 7266
rect 12922 7238 13062 7266
rect 13090 7238 13095 7266
rect 8185 7126 8190 7154
rect 8218 7126 8414 7154
rect 8442 7126 8918 7154
rect 8946 7126 9478 7154
rect 9506 7126 10374 7154
rect 10402 7126 10407 7154
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 8073 2086 8078 2114
rect 8106 2086 9254 2114
rect 9282 2086 9287 2114
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 12441 1806 12446 1834
rect 12474 1806 13062 1834
rect 13090 1806 13095 1834
rect 8577 1694 8582 1722
rect 8610 1694 9030 1722
rect 9058 1694 9063 1722
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 10150 9646 10178 9674
rect 10150 9422 10178 9450
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 10094 9366 10122 9394
rect 10150 9310 10178 9338
rect 10094 9198 10122 9226
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 10150 8470 10178 8498
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 10150 9674 10178 9679
rect 10150 9450 10178 9646
rect 10150 9417 10178 9422
rect 9904 8638 10064 9394
rect 10094 9394 10122 9399
rect 10094 9226 10122 9366
rect 10094 9193 10122 9198
rect 10150 9338 10178 9343
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 10150 8498 10178 9310
rect 10150 8465 10178 8470
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10808 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10248 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10920 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _116_
timestamp 1698175906
transform 1 0 11648 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform 1 0 7840 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7448 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _119_
timestamp 1698175906
transform -1 0 7616 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7784 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _121_
timestamp 1698175906
transform 1 0 7896 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _122_
timestamp 1698175906
transform 1 0 7504 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8456 0 1 11760
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1698175906
transform -1 0 9296 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11872 0 -1 13328
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _126_
timestamp 1698175906
transform 1 0 11144 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9912 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698175906
transform -1 0 8680 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_
timestamp 1698175906
transform 1 0 7168 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _130_
timestamp 1698175906
transform -1 0 8512 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform 1 0 7952 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _132_
timestamp 1698175906
transform 1 0 7952 0 -1 13328
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _133_
timestamp 1698175906
transform -1 0 7672 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _134_
timestamp 1698175906
transform -1 0 8008 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _135_
timestamp 1698175906
transform -1 0 10136 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _136_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8680 0 1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _137_
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _138_
timestamp 1698175906
transform 1 0 8960 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _139_
timestamp 1698175906
transform -1 0 8736 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _140_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _141_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7000 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _142_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7504 0 -1 9408
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _143_
timestamp 1698175906
transform 1 0 9912 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _144_
timestamp 1698175906
transform 1 0 9128 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _145_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9632 0 -1 7840
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _146_
timestamp 1698175906
transform -1 0 9352 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _147_
timestamp 1698175906
transform -1 0 8456 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _148_
timestamp 1698175906
transform -1 0 7952 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _149_
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _150_
timestamp 1698175906
transform 1 0 10192 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _151_
timestamp 1698175906
transform -1 0 10472 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _152_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8680 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _153_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7672 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _154_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7336 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _155_
timestamp 1698175906
transform -1 0 10472 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _156_
timestamp 1698175906
transform 1 0 9240 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _157_
timestamp 1698175906
transform -1 0 10080 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _158_
timestamp 1698175906
transform -1 0 9128 0 -1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _159_
timestamp 1698175906
transform -1 0 7672 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _160_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7336 0 -1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _161_
timestamp 1698175906
transform 1 0 9856 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _162_
timestamp 1698175906
transform 1 0 11144 0 -1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _163_
timestamp 1698175906
transform 1 0 13496 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _164_
timestamp 1698175906
transform -1 0 13496 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _165_
timestamp 1698175906
transform -1 0 8904 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _166_
timestamp 1698175906
transform -1 0 7952 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _167_
timestamp 1698175906
transform -1 0 13216 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _168_
timestamp 1698175906
transform -1 0 9128 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _169_
timestamp 1698175906
transform 1 0 9912 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _170_
timestamp 1698175906
transform -1 0 10920 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _171_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11480 0 1 10192
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _172_
timestamp 1698175906
transform -1 0 12824 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _173_
timestamp 1698175906
transform 1 0 12432 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _174_
timestamp 1698175906
transform 1 0 10696 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _175_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9744 0 1 10976
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _176_
timestamp 1698175906
transform -1 0 11200 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform -1 0 10472 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _178_
timestamp 1698175906
transform 1 0 10528 0 -1 11760
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _179_
timestamp 1698175906
transform -1 0 10248 0 -1 13328
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _180_
timestamp 1698175906
transform -1 0 10360 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _181_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10192 0 -1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _182_
timestamp 1698175906
transform 1 0 7616 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _183_
timestamp 1698175906
transform -1 0 7616 0 -1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _184_
timestamp 1698175906
transform 1 0 8064 0 1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _185_
timestamp 1698175906
transform 1 0 7896 0 -1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _186_
timestamp 1698175906
transform -1 0 11088 0 -1 13328
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _187_
timestamp 1698175906
transform -1 0 9520 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _188_
timestamp 1698175906
transform 1 0 10808 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _189_
timestamp 1698175906
transform -1 0 11648 0 1 8624
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _190_
timestamp 1698175906
transform 1 0 9072 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _191_
timestamp 1698175906
transform -1 0 7056 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _192_
timestamp 1698175906
transform -1 0 12432 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _193_
timestamp 1698175906
transform -1 0 7560 0 1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _194_
timestamp 1698175906
transform -1 0 12768 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _195_
timestamp 1698175906
transform 1 0 11984 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _196_
timestamp 1698175906
transform -1 0 12264 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _197_
timestamp 1698175906
transform 1 0 10080 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _198_
timestamp 1698175906
transform 1 0 10192 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _199_
timestamp 1698175906
transform 1 0 12320 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _200_
timestamp 1698175906
transform 1 0 10360 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _201_
timestamp 1698175906
transform 1 0 12040 0 1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _202_
timestamp 1698175906
transform 1 0 12544 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _203_
timestamp 1698175906
transform -1 0 13720 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _204_
timestamp 1698175906
transform 1 0 13216 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _205_
timestamp 1698175906
transform -1 0 13384 0 -1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _206_
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _207_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10752 0 1 9408
box -43 -43 1331 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _208_
timestamp 1698175906
transform 1 0 10808 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _209_
timestamp 1698175906
transform 1 0 9632 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _210_
timestamp 1698175906
transform 1 0 13496 0 1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _211_
timestamp 1698175906
transform -1 0 12320 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _212_
timestamp 1698175906
transform 1 0 13944 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _213_
timestamp 1698175906
transform -1 0 13496 0 1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _214_
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _215_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11200 0 -1 10192
box -43 -43 995 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _216_
timestamp 1698175906
transform 1 0 11256 0 -1 9408
box -43 -43 995 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _217_
timestamp 1698175906
transform 1 0 13272 0 1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _218_
timestamp 1698175906
transform -1 0 14112 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _219_
timestamp 1698175906
transform -1 0 13944 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _220_
timestamp 1698175906
transform -1 0 14168 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _221_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10920 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _222_
timestamp 1698175906
transform -1 0 12992 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _223_
timestamp 1698175906
transform 1 0 13048 0 -1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10808 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform -1 0 6496 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform 1 0 9352 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 8624 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 5936 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 5376 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform -1 0 8288 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 12768 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform 1 0 6888 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _236_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform -1 0 6552 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698175906
transform 1 0 6496 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform 1 0 8512 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _240_
timestamp 1698175906
transform -1 0 6552 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _241_
timestamp 1698175906
transform 1 0 11256 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _242_
timestamp 1698175906
transform 1 0 12768 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _243_
timestamp 1698175906
transform 1 0 13720 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _244_
timestamp 1698175906
transform 1 0 13664 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _245_
timestamp 1698175906
transform 1 0 13216 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _246_
timestamp 1698175906
transform 1 0 12768 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _247_
timestamp 1698175906
transform 1 0 12768 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _249_
timestamp 1698175906
transform 1 0 8120 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _250_
timestamp 1698175906
transform -1 0 11256 0 1 14112
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _251_
timestamp 1698175906
transform 1 0 14392 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _252_
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _253_
timestamp 1698175906
transform 1 0 12432 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12768 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 8400 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 7000 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 8904 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 10360 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 7672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 7000 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 8400 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 14616 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform -1 0 8848 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 14280 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 12320 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform -1 0 9184 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 6776 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform 1 0 8120 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform 1 0 10696 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__CLK
timestamp 1698175906
transform 1 0 6776 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__CLK
timestamp 1698175906
transform -1 0 13104 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__CLK
timestamp 1698175906
transform 1 0 14840 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__CLK
timestamp 1698175906
transform 1 0 13104 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__CLK
timestamp 1698175906
transform 1 0 13552 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__CLK
timestamp 1698175906
transform 1 0 14952 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__CLK
timestamp 1698175906
transform 1 0 14616 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__CLK
timestamp 1698175906
transform 1 0 14896 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 9520 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9632 0 -1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 11480 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_165 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9912 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698175906
transform 1 0 10136 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_206
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_210
timestamp 1698175906
transform 1 0 12432 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698175906
transform 1 0 13944 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_168
timestamp 1698175906
transform 1 0 10080 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_200 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11872 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_208
timestamp 1698175906
transform 1 0 12320 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 16128 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 10248 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_146
timestamp 1698175906
transform 1 0 8848 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_184 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10976 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_200
timestamp 1698175906
transform 1 0 11872 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698175906
transform 1 0 12320 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_123
timestamp 1698175906
transform 1 0 7560 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_131
timestamp 1698175906
transform 1 0 8008 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_135
timestamp 1698175906
transform 1 0 8232 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_139
timestamp 1698175906
transform 1 0 8456 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_141
timestamp 1698175906
transform 1 0 8568 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_171
timestamp 1698175906
transform 1 0 10248 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_185
timestamp 1698175906
transform 1 0 11032 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_218
timestamp 1698175906
transform 1 0 12880 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_222
timestamp 1698175906
transform 1 0 13104 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_238
timestamp 1698175906
transform 1 0 14000 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_242
timestamp 1698175906
transform 1 0 14224 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 14336 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698175906
transform 1 0 8456 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_146
timestamp 1698175906
transform 1 0 8848 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_160
timestamp 1698175906
transform 1 0 9632 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_168
timestamp 1698175906
transform 1 0 10080 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_172
timestamp 1698175906
transform 1 0 10304 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_174
timestamp 1698175906
transform 1 0 10416 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_189
timestamp 1698175906
transform 1 0 11256 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_205
timestamp 1698175906
transform 1 0 12152 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 12376 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_251
timestamp 1698175906
transform 1 0 14728 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_255
timestamp 1698175906
transform 1 0 14952 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_271
timestamp 1698175906
transform 1 0 15848 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 16296 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_136
timestamp 1698175906
transform 1 0 8288 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_140
timestamp 1698175906
transform 1 0 8512 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_156
timestamp 1698175906
transform 1 0 9408 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_164
timestamp 1698175906
transform 1 0 9856 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698175906
transform 1 0 10360 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_181
timestamp 1698175906
transform 1 0 10808 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_207
timestamp 1698175906
transform 1 0 12264 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_215
timestamp 1698175906
transform 1 0 12712 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_251
timestamp 1698175906
transform 1 0 14728 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 18648 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 2240 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 4032 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 4480 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_104
timestamp 1698175906
transform 1 0 6496 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_112
timestamp 1698175906
transform 1 0 6944 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_116
timestamp 1698175906
transform 1 0 7168 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_118
timestamp 1698175906
transform 1 0 7280 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 8456 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_151
timestamp 1698175906
transform 1 0 9128 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_159
timestamp 1698175906
transform 1 0 9576 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_169
timestamp 1698175906
transform 1 0 10136 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_177
timestamp 1698175906
transform 1 0 10584 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 12376 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_233
timestamp 1698175906
transform 1 0 13720 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_240
timestamp 1698175906
transform 1 0 14112 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_272
timestamp 1698175906
transform 1 0 15904 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_69
timestamp 1698175906
transform 1 0 4536 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_73
timestamp 1698175906
transform 1 0 4760 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1698175906
transform 1 0 6496 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_111
timestamp 1698175906
transform 1 0 6888 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_115
timestamp 1698175906
transform 1 0 7112 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_123
timestamp 1698175906
transform 1 0 7560 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_131
timestamp 1698175906
transform 1 0 8008 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_141
timestamp 1698175906
transform 1 0 8568 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_149
timestamp 1698175906
transform 1 0 9016 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_208
timestamp 1698175906
transform 1 0 12320 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_224
timestamp 1698175906
transform 1 0 13216 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_228
timestamp 1698175906
transform 1 0 13440 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_242
timestamp 1698175906
transform 1 0 14224 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 14336 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_104
timestamp 1698175906
transform 1 0 6496 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_112
timestamp 1698175906
transform 1 0 6944 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_121
timestamp 1698175906
transform 1 0 7448 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_133
timestamp 1698175906
transform 1 0 8120 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_137
timestamp 1698175906
transform 1 0 8344 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 8456 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_158
timestamp 1698175906
transform 1 0 9520 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698175906
transform 1 0 12208 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_216
timestamp 1698175906
transform 1 0 12768 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_227
timestamp 1698175906
transform 1 0 13384 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_229
timestamp 1698175906
transform 1 0 13496 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_261
timestamp 1698175906
transform 1 0 15288 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698175906
transform 1 0 16184 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 16296 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 18256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 18704 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 4536 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698175906
transform 1 0 4760 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_75
timestamp 1698175906
transform 1 0 4872 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_111
timestamp 1698175906
transform 1 0 6888 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_113
timestamp 1698175906
transform 1 0 7000 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_123
timestamp 1698175906
transform 1 0 7560 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_131
timestamp 1698175906
transform 1 0 8008 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_135
timestamp 1698175906
transform 1 0 8232 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_168
timestamp 1698175906
transform 1 0 10080 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_179
timestamp 1698175906
transform 1 0 10696 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_210
timestamp 1698175906
transform 1 0 12432 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_217
timestamp 1698175906
transform 1 0 12824 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_219
timestamp 1698175906
transform 1 0 12936 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_238
timestamp 1698175906
transform 1 0 14000 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_242
timestamp 1698175906
transform 1 0 14224 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 14336 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_252
timestamp 1698175906
transform 1 0 14784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_284
timestamp 1698175906
transform 1 0 16576 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_300
timestamp 1698175906
transform 1 0 17472 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_308
timestamp 1698175906
transform 1 0 17920 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698175906
transform 1 0 18144 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698175906
transform 1 0 18256 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 2240 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 4032 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 4480 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_104
timestamp 1698175906
transform 1 0 6496 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_108
timestamp 1698175906
transform 1 0 6720 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_132
timestamp 1698175906
transform 1 0 8064 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_155
timestamp 1698175906
transform 1 0 9352 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_159
timestamp 1698175906
transform 1 0 9576 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_175
timestamp 1698175906
transform 1 0 10472 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_220
timestamp 1698175906
transform 1 0 12992 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_230
timestamp 1698175906
transform 1 0 13552 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_232
timestamp 1698175906
transform 1 0 13664 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_262
timestamp 1698175906
transform 1 0 15344 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 16240 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 18256 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 18704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698175906
transform 1 0 2240 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698175906
transform 1 0 2464 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 4536 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 4760 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 4872 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_111
timestamp 1698175906
transform 1 0 6888 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698175906
transform 1 0 14280 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_104
timestamp 1698175906
transform 1 0 6496 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_112
timestamp 1698175906
transform 1 0 6944 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_116
timestamp 1698175906
transform 1 0 7168 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_118
timestamp 1698175906
transform 1 0 7280 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_135
timestamp 1698175906
transform 1 0 8232 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698175906
transform 1 0 8456 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_142
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_146
timestamp 1698175906
transform 1 0 8848 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_156
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_217
timestamp 1698175906
transform 1 0 12824 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_230
timestamp 1698175906
transform 1 0 13552 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_234
timestamp 1698175906
transform 1 0 13776 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_241
timestamp 1698175906
transform 1 0 14168 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_273
timestamp 1698175906
transform 1 0 15960 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698175906
transform 1 0 16184 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 16296 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 20048 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 20160 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_111
timestamp 1698175906
transform 1 0 6888 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_115
timestamp 1698175906
transform 1 0 7112 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_117
timestamp 1698175906
transform 1 0 7224 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_144
timestamp 1698175906
transform 1 0 8736 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_151
timestamp 1698175906
transform 1 0 9128 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_159
timestamp 1698175906
transform 1 0 9576 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_161
timestamp 1698175906
transform 1 0 9688 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_191
timestamp 1698175906
transform 1 0 11368 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_199
timestamp 1698175906
transform 1 0 11816 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_214
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_252
timestamp 1698175906
transform 1 0 14784 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_256
timestamp 1698175906
transform 1 0 15008 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_288
timestamp 1698175906
transform 1 0 16800 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_304
timestamp 1698175906
transform 1 0 17696 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_312
timestamp 1698175906
transform 1 0 18144 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698175906
transform 1 0 18256 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_80
timestamp 1698175906
transform 1 0 5152 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_113
timestamp 1698175906
transform 1 0 7000 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_115
timestamp 1698175906
transform 1 0 7112 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_158
timestamp 1698175906
transform 1 0 9520 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_162
timestamp 1698175906
transform 1 0 9744 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_186
timestamp 1698175906
transform 1 0 11088 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_202
timestamp 1698175906
transform 1 0 11984 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_220
timestamp 1698175906
transform 1 0 12992 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_253
timestamp 1698175906
transform 1 0 14840 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_257
timestamp 1698175906
transform 1 0 15064 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698175906
transform 1 0 15960 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 16184 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 16296 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_115
timestamp 1698175906
transform 1 0 7112 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_119
timestamp 1698175906
transform 1 0 7336 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_149
timestamp 1698175906
transform 1 0 9016 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_165
timestamp 1698175906
transform 1 0 9912 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_206
timestamp 1698175906
transform 1 0 12208 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_210
timestamp 1698175906
transform 1 0 12432 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_218
timestamp 1698175906
transform 1 0 12880 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_222
timestamp 1698175906
transform 1 0 13104 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_224
timestamp 1698175906
transform 1 0 13216 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_234
timestamp 1698175906
transform 1 0 13776 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698175906
transform 1 0 14224 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 14336 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_88
timestamp 1698175906
transform 1 0 5600 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_92
timestamp 1698175906
transform 1 0 5824 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_123
timestamp 1698175906
transform 1 0 7560 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_127
timestamp 1698175906
transform 1 0 7784 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_133
timestamp 1698175906
transform 1 0 8120 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_137
timestamp 1698175906
transform 1 0 8344 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 8456 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_174
timestamp 1698175906
transform 1 0 10416 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_178
timestamp 1698175906
transform 1 0 10640 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_192
timestamp 1698175906
transform 1 0 11424 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698175906
transform 1 0 12320 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 16128 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_123
timestamp 1698175906
transform 1 0 7560 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_131
timestamp 1698175906
transform 1 0 8008 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_135
timestamp 1698175906
transform 1 0 8232 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_137
timestamp 1698175906
transform 1 0 8344 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_143
timestamp 1698175906
transform 1 0 8680 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_177
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_209
timestamp 1698175906
transform 1 0 12376 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_215
timestamp 1698175906
transform 1 0 12712 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_251
timestamp 1698175906
transform 1 0 14728 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_104
timestamp 1698175906
transform 1 0 6496 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_120
timestamp 1698175906
transform 1 0 7392 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 8456 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_147
timestamp 1698175906
transform 1 0 8904 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_158
timestamp 1698175906
transform 1 0 9520 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_171
timestamp 1698175906
transform 1 0 10248 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_175
timestamp 1698175906
transform 1 0 10472 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_186
timestamp 1698175906
transform 1 0 11088 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_200
timestamp 1698175906
transform 1 0 11872 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698175906
transform 1 0 12320 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_241
timestamp 1698175906
transform 1 0 14168 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_245
timestamp 1698175906
transform 1 0 14392 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 16184 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 16296 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_136
timestamp 1698175906
transform 1 0 8288 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698175906
transform 1 0 10360 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_216
timestamp 1698175906
transform 1 0 12768 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_218
timestamp 1698175906
transform 1 0 12880 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_234
timestamp 1698175906
transform 1 0 13776 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 14224 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 18648 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_104
timestamp 1698175906
transform 1 0 6496 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_108
timestamp 1698175906
transform 1 0 6720 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_110
timestamp 1698175906
transform 1 0 6832 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_146
timestamp 1698175906
transform 1 0 8848 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_183
timestamp 1698175906
transform 1 0 10920 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_199
timestamp 1698175906
transform 1 0 11816 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698175906
transform 1 0 12264 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 12376 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_216
timestamp 1698175906
transform 1 0 12768 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_189
timestamp 1698175906
transform 1 0 11256 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_221
timestamp 1698175906
transform 1 0 13048 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_237
timestamp 1698175906
transform 1 0 13944 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_333
timestamp 1698175906
transform 1 0 19320 0 1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_341
timestamp 1698175906
transform 1 0 19768 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_123
timestamp 1698175906
transform 1 0 7560 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_131
timestamp 1698175906
transform 1 0 8008 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_159
timestamp 1698175906
transform 1 0 9576 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_203
timestamp 1698175906
transform 1 0 12040 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_237
timestamp 1698175906
transform 1 0 13944 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_150
timestamp 1698175906
transform 1 0 9072 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_154
timestamp 1698175906
transform 1 0 9296 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 14000 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 15792 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 16240 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita13_26 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19992 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18760 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 18760 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 8456 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 10640 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 12488 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 18760 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 18760 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 18760 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform -1 0 2240 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 10808 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform -1 0 2240 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 12488 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 8736 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 18760 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 2240 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 8120 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform -1 0 10808 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13776 400 13832 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 20600 17136 21000 17192 0 FreeSans 224 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 20600 9072 21000 9128 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 20600 8400 21000 8456 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 8400 0 8456 400 0 FreeSans 224 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 12432 20600 12488 21000 0 FreeSans 224 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 8064 0 8120 400 0 FreeSans 224 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 10416 20600 10472 21000 0 FreeSans 224 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 20600 7728 21000 7784 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 20600 8064 21000 8120 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 20600 9744 21000 9800 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 0 10080 400 10136 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 10752 20600 10808 21000 0 FreeSans 224 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 9744 400 9800 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 12432 0 12488 400 0 FreeSans 224 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 11760 20600 11816 21000 0 FreeSans 224 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 8736 20600 8792 21000 0 FreeSans 224 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 8400 400 8456 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 0 8736 400 8792 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 8064 20600 8120 21000 0 FreeSans 224 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 10080 20600 10136 21000 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 12096 20600 12152 21000 0 FreeSans 224 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 11284 13356 11284 13356 0 _000_
rlabel metal2 7420 13132 7420 13132 0 _001_
rlabel metal2 6020 9100 6020 9100 0 _002_
rlabel metal2 9828 9240 9828 9240 0 _003_
rlabel metal2 9100 7084 9100 7084 0 _004_
rlabel metal2 7812 12152 7812 12152 0 _005_
rlabel metal3 6664 10836 6664 10836 0 _006_
rlabel metal2 7812 8316 7812 8316 0 _007_
rlabel metal2 13244 13104 13244 13104 0 _008_
rlabel metal2 7532 13636 7532 13636 0 _009_
rlabel metal3 12852 12628 12852 12628 0 _010_
rlabel metal2 11032 11900 11032 11900 0 _011_
rlabel metal2 9660 13748 9660 13748 0 _012_
rlabel metal2 6076 10220 6076 10220 0 _013_
rlabel metal2 6972 7868 6972 7868 0 _014_
rlabel metal3 9184 13244 9184 13244 0 _015_
rlabel metal2 7196 9632 7196 9632 0 _016_
rlabel metal2 11732 7434 11732 7434 0 _017_
rlabel metal2 13216 7700 13216 7700 0 _018_
rlabel metal2 13748 9870 13748 9870 0 _019_
rlabel metal2 13244 9352 13244 9352 0 _020_
rlabel metal2 13692 11816 13692 11816 0 _021_
rlabel metal2 13244 8400 13244 8400 0 _022_
rlabel metal2 13272 10892 13272 10892 0 _023_
rlabel metal2 13524 13636 13524 13636 0 _024_
rlabel metal3 8260 13188 8260 13188 0 _025_
rlabel metal3 12768 13468 12768 13468 0 _026_
rlabel metal3 8680 11116 8680 11116 0 _027_
rlabel metal2 10948 9436 10948 9436 0 _028_
rlabel metal2 11032 11284 11032 11284 0 _029_
rlabel metal2 12348 10164 12348 10164 0 _030_
rlabel metal2 12656 10668 12656 10668 0 _031_
rlabel metal2 10836 11928 10836 11928 0 _032_
rlabel metal2 10332 9856 10332 9856 0 _033_
rlabel metal3 10668 9996 10668 9996 0 _034_
rlabel metal2 10220 10500 10220 10500 0 _035_
rlabel metal2 10192 13468 10192 13468 0 _036_
rlabel metal2 8036 9968 8036 9968 0 _037_
rlabel metal3 7532 9940 7532 9940 0 _038_
rlabel metal2 8288 8316 8288 8316 0 _039_
rlabel metal3 10108 13076 10108 13076 0 _040_
rlabel metal2 11172 8204 11172 8204 0 _041_
rlabel metal2 11620 9576 11620 9576 0 _042_
rlabel metal2 13580 11396 13580 11396 0 _043_
rlabel metal2 7364 9744 7364 9744 0 _044_
rlabel metal2 7476 10108 7476 10108 0 _045_
rlabel metal2 12628 7868 12628 7868 0 _046_
rlabel metal3 13832 8484 13832 8484 0 _047_
rlabel metal2 10276 9828 10276 9828 0 _048_
rlabel metal2 12796 10052 12796 10052 0 _049_
rlabel metal3 14336 10780 14336 10780 0 _050_
rlabel metal2 11256 9996 11256 9996 0 _051_
rlabel metal3 12768 9604 12768 9604 0 _052_
rlabel metal2 12964 9352 12964 9352 0 _053_
rlabel metal2 13188 8876 13188 8876 0 _054_
rlabel metal2 13804 9156 13804 9156 0 _055_
rlabel metal3 14336 9604 14336 9604 0 _056_
rlabel metal2 11676 9492 11676 9492 0 _057_
rlabel metal3 12096 9492 12096 9492 0 _058_
rlabel metal3 13524 9128 13524 9128 0 _059_
rlabel metal3 12656 10836 12656 10836 0 _060_
rlabel metal2 14056 8932 14056 8932 0 _061_
rlabel metal2 14728 11172 14728 11172 0 _062_
rlabel metal2 11816 9212 11816 9212 0 _063_
rlabel metal2 13468 11368 13468 11368 0 _064_
rlabel metal2 13860 8652 13860 8652 0 _065_
rlabel metal2 13692 10780 13692 10780 0 _066_
rlabel metal2 11284 10836 11284 10836 0 _067_
rlabel metal3 13048 10052 13048 10052 0 _068_
rlabel metal2 10220 8848 10220 8848 0 _069_
rlabel metal2 10920 8820 10920 8820 0 _070_
rlabel metal2 11396 9072 11396 9072 0 _071_
rlabel metal2 12124 11480 12124 11480 0 _072_
rlabel metal2 7364 11396 7364 11396 0 _073_
rlabel metal2 7532 11480 7532 11480 0 _074_
rlabel metal2 7532 10920 7532 10920 0 _075_
rlabel metal2 8092 9968 8092 9968 0 _076_
rlabel metal3 8204 11956 8204 11956 0 _077_
rlabel metal2 9324 10332 9324 10332 0 _078_
rlabel metal2 8372 13048 8372 13048 0 _079_
rlabel metal3 12404 13524 12404 13524 0 _080_
rlabel metal2 11284 13132 11284 13132 0 _081_
rlabel metal2 9156 9464 9156 9464 0 _082_
rlabel metal3 8344 12684 8344 12684 0 _083_
rlabel metal2 7420 11536 7420 11536 0 _084_
rlabel metal2 7924 8736 7924 8736 0 _085_
rlabel metal3 7924 11060 7924 11060 0 _086_
rlabel metal3 7896 13132 7896 13132 0 _087_
rlabel metal2 7532 9660 7532 9660 0 _088_
rlabel metal2 10164 9520 10164 9520 0 _089_
rlabel metal2 7756 9436 7756 9436 0 _090_
rlabel metal2 6804 9044 6804 9044 0 _091_
rlabel metal2 11144 10388 11144 10388 0 _092_
rlabel metal2 11900 10080 11900 10080 0 _093_
rlabel metal2 7196 9240 7196 9240 0 _094_
rlabel metal2 7588 9184 7588 9184 0 _095_
rlabel metal2 10220 7868 10220 7868 0 _096_
rlabel metal2 9380 8988 9380 8988 0 _097_
rlabel metal2 9212 7210 9212 7210 0 _098_
rlabel metal2 8204 11956 8204 11956 0 _099_
rlabel metal2 7364 10864 7364 10864 0 _100_
rlabel metal2 10808 11116 10808 11116 0 _101_
rlabel metal2 10388 12152 10388 12152 0 _102_
rlabel metal2 10192 11844 10192 11844 0 _103_
rlabel metal2 8428 12796 8428 12796 0 _104_
rlabel metal2 9996 9688 9996 9688 0 _105_
rlabel metal2 9716 10052 9716 10052 0 _106_
rlabel metal2 8932 8960 8932 8960 0 _107_
rlabel metal3 8260 8372 8260 8372 0 _108_
rlabel metal2 7420 10178 7420 10178 0 _109_
rlabel metal2 10864 13188 10864 13188 0 _110_
rlabel metal3 12376 12460 12376 12460 0 _111_
rlabel metal2 5796 12348 5796 12348 0 clk
rlabel metal2 11564 10556 11564 10556 0 clknet_0_clk
rlabel metal2 10696 13580 10696 13580 0 clknet_1_0__leaf_clk
rlabel metal2 14644 12964 14644 12964 0 clknet_1_1__leaf_clk
rlabel metal2 10808 7644 10808 7644 0 dut13.count\[0\]
rlabel metal2 10164 7434 10164 7434 0 dut13.count\[1\]
rlabel metal2 7476 12264 7476 12264 0 dut13.count\[2\]
rlabel metal2 7308 11732 7308 11732 0 dut13.count\[3\]
rlabel metal2 15204 8960 15204 8960 0 net1
rlabel metal2 18844 7868 18844 7868 0 net10
rlabel metal2 14532 8036 14532 8036 0 net11
rlabel metal2 14644 9744 14644 9744 0 net12
rlabel metal3 3178 10388 3178 10388 0 net13
rlabel metal2 10836 14672 10836 14672 0 net14
rlabel metal3 3178 9996 3178 9996 0 net15
rlabel metal2 12628 2982 12628 2982 0 net16
rlabel metal2 12208 15960 12208 15960 0 net17
rlabel metal2 14084 13048 14084 13048 0 net18
rlabel metal2 8680 13804 8680 13804 0 net19
rlabel metal2 14644 11312 14644 11312 0 net2
rlabel metal2 14336 12796 14336 12796 0 net20
rlabel metal2 6748 8204 6748 8204 0 net21
rlabel metal3 3178 8820 3178 8820 0 net22
rlabel metal2 8232 13580 8232 13580 0 net23
rlabel metal2 10724 13860 10724 13860 0 net24
rlabel metal2 12684 16044 12684 16044 0 net25
rlabel metal2 20132 17248 20132 17248 0 net26
rlabel metal2 13972 8680 13972 8680 0 net3
rlabel metal2 14028 11060 14028 11060 0 net4
rlabel metal2 8456 1764 8456 1764 0 net5
rlabel metal2 10948 19012 10948 19012 0 net6
rlabel metal2 12432 13580 12432 13580 0 net7
rlabel metal2 8204 8288 8204 8288 0 net8
rlabel metal2 10780 14168 10780 14168 0 net9
rlabel metal3 20321 9100 20321 9100 0 segm[10]
rlabel metal3 20321 11452 20321 11452 0 segm[11]
rlabel metal2 20020 8652 20020 8652 0 segm[12]
rlabel metal2 20020 11172 20020 11172 0 segm[13]
rlabel metal2 8428 427 8428 427 0 segm[1]
rlabel metal2 11116 19873 11116 19873 0 segm[2]
rlabel metal2 12460 19481 12460 19481 0 segm[3]
rlabel metal2 8092 1239 8092 1239 0 segm[4]
rlabel metal2 10444 19481 10444 19481 0 segm[5]
rlabel metal2 20020 7924 20020 7924 0 segm[6]
rlabel metal2 19964 8232 19964 8232 0 segm[7]
rlabel metal2 20020 9828 20020 9828 0 segm[8]
rlabel metal3 679 10108 679 10108 0 segm[9]
rlabel metal2 10780 19677 10780 19677 0 sel[0]
rlabel metal3 679 9772 679 9772 0 sel[10]
rlabel metal2 12460 1099 12460 1099 0 sel[11]
rlabel metal2 11788 19873 11788 19873 0 sel[1]
rlabel metal2 20020 12908 20020 12908 0 sel[2]
rlabel metal2 8764 19873 8764 19873 0 sel[3]
rlabel metal2 20020 13356 20020 13356 0 sel[4]
rlabel metal3 679 8428 679 8428 0 sel[5]
rlabel metal3 679 8764 679 8764 0 sel[6]
rlabel metal2 8092 19481 8092 19481 0 sel[7]
rlabel metal2 10108 19593 10108 19593 0 sel[8]
rlabel metal2 12124 19677 12124 19677 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
