magic
tech gf180mcuD
magscale 1 5
timestamp 1699643347
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9031 19137 9057 19143
rect 9031 19105 9057 19111
rect 11215 19137 11241 19143
rect 11215 19105 11241 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 8521 18999 8527 19025
rect 8553 18999 8559 19025
rect 10873 18999 10879 19025
rect 10905 18999 10911 19025
rect 12385 18999 12391 19025
rect 12417 18999 12423 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 9927 18745 9953 18751
rect 9927 18713 9953 18719
rect 11383 18745 11409 18751
rect 11383 18713 11409 18719
rect 9417 18607 9423 18633
rect 9449 18607 9455 18633
rect 10985 18607 10991 18633
rect 11017 18607 11023 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 7967 13873 7993 13879
rect 7967 13841 7993 13847
rect 9311 13873 9337 13879
rect 9311 13841 9337 13847
rect 7911 13817 7937 13823
rect 7911 13785 7937 13791
rect 9255 13817 9281 13823
rect 9255 13785 9281 13791
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 967 13593 993 13599
rect 7345 13567 7351 13593
rect 7377 13567 7383 13593
rect 8409 13567 8415 13593
rect 8441 13567 8447 13593
rect 8969 13567 8975 13593
rect 9001 13567 9007 13593
rect 10033 13567 10039 13593
rect 10065 13567 10071 13593
rect 967 13561 993 13567
rect 2137 13511 2143 13537
rect 2169 13511 2175 13537
rect 7009 13511 7015 13537
rect 7041 13511 7047 13537
rect 8633 13511 8639 13537
rect 8665 13511 8671 13537
rect 10985 13511 10991 13537
rect 11017 13511 11023 13537
rect 10263 13481 10289 13487
rect 10873 13455 10879 13481
rect 10905 13455 10911 13481
rect 10263 13449 10289 13455
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 8247 13257 8273 13263
rect 8247 13225 8273 13231
rect 8303 13257 8329 13263
rect 8303 13225 8329 13231
rect 9255 13257 9281 13263
rect 9255 13225 9281 13231
rect 9311 13257 9337 13263
rect 9311 13225 9337 13231
rect 13063 13201 13089 13207
rect 13063 13169 13089 13175
rect 7463 13145 7489 13151
rect 2137 13119 2143 13145
rect 2169 13119 2175 13145
rect 7233 13119 7239 13145
rect 7265 13119 7271 13145
rect 7463 13113 7489 13119
rect 8135 13145 8161 13151
rect 8135 13113 8161 13119
rect 8191 13145 8217 13151
rect 9143 13145 9169 13151
rect 8409 13119 8415 13145
rect 8441 13119 8447 13145
rect 8191 13113 8217 13119
rect 9143 13113 9169 13119
rect 9199 13145 9225 13151
rect 9199 13113 9225 13119
rect 9367 13145 9393 13151
rect 13119 13145 13145 13151
rect 9585 13119 9591 13145
rect 9617 13119 9623 13145
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 9367 13113 9393 13119
rect 13119 13113 13145 13119
rect 8751 13089 8777 13095
rect 11271 13089 11297 13095
rect 5777 13063 5783 13089
rect 5809 13063 5815 13089
rect 6841 13063 6847 13089
rect 6873 13063 6879 13089
rect 9977 13063 9983 13089
rect 10009 13063 10015 13089
rect 11041 13063 11047 13089
rect 11073 13063 11079 13089
rect 8751 13057 8777 13063
rect 11271 13057 11297 13063
rect 11495 13089 11521 13095
rect 11495 13057 11521 13063
rect 12671 13089 12697 13095
rect 12671 13057 12697 13063
rect 13343 13089 13369 13095
rect 13343 13057 13369 13063
rect 967 13033 993 13039
rect 967 13001 993 13007
rect 13063 13033 13089 13039
rect 13063 13001 13089 13007
rect 20007 13033 20033 13039
rect 20007 13001 20033 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 10039 12809 10065 12815
rect 9809 12783 9815 12809
rect 9841 12783 9847 12809
rect 12385 12783 12391 12809
rect 12417 12783 12423 12809
rect 14009 12783 14015 12809
rect 14041 12783 14047 12809
rect 10039 12777 10065 12783
rect 6903 12753 6929 12759
rect 6903 12721 6929 12727
rect 7183 12753 7209 12759
rect 7183 12721 7209 12727
rect 7351 12753 7377 12759
rect 7351 12721 7377 12727
rect 7519 12753 7545 12759
rect 7519 12721 7545 12727
rect 9983 12753 10009 12759
rect 9983 12721 10009 12727
rect 10319 12753 10345 12759
rect 10319 12721 10345 12727
rect 10599 12753 10625 12759
rect 10929 12727 10935 12753
rect 10961 12727 10967 12753
rect 12609 12727 12615 12753
rect 12641 12727 12647 12753
rect 10599 12721 10625 12727
rect 7015 12697 7041 12703
rect 7015 12665 7041 12671
rect 7071 12697 7097 12703
rect 7071 12665 7097 12671
rect 7295 12697 7321 12703
rect 7295 12665 7321 12671
rect 9647 12697 9673 12703
rect 9647 12665 9673 12671
rect 10711 12697 10737 12703
rect 10711 12665 10737 12671
rect 10767 12697 10793 12703
rect 11321 12671 11327 12697
rect 11353 12671 11359 12697
rect 12945 12671 12951 12697
rect 12977 12671 12983 12697
rect 10767 12665 10793 12671
rect 7575 12641 7601 12647
rect 7575 12609 7601 12615
rect 7687 12641 7713 12647
rect 7687 12609 7713 12615
rect 9759 12641 9785 12647
rect 9759 12609 9785 12615
rect 10095 12641 10121 12647
rect 10095 12609 10121 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 11271 12473 11297 12479
rect 9305 12447 9311 12473
rect 9337 12447 9343 12473
rect 11271 12441 11297 12447
rect 11775 12473 11801 12479
rect 11775 12441 11801 12447
rect 12671 12473 12697 12479
rect 12671 12441 12697 12447
rect 10319 12417 10345 12423
rect 10319 12385 10345 12391
rect 11439 12417 11465 12423
rect 11439 12385 11465 12391
rect 11943 12417 11969 12423
rect 11943 12385 11969 12391
rect 7855 12361 7881 12367
rect 7457 12335 7463 12361
rect 7489 12335 7495 12361
rect 7681 12335 7687 12361
rect 7713 12335 7719 12361
rect 7855 12329 7881 12335
rect 7967 12361 7993 12367
rect 11103 12361 11129 12367
rect 9417 12335 9423 12361
rect 9449 12335 9455 12361
rect 7967 12329 7993 12335
rect 11103 12329 11129 12335
rect 11271 12361 11297 12367
rect 11271 12329 11297 12335
rect 11663 12361 11689 12367
rect 11663 12329 11689 12335
rect 11719 12361 11745 12367
rect 11719 12329 11745 12335
rect 11831 12361 11857 12367
rect 12833 12335 12839 12361
rect 12865 12335 12871 12361
rect 18825 12335 18831 12361
rect 18857 12335 18863 12361
rect 11831 12329 11857 12335
rect 7911 12305 7937 12311
rect 6057 12279 6063 12305
rect 6089 12279 6095 12305
rect 7121 12279 7127 12305
rect 7153 12279 7159 12305
rect 7911 12273 7937 12279
rect 8191 12305 8217 12311
rect 8191 12273 8217 12279
rect 10207 12305 10233 12311
rect 10879 12305 10905 12311
rect 10369 12279 10375 12305
rect 10401 12279 10407 12305
rect 13225 12279 13231 12305
rect 13257 12279 13263 12305
rect 14289 12279 14295 12305
rect 14321 12279 14327 12305
rect 10207 12273 10233 12279
rect 10879 12273 10905 12279
rect 20007 12249 20033 12255
rect 20007 12217 20033 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 11215 12081 11241 12087
rect 11215 12049 11241 12055
rect 20007 12025 20033 12031
rect 12889 11999 12895 12025
rect 12921 11999 12927 12025
rect 20007 11993 20033 11999
rect 9591 11969 9617 11975
rect 8801 11943 8807 11969
rect 8833 11943 8839 11969
rect 9473 11943 9479 11969
rect 9505 11943 9511 11969
rect 9591 11937 9617 11943
rect 9983 11969 10009 11975
rect 9983 11937 10009 11943
rect 10095 11969 10121 11975
rect 12727 11969 12753 11975
rect 13063 11969 13089 11975
rect 10985 11943 10991 11969
rect 11017 11943 11023 11969
rect 11545 11943 11551 11969
rect 11577 11943 11583 11969
rect 12945 11943 12951 11969
rect 12977 11943 12983 11969
rect 10095 11937 10121 11943
rect 12727 11937 12753 11943
rect 13063 11937 13089 11943
rect 13399 11969 13425 11975
rect 13399 11937 13425 11943
rect 13623 11969 13649 11975
rect 13623 11937 13649 11943
rect 13735 11969 13761 11975
rect 14065 11943 14071 11969
rect 14097 11943 14103 11969
rect 18825 11943 18831 11969
rect 18857 11943 18863 11969
rect 13735 11937 13761 11943
rect 9647 11913 9673 11919
rect 9647 11881 9673 11887
rect 10375 11913 10401 11919
rect 12615 11913 12641 11919
rect 11265 11887 11271 11913
rect 11297 11887 11303 11913
rect 10375 11881 10401 11887
rect 12615 11881 12641 11887
rect 12839 11913 12865 11919
rect 12839 11881 12865 11887
rect 13287 11913 13313 11919
rect 13287 11881 13313 11887
rect 13567 11913 13593 11919
rect 13567 11881 13593 11887
rect 13847 11913 13873 11919
rect 14177 11887 14183 11913
rect 14209 11887 14215 11913
rect 13847 11881 13873 11887
rect 7631 11857 7657 11863
rect 10207 11857 10233 11863
rect 8689 11831 8695 11857
rect 8721 11831 8727 11857
rect 9809 11831 9815 11857
rect 9841 11831 9847 11857
rect 7631 11825 7657 11831
rect 10207 11825 10233 11831
rect 10319 11857 10345 11863
rect 13231 11857 13257 11863
rect 11433 11831 11439 11857
rect 11465 11831 11471 11857
rect 10319 11825 10345 11831
rect 13231 11825 13257 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 13399 11689 13425 11695
rect 13399 11657 13425 11663
rect 7183 11633 7209 11639
rect 9081 11607 9087 11633
rect 9113 11607 9119 11633
rect 9305 11607 9311 11633
rect 9337 11607 9343 11633
rect 7183 11601 7209 11607
rect 7687 11577 7713 11583
rect 7569 11551 7575 11577
rect 7601 11551 7607 11577
rect 7687 11545 7713 11551
rect 7743 11577 7769 11583
rect 7743 11545 7769 11551
rect 7799 11577 7825 11583
rect 7905 11551 7911 11577
rect 7937 11551 7943 11577
rect 9361 11551 9367 11577
rect 9393 11551 9399 11577
rect 11881 11551 11887 11577
rect 11913 11551 11919 11577
rect 7799 11545 7825 11551
rect 8303 11521 8329 11527
rect 8303 11489 8329 11495
rect 8751 11521 8777 11527
rect 10089 11495 10095 11521
rect 10121 11495 10127 11521
rect 8751 11489 8777 11495
rect 7127 11465 7153 11471
rect 7127 11433 7153 11439
rect 7295 11465 7321 11471
rect 7295 11433 7321 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 8863 11297 8889 11303
rect 8863 11265 8889 11271
rect 967 11241 993 11247
rect 8415 11241 8441 11247
rect 13343 11241 13369 11247
rect 8185 11215 8191 11241
rect 8217 11215 8223 11241
rect 12609 11215 12615 11241
rect 12641 11215 12647 11241
rect 967 11209 993 11215
rect 8415 11209 8441 11215
rect 13343 11209 13369 11215
rect 8359 11185 8385 11191
rect 9087 11185 9113 11191
rect 9983 11185 10009 11191
rect 2137 11159 2143 11185
rect 2169 11159 2175 11185
rect 6785 11159 6791 11185
rect 6817 11159 6823 11185
rect 8633 11159 8639 11185
rect 8665 11159 8671 11185
rect 9305 11159 9311 11185
rect 9337 11159 9343 11185
rect 9697 11159 9703 11185
rect 9729 11159 9735 11185
rect 9921 11159 9927 11185
rect 9953 11159 9959 11185
rect 8359 11153 8385 11159
rect 9087 11153 9113 11159
rect 9983 11153 10009 11159
rect 10823 11185 10849 11191
rect 10823 11153 10849 11159
rect 11047 11185 11073 11191
rect 11047 11153 11073 11159
rect 12895 11185 12921 11191
rect 12895 11153 12921 11159
rect 13007 11185 13033 11191
rect 13007 11153 13033 11159
rect 8807 11129 8833 11135
rect 7121 11103 7127 11129
rect 7153 11103 7159 11129
rect 8807 11097 8833 11103
rect 10207 11129 10233 11135
rect 10207 11097 10233 11103
rect 10655 11129 10681 11135
rect 11377 11103 11383 11129
rect 11409 11103 11415 11129
rect 10655 11097 10681 11103
rect 8471 11073 8497 11079
rect 8471 11041 8497 11047
rect 10263 11073 10289 11079
rect 10263 11041 10289 11047
rect 11215 11073 11241 11079
rect 11215 11041 11241 11047
rect 11551 11073 11577 11079
rect 12615 11073 12641 11079
rect 11713 11047 11719 11073
rect 11745 11047 11751 11073
rect 11551 11041 11577 11047
rect 12615 11041 12641 11047
rect 12727 11073 12753 11079
rect 12727 11041 12753 11047
rect 13063 11073 13089 11079
rect 13063 11041 13089 11047
rect 13175 11073 13201 11079
rect 13175 11041 13201 11047
rect 20119 11073 20145 11079
rect 20119 11041 20145 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 8023 10905 8049 10911
rect 8023 10873 8049 10879
rect 8079 10905 8105 10911
rect 8079 10873 8105 10879
rect 9087 10905 9113 10911
rect 9087 10873 9113 10879
rect 7911 10849 7937 10855
rect 13063 10849 13089 10855
rect 6673 10823 6679 10849
rect 6705 10823 6711 10849
rect 8913 10823 8919 10849
rect 8945 10823 8951 10849
rect 10425 10823 10431 10849
rect 10457 10823 10463 10849
rect 10817 10823 10823 10849
rect 10849 10823 10855 10849
rect 7911 10817 7937 10823
rect 13063 10817 13089 10823
rect 7239 10793 7265 10799
rect 2137 10767 2143 10793
rect 2169 10767 2175 10793
rect 7009 10767 7015 10793
rect 7041 10767 7047 10793
rect 7239 10761 7265 10767
rect 7351 10793 7377 10799
rect 7351 10761 7377 10767
rect 7463 10793 7489 10799
rect 7743 10793 7769 10799
rect 7569 10767 7575 10793
rect 7601 10767 7607 10793
rect 7463 10761 7489 10767
rect 7743 10761 7769 10767
rect 8135 10793 8161 10799
rect 8135 10761 8161 10767
rect 9871 10793 9897 10799
rect 11719 10793 11745 10799
rect 10649 10767 10655 10793
rect 10681 10767 10687 10793
rect 10873 10767 10879 10793
rect 10905 10767 10911 10793
rect 9871 10761 9897 10767
rect 11719 10761 11745 10767
rect 12727 10793 12753 10799
rect 12727 10761 12753 10767
rect 12839 10793 12865 10799
rect 12839 10761 12865 10767
rect 12951 10793 12977 10799
rect 13281 10767 13287 10793
rect 13313 10767 13319 10793
rect 18825 10767 18831 10793
rect 18857 10767 18863 10793
rect 12951 10761 12977 10767
rect 7295 10737 7321 10743
rect 5609 10711 5615 10737
rect 5641 10711 5647 10737
rect 7295 10705 7321 10711
rect 9591 10737 9617 10743
rect 13617 10711 13623 10737
rect 13649 10711 13655 10737
rect 14681 10711 14687 10737
rect 14713 10711 14719 10737
rect 9591 10705 9617 10711
rect 967 10681 993 10687
rect 967 10649 993 10655
rect 13007 10681 13033 10687
rect 13007 10649 13033 10655
rect 20007 10681 20033 10687
rect 20007 10649 20033 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 7015 10513 7041 10519
rect 7015 10481 7041 10487
rect 7463 10513 7489 10519
rect 7463 10481 7489 10487
rect 9927 10513 9953 10519
rect 9927 10481 9953 10487
rect 6791 10457 6817 10463
rect 4993 10431 4999 10457
rect 5025 10431 5031 10457
rect 6057 10431 6063 10457
rect 6089 10431 6095 10457
rect 6791 10425 6817 10431
rect 6959 10457 6985 10463
rect 6959 10425 6985 10431
rect 9871 10457 9897 10463
rect 10145 10431 10151 10457
rect 10177 10431 10183 10457
rect 9871 10425 9897 10431
rect 7239 10401 7265 10407
rect 6449 10375 6455 10401
rect 6481 10375 6487 10401
rect 7239 10369 7265 10375
rect 7519 10401 7545 10407
rect 7519 10369 7545 10375
rect 8247 10401 8273 10407
rect 13735 10401 13761 10407
rect 10313 10375 10319 10401
rect 10345 10375 10351 10401
rect 10929 10375 10935 10401
rect 10961 10375 10967 10401
rect 8247 10369 8273 10375
rect 13735 10369 13761 10375
rect 7463 10345 7489 10351
rect 7463 10313 7489 10319
rect 9815 10345 9841 10351
rect 13455 10345 13481 10351
rect 11881 10319 11887 10345
rect 11913 10319 11919 10345
rect 9815 10313 9841 10319
rect 13455 10313 13481 10319
rect 13847 10345 13873 10351
rect 13847 10313 13873 10319
rect 13903 10345 13929 10351
rect 13903 10313 13929 10319
rect 13623 10289 13649 10295
rect 8409 10263 8415 10289
rect 8441 10263 8447 10289
rect 13623 10257 13649 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 12839 10121 12865 10127
rect 10201 10095 10207 10121
rect 10233 10095 10239 10121
rect 10537 10095 10543 10121
rect 10569 10095 10575 10121
rect 12839 10089 12865 10095
rect 7967 10065 7993 10071
rect 7967 10033 7993 10039
rect 8079 10065 8105 10071
rect 9871 10065 9897 10071
rect 8969 10039 8975 10065
rect 9001 10039 9007 10065
rect 8079 10033 8105 10039
rect 9871 10033 9897 10039
rect 13287 10065 13313 10071
rect 13287 10033 13313 10039
rect 8023 10009 8049 10015
rect 8023 9977 8049 9983
rect 8135 10009 8161 10015
rect 8695 10009 8721 10015
rect 8241 9983 8247 10009
rect 8273 9983 8279 10009
rect 8135 9977 8161 9983
rect 8695 9977 8721 9983
rect 9143 10009 9169 10015
rect 9143 9977 9169 9983
rect 10039 10009 10065 10015
rect 10711 10009 10737 10015
rect 12727 10009 12753 10015
rect 10313 9983 10319 10009
rect 10345 9983 10351 10009
rect 10873 9983 10879 10009
rect 10905 9983 10911 10009
rect 10039 9977 10065 9983
rect 10711 9977 10737 9983
rect 12727 9977 12753 9983
rect 12839 10009 12865 10015
rect 12839 9977 12865 9983
rect 13007 10009 13033 10015
rect 13007 9977 13033 9983
rect 13175 10009 13201 10015
rect 13175 9977 13201 9983
rect 13511 10009 13537 10015
rect 13511 9977 13537 9983
rect 9423 9953 9449 9959
rect 13231 9953 13257 9959
rect 11265 9927 11271 9953
rect 11297 9927 11303 9953
rect 12329 9927 12335 9953
rect 12361 9927 12367 9953
rect 9423 9921 9449 9927
rect 13231 9921 13257 9927
rect 8807 9897 8833 9903
rect 8807 9865 8833 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 8303 9729 8329 9735
rect 8303 9697 8329 9703
rect 8471 9729 8497 9735
rect 9255 9729 9281 9735
rect 8969 9703 8975 9729
rect 9001 9703 9007 9729
rect 8471 9697 8497 9703
rect 9255 9697 9281 9703
rect 10935 9729 10961 9735
rect 10935 9697 10961 9703
rect 11215 9729 11241 9735
rect 12329 9703 12335 9729
rect 12361 9703 12367 9729
rect 11215 9697 11241 9703
rect 967 9673 993 9679
rect 967 9641 993 9647
rect 7687 9673 7713 9679
rect 7687 9641 7713 9647
rect 10655 9673 10681 9679
rect 10655 9641 10681 9647
rect 11159 9673 11185 9679
rect 11159 9641 11185 9647
rect 11607 9673 11633 9679
rect 20007 9673 20033 9679
rect 12441 9647 12447 9673
rect 12473 9647 12479 9673
rect 14289 9647 14295 9673
rect 14321 9647 14327 9673
rect 11607 9641 11633 9647
rect 20007 9641 20033 9647
rect 7183 9617 7209 9623
rect 2137 9591 2143 9617
rect 2169 9591 2175 9617
rect 7183 9585 7209 9591
rect 7239 9617 7265 9623
rect 8639 9617 8665 9623
rect 7457 9591 7463 9617
rect 7489 9591 7495 9617
rect 8073 9591 8079 9617
rect 8105 9591 8111 9617
rect 7239 9585 7265 9591
rect 8639 9585 8665 9591
rect 8863 9617 8889 9623
rect 9983 9617 10009 9623
rect 9305 9591 9311 9617
rect 9337 9591 9343 9617
rect 8863 9585 8889 9591
rect 9983 9585 10009 9591
rect 10039 9617 10065 9623
rect 10767 9617 10793 9623
rect 10257 9591 10263 9617
rect 10289 9591 10295 9617
rect 11657 9591 11663 9617
rect 11689 9591 11695 9617
rect 12161 9591 12167 9617
rect 12193 9591 12199 9617
rect 12833 9591 12839 9617
rect 12865 9591 12871 9617
rect 18825 9591 18831 9617
rect 18857 9591 18863 9617
rect 10039 9585 10065 9591
rect 10767 9585 10793 9591
rect 9703 9561 9729 9567
rect 9361 9535 9367 9561
rect 9393 9535 9399 9561
rect 9703 9529 9729 9535
rect 9759 9561 9785 9567
rect 9759 9529 9785 9535
rect 11439 9561 11465 9567
rect 13225 9535 13231 9561
rect 13257 9535 13263 9561
rect 11439 9529 11465 9535
rect 7295 9505 7321 9511
rect 7295 9473 7321 9479
rect 7351 9505 7377 9511
rect 8359 9505 8385 9511
rect 7961 9479 7967 9505
rect 7993 9479 7999 9505
rect 7351 9473 7377 9479
rect 8359 9473 8385 9479
rect 10095 9505 10121 9511
rect 10095 9473 10121 9479
rect 11551 9505 11577 9511
rect 11551 9473 11577 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 7799 9337 7825 9343
rect 7799 9305 7825 9311
rect 7911 9337 7937 9343
rect 7911 9305 7937 9311
rect 11831 9337 11857 9343
rect 11831 9305 11857 9311
rect 12671 9337 12697 9343
rect 12671 9305 12697 9311
rect 13343 9337 13369 9343
rect 13343 9305 13369 9311
rect 13735 9337 13761 9343
rect 13735 9305 13761 9311
rect 14127 9337 14153 9343
rect 14127 9305 14153 9311
rect 7631 9281 7657 9287
rect 7569 9255 7575 9281
rect 7601 9255 7607 9281
rect 7631 9249 7657 9255
rect 7687 9281 7713 9287
rect 7687 9249 7713 9255
rect 8023 9281 8049 9287
rect 8023 9249 8049 9255
rect 8079 9281 8105 9287
rect 8079 9249 8105 9255
rect 8415 9281 8441 9287
rect 12167 9281 12193 9287
rect 9753 9255 9759 9281
rect 9785 9255 9791 9281
rect 9977 9255 9983 9281
rect 10009 9255 10015 9281
rect 8415 9249 8441 9255
rect 12167 9249 12193 9255
rect 13287 9281 13313 9287
rect 13287 9249 13313 9255
rect 13623 9281 13649 9287
rect 13623 9249 13649 9255
rect 14071 9281 14097 9287
rect 14071 9249 14097 9255
rect 8247 9225 8273 9231
rect 9031 9225 9057 9231
rect 10487 9225 10513 9231
rect 6673 9199 6679 9225
rect 6705 9199 6711 9225
rect 7065 9199 7071 9225
rect 7097 9199 7103 9225
rect 8801 9199 8807 9225
rect 8833 9199 8839 9225
rect 9249 9199 9255 9225
rect 9281 9199 9287 9225
rect 9585 9199 9591 9225
rect 9617 9199 9623 9225
rect 8247 9193 8273 9199
rect 9031 9193 9057 9199
rect 10487 9193 10513 9199
rect 10711 9225 10737 9231
rect 10711 9193 10737 9199
rect 11775 9225 11801 9231
rect 11775 9193 11801 9199
rect 11943 9225 11969 9231
rect 11943 9193 11969 9199
rect 13175 9225 13201 9231
rect 13175 9193 13201 9199
rect 13455 9225 13481 9231
rect 13455 9193 13481 9199
rect 13679 9225 13705 9231
rect 13679 9193 13705 9199
rect 13959 9225 13985 9231
rect 13959 9193 13985 9199
rect 5609 9143 5615 9169
rect 5641 9143 5647 9169
rect 7401 9143 7407 9169
rect 7433 9143 7439 9169
rect 9641 9143 9647 9169
rect 9673 9143 9679 9169
rect 10767 9113 10793 9119
rect 10033 9087 10039 9113
rect 10065 9087 10071 9113
rect 10767 9081 10793 9087
rect 12111 9113 12137 9119
rect 12111 9081 12137 9087
rect 14127 9113 14153 9119
rect 14127 9081 14153 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 7183 8945 7209 8951
rect 7183 8913 7209 8919
rect 9031 8945 9057 8951
rect 9031 8913 9057 8919
rect 7463 8889 7489 8895
rect 7463 8857 7489 8863
rect 7967 8889 7993 8895
rect 7967 8857 7993 8863
rect 8919 8889 8945 8895
rect 13511 8889 13537 8895
rect 10313 8863 10319 8889
rect 10345 8863 10351 8889
rect 11097 8863 11103 8889
rect 11129 8863 11135 8889
rect 8919 8857 8945 8863
rect 13511 8857 13537 8863
rect 20007 8889 20033 8895
rect 20007 8857 20033 8863
rect 7239 8833 7265 8839
rect 9367 8833 9393 8839
rect 10263 8833 10289 8839
rect 8353 8807 8359 8833
rect 8385 8807 8391 8833
rect 9809 8807 9815 8833
rect 9841 8807 9847 8833
rect 10033 8807 10039 8833
rect 10065 8807 10071 8833
rect 12553 8807 12559 8833
rect 12585 8807 12591 8833
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 7239 8801 7265 8807
rect 9367 8801 9393 8807
rect 10263 8801 10289 8807
rect 7183 8777 7209 8783
rect 8241 8751 8247 8777
rect 8273 8751 8279 8777
rect 9529 8751 9535 8777
rect 9561 8751 9567 8777
rect 12161 8751 12167 8777
rect 12193 8751 12199 8777
rect 7183 8745 7209 8751
rect 10151 8721 10177 8727
rect 9193 8695 9199 8721
rect 9225 8695 9231 8721
rect 9697 8695 9703 8721
rect 9729 8695 9735 8721
rect 10151 8689 10177 8695
rect 10319 8721 10345 8727
rect 10319 8689 10345 8695
rect 10935 8721 10961 8727
rect 10935 8689 10961 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 7239 8553 7265 8559
rect 7239 8521 7265 8527
rect 13119 8553 13145 8559
rect 13119 8521 13145 8527
rect 7631 8497 7657 8503
rect 7631 8465 7657 8471
rect 7743 8497 7769 8503
rect 10929 8471 10935 8497
rect 10961 8471 10967 8497
rect 13673 8471 13679 8497
rect 13705 8471 13711 8497
rect 7743 8465 7769 8471
rect 7127 8441 7153 8447
rect 2137 8415 2143 8441
rect 2169 8415 2175 8441
rect 7127 8409 7153 8415
rect 7463 8441 7489 8447
rect 11881 8415 11887 8441
rect 11913 8415 11919 8441
rect 13281 8415 13287 8441
rect 13313 8415 13319 8441
rect 7463 8409 7489 8415
rect 7183 8385 7209 8391
rect 7569 8359 7575 8385
rect 7601 8359 7607 8385
rect 14737 8359 14743 8385
rect 14769 8359 14775 8385
rect 7183 8353 7209 8359
rect 967 8329 993 8335
rect 967 8297 993 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 12391 8161 12417 8167
rect 10929 8135 10935 8161
rect 10961 8135 10967 8161
rect 12391 8129 12417 8135
rect 12503 8105 12529 8111
rect 12503 8073 12529 8079
rect 9199 8049 9225 8055
rect 9199 8017 9225 8023
rect 10655 8049 10681 8055
rect 10655 8017 10681 8023
rect 10823 8049 10849 8055
rect 11327 8049 11353 8055
rect 11041 8023 11047 8049
rect 11073 8023 11079 8049
rect 10823 8017 10849 8023
rect 11327 8017 11353 8023
rect 13287 8049 13313 8055
rect 13287 8017 13313 8023
rect 9143 7993 9169 7999
rect 9143 7961 9169 7967
rect 11215 7993 11241 7999
rect 11215 7961 11241 7967
rect 11495 7993 11521 7999
rect 11495 7961 11521 7967
rect 9031 7937 9057 7943
rect 9031 7905 9057 7911
rect 10711 7937 10737 7943
rect 10711 7905 10737 7911
rect 11271 7937 11297 7943
rect 12217 7911 12223 7937
rect 12249 7911 12255 7937
rect 13113 7911 13119 7937
rect 13145 7911 13151 7937
rect 11271 7905 11297 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 8695 7769 8721 7775
rect 8695 7737 8721 7743
rect 8807 7769 8833 7775
rect 8807 7737 8833 7743
rect 11439 7769 11465 7775
rect 11439 7737 11465 7743
rect 12671 7769 12697 7775
rect 12671 7737 12697 7743
rect 13343 7769 13369 7775
rect 13343 7737 13369 7743
rect 13623 7769 13649 7775
rect 13623 7737 13649 7743
rect 7631 7713 7657 7719
rect 13567 7713 13593 7719
rect 7009 7687 7015 7713
rect 7041 7687 7047 7713
rect 10145 7687 10151 7713
rect 10177 7687 10183 7713
rect 7631 7681 7657 7687
rect 13567 7681 13593 7687
rect 9031 7657 9057 7663
rect 13231 7657 13257 7663
rect 7401 7631 7407 7657
rect 7433 7631 7439 7657
rect 8017 7631 8023 7657
rect 8049 7631 8055 7657
rect 9753 7631 9759 7657
rect 9785 7631 9791 7657
rect 9031 7625 9057 7631
rect 13231 7625 13257 7631
rect 13399 7657 13425 7663
rect 13399 7625 13425 7631
rect 13735 7657 13761 7663
rect 18825 7631 18831 7657
rect 18857 7631 18863 7657
rect 13735 7625 13761 7631
rect 7855 7601 7881 7607
rect 5945 7575 5951 7601
rect 5977 7575 5983 7601
rect 7855 7569 7881 7575
rect 7911 7601 7937 7607
rect 7911 7569 7937 7575
rect 8751 7601 8777 7607
rect 13063 7601 13089 7607
rect 11209 7575 11215 7601
rect 11241 7575 11247 7601
rect 8751 7569 8777 7575
rect 13063 7569 13089 7575
rect 13119 7601 13145 7607
rect 13119 7569 13145 7575
rect 20007 7601 20033 7607
rect 20007 7569 20033 7575
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 7463 7377 7489 7383
rect 7463 7345 7489 7351
rect 7631 7377 7657 7383
rect 7631 7345 7657 7351
rect 7793 7295 7799 7321
rect 7825 7295 7831 7321
rect 8857 7295 8863 7321
rect 8889 7295 8895 7321
rect 13225 7295 13231 7321
rect 13257 7295 13263 7321
rect 14289 7295 14295 7321
rect 14321 7295 14327 7321
rect 9479 7265 9505 7271
rect 9249 7239 9255 7265
rect 9281 7239 9287 7265
rect 9479 7233 9505 7239
rect 10263 7265 10289 7271
rect 10767 7265 10793 7271
rect 10649 7239 10655 7265
rect 10681 7239 10687 7265
rect 10263 7233 10289 7239
rect 10767 7233 10793 7239
rect 10935 7265 10961 7271
rect 12447 7265 12473 7271
rect 12329 7239 12335 7265
rect 12361 7239 12367 7265
rect 10935 7233 10961 7239
rect 12447 7233 12473 7239
rect 12559 7265 12585 7271
rect 12559 7233 12585 7239
rect 12615 7265 12641 7271
rect 12833 7239 12839 7265
rect 12865 7239 12871 7265
rect 12615 7233 12641 7239
rect 11215 7209 11241 7215
rect 11215 7177 11241 7183
rect 7519 7153 7545 7159
rect 7519 7121 7545 7127
rect 10095 7153 10121 7159
rect 10095 7121 10121 7127
rect 10207 7153 10233 7159
rect 10207 7121 10233 7127
rect 10823 7153 10849 7159
rect 10823 7121 10849 7127
rect 10879 7153 10905 7159
rect 10879 7121 10905 7127
rect 11159 7153 11185 7159
rect 11159 7121 11185 7127
rect 12503 7153 12529 7159
rect 12503 7121 12529 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 8359 6985 8385 6991
rect 8359 6953 8385 6959
rect 9367 6985 9393 6991
rect 9367 6953 9393 6959
rect 11831 6985 11857 6991
rect 11831 6953 11857 6959
rect 12335 6985 12361 6991
rect 12335 6953 12361 6959
rect 9423 6929 9449 6935
rect 7737 6903 7743 6929
rect 7769 6903 7775 6929
rect 10537 6903 10543 6929
rect 10569 6903 10575 6929
rect 13001 6903 13007 6929
rect 13033 6903 13039 6929
rect 9423 6897 9449 6903
rect 9255 6873 9281 6879
rect 8073 6847 8079 6873
rect 8105 6847 8111 6873
rect 10201 6847 10207 6873
rect 10233 6847 10239 6873
rect 12665 6847 12671 6873
rect 12697 6847 12703 6873
rect 9255 6841 9281 6847
rect 6673 6791 6679 6817
rect 6705 6791 6711 6817
rect 11601 6791 11607 6817
rect 11633 6791 11639 6817
rect 14065 6791 14071 6817
rect 14097 6791 14103 6817
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 10767 6537 10793 6543
rect 9249 6511 9255 6537
rect 9281 6511 9287 6537
rect 10313 6511 10319 6537
rect 10345 6511 10351 6537
rect 10767 6505 10793 6511
rect 8857 6455 8863 6481
rect 8889 6455 8895 6481
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 10537 2143 10543 2169
rect 10569 2143 10575 2169
rect 14289 2143 14295 2169
rect 14321 2143 14327 2169
rect 11047 2057 11073 2063
rect 11047 2025 11073 2031
rect 13343 2057 13369 2063
rect 13343 2025 13369 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 10823 1833 10849 1839
rect 10823 1801 10849 1807
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 8465 1751 8471 1777
rect 8497 1751 8503 1777
rect 11769 1751 11775 1777
rect 11801 1751 11807 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 9249 1695 9255 1721
rect 9281 1695 9287 1721
rect 7183 1665 7209 1671
rect 7183 1633 7209 1639
rect 14239 1665 14265 1671
rect 14239 1633 14265 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9031 19111 9057 19137
rect 11215 19111 11241 19137
rect 12783 19111 12809 19137
rect 8527 18999 8553 19025
rect 10879 18999 10905 19025
rect 12391 18999 12417 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 9927 18719 9953 18745
rect 11383 18719 11409 18745
rect 9423 18607 9449 18633
rect 10991 18607 11017 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 7967 13847 7993 13873
rect 9311 13847 9337 13873
rect 7911 13791 7937 13817
rect 9255 13791 9281 13817
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 967 13567 993 13593
rect 7351 13567 7377 13593
rect 8415 13567 8441 13593
rect 8975 13567 9001 13593
rect 10039 13567 10065 13593
rect 2143 13511 2169 13537
rect 7015 13511 7041 13537
rect 8639 13511 8665 13537
rect 10991 13511 11017 13537
rect 10263 13455 10289 13481
rect 10879 13455 10905 13481
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 8247 13231 8273 13257
rect 8303 13231 8329 13257
rect 9255 13231 9281 13257
rect 9311 13231 9337 13257
rect 13063 13175 13089 13201
rect 2143 13119 2169 13145
rect 7239 13119 7265 13145
rect 7463 13119 7489 13145
rect 8135 13119 8161 13145
rect 8191 13119 8217 13145
rect 8415 13119 8441 13145
rect 9143 13119 9169 13145
rect 9199 13119 9225 13145
rect 9367 13119 9393 13145
rect 9591 13119 9617 13145
rect 13119 13119 13145 13145
rect 18831 13119 18857 13145
rect 5783 13063 5809 13089
rect 6847 13063 6873 13089
rect 8751 13063 8777 13089
rect 9983 13063 10009 13089
rect 11047 13063 11073 13089
rect 11271 13063 11297 13089
rect 11495 13063 11521 13089
rect 12671 13063 12697 13089
rect 13343 13063 13369 13089
rect 967 13007 993 13033
rect 13063 13007 13089 13033
rect 20007 13007 20033 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 9815 12783 9841 12809
rect 10039 12783 10065 12809
rect 12391 12783 12417 12809
rect 14015 12783 14041 12809
rect 6903 12727 6929 12753
rect 7183 12727 7209 12753
rect 7351 12727 7377 12753
rect 7519 12727 7545 12753
rect 9983 12727 10009 12753
rect 10319 12727 10345 12753
rect 10599 12727 10625 12753
rect 10935 12727 10961 12753
rect 12615 12727 12641 12753
rect 7015 12671 7041 12697
rect 7071 12671 7097 12697
rect 7295 12671 7321 12697
rect 9647 12671 9673 12697
rect 10711 12671 10737 12697
rect 10767 12671 10793 12697
rect 11327 12671 11353 12697
rect 12951 12671 12977 12697
rect 7575 12615 7601 12641
rect 7687 12615 7713 12641
rect 9759 12615 9785 12641
rect 10095 12615 10121 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 9311 12447 9337 12473
rect 11271 12447 11297 12473
rect 11775 12447 11801 12473
rect 12671 12447 12697 12473
rect 10319 12391 10345 12417
rect 11439 12391 11465 12417
rect 11943 12391 11969 12417
rect 7463 12335 7489 12361
rect 7687 12335 7713 12361
rect 7855 12335 7881 12361
rect 7967 12335 7993 12361
rect 9423 12335 9449 12361
rect 11103 12335 11129 12361
rect 11271 12335 11297 12361
rect 11663 12335 11689 12361
rect 11719 12335 11745 12361
rect 11831 12335 11857 12361
rect 12839 12335 12865 12361
rect 18831 12335 18857 12361
rect 6063 12279 6089 12305
rect 7127 12279 7153 12305
rect 7911 12279 7937 12305
rect 8191 12279 8217 12305
rect 10207 12279 10233 12305
rect 10375 12279 10401 12305
rect 10879 12279 10905 12305
rect 13231 12279 13257 12305
rect 14295 12279 14321 12305
rect 20007 12223 20033 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 11215 12055 11241 12081
rect 12895 11999 12921 12025
rect 20007 11999 20033 12025
rect 8807 11943 8833 11969
rect 9479 11943 9505 11969
rect 9591 11943 9617 11969
rect 9983 11943 10009 11969
rect 10095 11943 10121 11969
rect 10991 11943 11017 11969
rect 11551 11943 11577 11969
rect 12727 11943 12753 11969
rect 12951 11943 12977 11969
rect 13063 11943 13089 11969
rect 13399 11943 13425 11969
rect 13623 11943 13649 11969
rect 13735 11943 13761 11969
rect 14071 11943 14097 11969
rect 18831 11943 18857 11969
rect 9647 11887 9673 11913
rect 10375 11887 10401 11913
rect 11271 11887 11297 11913
rect 12615 11887 12641 11913
rect 12839 11887 12865 11913
rect 13287 11887 13313 11913
rect 13567 11887 13593 11913
rect 13847 11887 13873 11913
rect 14183 11887 14209 11913
rect 7631 11831 7657 11857
rect 8695 11831 8721 11857
rect 9815 11831 9841 11857
rect 10207 11831 10233 11857
rect 10319 11831 10345 11857
rect 11439 11831 11465 11857
rect 13231 11831 13257 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 13399 11663 13425 11689
rect 7183 11607 7209 11633
rect 9087 11607 9113 11633
rect 9311 11607 9337 11633
rect 7575 11551 7601 11577
rect 7687 11551 7713 11577
rect 7743 11551 7769 11577
rect 7799 11551 7825 11577
rect 7911 11551 7937 11577
rect 9367 11551 9393 11577
rect 11887 11551 11913 11577
rect 8303 11495 8329 11521
rect 8751 11495 8777 11521
rect 10095 11495 10121 11521
rect 7127 11439 7153 11465
rect 7295 11439 7321 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 8863 11271 8889 11297
rect 967 11215 993 11241
rect 8191 11215 8217 11241
rect 8415 11215 8441 11241
rect 12615 11215 12641 11241
rect 13343 11215 13369 11241
rect 2143 11159 2169 11185
rect 6791 11159 6817 11185
rect 8359 11159 8385 11185
rect 8639 11159 8665 11185
rect 9087 11159 9113 11185
rect 9311 11159 9337 11185
rect 9703 11159 9729 11185
rect 9927 11159 9953 11185
rect 9983 11159 10009 11185
rect 10823 11159 10849 11185
rect 11047 11159 11073 11185
rect 12895 11159 12921 11185
rect 13007 11159 13033 11185
rect 7127 11103 7153 11129
rect 8807 11103 8833 11129
rect 10207 11103 10233 11129
rect 10655 11103 10681 11129
rect 11383 11103 11409 11129
rect 8471 11047 8497 11073
rect 10263 11047 10289 11073
rect 11215 11047 11241 11073
rect 11551 11047 11577 11073
rect 11719 11047 11745 11073
rect 12615 11047 12641 11073
rect 12727 11047 12753 11073
rect 13063 11047 13089 11073
rect 13175 11047 13201 11073
rect 20119 11047 20145 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 8023 10879 8049 10905
rect 8079 10879 8105 10905
rect 9087 10879 9113 10905
rect 6679 10823 6705 10849
rect 7911 10823 7937 10849
rect 8919 10823 8945 10849
rect 10431 10823 10457 10849
rect 10823 10823 10849 10849
rect 13063 10823 13089 10849
rect 2143 10767 2169 10793
rect 7015 10767 7041 10793
rect 7239 10767 7265 10793
rect 7351 10767 7377 10793
rect 7463 10767 7489 10793
rect 7575 10767 7601 10793
rect 7743 10767 7769 10793
rect 8135 10767 8161 10793
rect 9871 10767 9897 10793
rect 10655 10767 10681 10793
rect 10879 10767 10905 10793
rect 11719 10767 11745 10793
rect 12727 10767 12753 10793
rect 12839 10767 12865 10793
rect 12951 10767 12977 10793
rect 13287 10767 13313 10793
rect 18831 10767 18857 10793
rect 5615 10711 5641 10737
rect 7295 10711 7321 10737
rect 9591 10711 9617 10737
rect 13623 10711 13649 10737
rect 14687 10711 14713 10737
rect 967 10655 993 10681
rect 13007 10655 13033 10681
rect 20007 10655 20033 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 7015 10487 7041 10513
rect 7463 10487 7489 10513
rect 9927 10487 9953 10513
rect 4999 10431 5025 10457
rect 6063 10431 6089 10457
rect 6791 10431 6817 10457
rect 6959 10431 6985 10457
rect 9871 10431 9897 10457
rect 10151 10431 10177 10457
rect 6455 10375 6481 10401
rect 7239 10375 7265 10401
rect 7519 10375 7545 10401
rect 8247 10375 8273 10401
rect 10319 10375 10345 10401
rect 10935 10375 10961 10401
rect 13735 10375 13761 10401
rect 7463 10319 7489 10345
rect 9815 10319 9841 10345
rect 11887 10319 11913 10345
rect 13455 10319 13481 10345
rect 13847 10319 13873 10345
rect 13903 10319 13929 10345
rect 8415 10263 8441 10289
rect 13623 10263 13649 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 10207 10095 10233 10121
rect 10543 10095 10569 10121
rect 12839 10095 12865 10121
rect 7967 10039 7993 10065
rect 8079 10039 8105 10065
rect 8975 10039 9001 10065
rect 9871 10039 9897 10065
rect 13287 10039 13313 10065
rect 8023 9983 8049 10009
rect 8135 9983 8161 10009
rect 8247 9983 8273 10009
rect 8695 9983 8721 10009
rect 9143 9983 9169 10009
rect 10039 9983 10065 10009
rect 10319 9983 10345 10009
rect 10711 9983 10737 10009
rect 10879 9983 10905 10009
rect 12727 9983 12753 10009
rect 12839 9983 12865 10009
rect 13007 9983 13033 10009
rect 13175 9983 13201 10009
rect 13511 9983 13537 10009
rect 9423 9927 9449 9953
rect 11271 9927 11297 9953
rect 12335 9927 12361 9953
rect 13231 9927 13257 9953
rect 8807 9871 8833 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 8303 9703 8329 9729
rect 8471 9703 8497 9729
rect 8975 9703 9001 9729
rect 9255 9703 9281 9729
rect 10935 9703 10961 9729
rect 11215 9703 11241 9729
rect 12335 9703 12361 9729
rect 967 9647 993 9673
rect 7687 9647 7713 9673
rect 10655 9647 10681 9673
rect 11159 9647 11185 9673
rect 11607 9647 11633 9673
rect 12447 9647 12473 9673
rect 14295 9647 14321 9673
rect 20007 9647 20033 9673
rect 2143 9591 2169 9617
rect 7183 9591 7209 9617
rect 7239 9591 7265 9617
rect 7463 9591 7489 9617
rect 8079 9591 8105 9617
rect 8639 9591 8665 9617
rect 8863 9591 8889 9617
rect 9311 9591 9337 9617
rect 9983 9591 10009 9617
rect 10039 9591 10065 9617
rect 10263 9591 10289 9617
rect 10767 9591 10793 9617
rect 11663 9591 11689 9617
rect 12167 9591 12193 9617
rect 12839 9591 12865 9617
rect 18831 9591 18857 9617
rect 9367 9535 9393 9561
rect 9703 9535 9729 9561
rect 9759 9535 9785 9561
rect 11439 9535 11465 9561
rect 13231 9535 13257 9561
rect 7295 9479 7321 9505
rect 7351 9479 7377 9505
rect 7967 9479 7993 9505
rect 8359 9479 8385 9505
rect 10095 9479 10121 9505
rect 11551 9479 11577 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 7799 9311 7825 9337
rect 7911 9311 7937 9337
rect 11831 9311 11857 9337
rect 12671 9311 12697 9337
rect 13343 9311 13369 9337
rect 13735 9311 13761 9337
rect 14127 9311 14153 9337
rect 7575 9255 7601 9281
rect 7631 9255 7657 9281
rect 7687 9255 7713 9281
rect 8023 9255 8049 9281
rect 8079 9255 8105 9281
rect 8415 9255 8441 9281
rect 9759 9255 9785 9281
rect 9983 9255 10009 9281
rect 12167 9255 12193 9281
rect 13287 9255 13313 9281
rect 13623 9255 13649 9281
rect 14071 9255 14097 9281
rect 6679 9199 6705 9225
rect 7071 9199 7097 9225
rect 8247 9199 8273 9225
rect 8807 9199 8833 9225
rect 9031 9199 9057 9225
rect 9255 9199 9281 9225
rect 9591 9199 9617 9225
rect 10487 9199 10513 9225
rect 10711 9199 10737 9225
rect 11775 9199 11801 9225
rect 11943 9199 11969 9225
rect 13175 9199 13201 9225
rect 13455 9199 13481 9225
rect 13679 9199 13705 9225
rect 13959 9199 13985 9225
rect 5615 9143 5641 9169
rect 7407 9143 7433 9169
rect 9647 9143 9673 9169
rect 10039 9087 10065 9113
rect 10767 9087 10793 9113
rect 12111 9087 12137 9113
rect 14127 9087 14153 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 7183 8919 7209 8945
rect 9031 8919 9057 8945
rect 7463 8863 7489 8889
rect 7967 8863 7993 8889
rect 8919 8863 8945 8889
rect 10319 8863 10345 8889
rect 11103 8863 11129 8889
rect 13511 8863 13537 8889
rect 20007 8863 20033 8889
rect 7239 8807 7265 8833
rect 8359 8807 8385 8833
rect 9367 8807 9393 8833
rect 9815 8807 9841 8833
rect 10039 8807 10065 8833
rect 10263 8807 10289 8833
rect 12559 8807 12585 8833
rect 18831 8807 18857 8833
rect 7183 8751 7209 8777
rect 8247 8751 8273 8777
rect 9535 8751 9561 8777
rect 12167 8751 12193 8777
rect 9199 8695 9225 8721
rect 9703 8695 9729 8721
rect 10151 8695 10177 8721
rect 10319 8695 10345 8721
rect 10935 8695 10961 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7239 8527 7265 8553
rect 13119 8527 13145 8553
rect 7631 8471 7657 8497
rect 7743 8471 7769 8497
rect 10935 8471 10961 8497
rect 13679 8471 13705 8497
rect 2143 8415 2169 8441
rect 7127 8415 7153 8441
rect 7463 8415 7489 8441
rect 11887 8415 11913 8441
rect 13287 8415 13313 8441
rect 7183 8359 7209 8385
rect 7575 8359 7601 8385
rect 14743 8359 14769 8385
rect 967 8303 993 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 10935 8135 10961 8161
rect 12391 8135 12417 8161
rect 12503 8079 12529 8105
rect 9199 8023 9225 8049
rect 10655 8023 10681 8049
rect 10823 8023 10849 8049
rect 11047 8023 11073 8049
rect 11327 8023 11353 8049
rect 13287 8023 13313 8049
rect 9143 7967 9169 7993
rect 11215 7967 11241 7993
rect 11495 7967 11521 7993
rect 9031 7911 9057 7937
rect 10711 7911 10737 7937
rect 11271 7911 11297 7937
rect 12223 7911 12249 7937
rect 13119 7911 13145 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 8695 7743 8721 7769
rect 8807 7743 8833 7769
rect 11439 7743 11465 7769
rect 12671 7743 12697 7769
rect 13343 7743 13369 7769
rect 13623 7743 13649 7769
rect 7015 7687 7041 7713
rect 7631 7687 7657 7713
rect 10151 7687 10177 7713
rect 13567 7687 13593 7713
rect 7407 7631 7433 7657
rect 8023 7631 8049 7657
rect 9031 7631 9057 7657
rect 9759 7631 9785 7657
rect 13231 7631 13257 7657
rect 13399 7631 13425 7657
rect 13735 7631 13761 7657
rect 18831 7631 18857 7657
rect 5951 7575 5977 7601
rect 7855 7575 7881 7601
rect 7911 7575 7937 7601
rect 8751 7575 8777 7601
rect 11215 7575 11241 7601
rect 13063 7575 13089 7601
rect 13119 7575 13145 7601
rect 20007 7575 20033 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 7463 7351 7489 7377
rect 7631 7351 7657 7377
rect 7799 7295 7825 7321
rect 8863 7295 8889 7321
rect 13231 7295 13257 7321
rect 14295 7295 14321 7321
rect 9255 7239 9281 7265
rect 9479 7239 9505 7265
rect 10263 7239 10289 7265
rect 10655 7239 10681 7265
rect 10767 7239 10793 7265
rect 10935 7239 10961 7265
rect 12335 7239 12361 7265
rect 12447 7239 12473 7265
rect 12559 7239 12585 7265
rect 12615 7239 12641 7265
rect 12839 7239 12865 7265
rect 11215 7183 11241 7209
rect 7519 7127 7545 7153
rect 10095 7127 10121 7153
rect 10207 7127 10233 7153
rect 10823 7127 10849 7153
rect 10879 7127 10905 7153
rect 11159 7127 11185 7153
rect 12503 7127 12529 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 8359 6959 8385 6985
rect 9367 6959 9393 6985
rect 11831 6959 11857 6985
rect 12335 6959 12361 6985
rect 7743 6903 7769 6929
rect 9423 6903 9449 6929
rect 10543 6903 10569 6929
rect 13007 6903 13033 6929
rect 8079 6847 8105 6873
rect 9255 6847 9281 6873
rect 10207 6847 10233 6873
rect 12671 6847 12697 6873
rect 6679 6791 6705 6817
rect 11607 6791 11633 6817
rect 14071 6791 14097 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9255 6511 9281 6537
rect 10319 6511 10345 6537
rect 10767 6511 10793 6537
rect 8863 6455 8889 6481
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 10543 2143 10569 2169
rect 14295 2143 14321 2169
rect 11047 2031 11073 2057
rect 13343 2031 13369 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 10823 1807 10849 1833
rect 12783 1807 12809 1833
rect 8471 1751 8497 1777
rect 11775 1751 11801 1777
rect 12279 1751 12305 1777
rect 9255 1695 9281 1721
rect 7183 1639 7209 1665
rect 14239 1639 14265 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8400 20600 8456 21000
rect 9744 20600 9800 21000
rect 10752 20600 10808 21000
rect 11088 20600 11144 21000
rect 12096 20600 12152 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 8414 19138 8442 20600
rect 8414 19105 8442 19110
rect 9030 19138 9058 19143
rect 9030 19091 9058 19110
rect 8526 19025 8554 19031
rect 8526 18999 8527 19025
rect 8553 18999 8554 19025
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 8526 15974 8554 18999
rect 9758 18802 9786 20600
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9758 18774 9842 18802
rect 9918 18797 10050 18802
rect 9814 18746 9842 18774
rect 9926 18746 9954 18751
rect 9814 18745 9954 18746
rect 9814 18719 9927 18745
rect 9953 18719 9954 18745
rect 9814 18718 9954 18719
rect 9926 18713 9954 18718
rect 10766 18746 10794 20600
rect 11102 19138 11130 20600
rect 11214 19138 11242 19143
rect 11102 19137 11242 19138
rect 11102 19111 11215 19137
rect 11241 19111 11242 19137
rect 11102 19110 11242 19111
rect 11214 19105 11242 19110
rect 12110 19138 12138 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 12110 19105 12138 19110
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 10766 18713 10794 18718
rect 10878 19025 10906 19031
rect 10878 18999 10879 19025
rect 10905 18999 10906 19025
rect 8414 15946 8554 15974
rect 9422 18633 9450 18639
rect 9422 18607 9423 18633
rect 9449 18607 9450 18633
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 7966 13874 7994 13879
rect 7966 13873 8274 13874
rect 7966 13847 7967 13873
rect 7993 13847 8274 13873
rect 7966 13846 8274 13847
rect 7966 13841 7994 13846
rect 7350 13818 7378 13823
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 966 13593 994 13599
rect 966 13567 967 13593
rect 993 13567 994 13593
rect 966 13146 994 13567
rect 7350 13593 7378 13790
rect 7910 13818 7938 13823
rect 7910 13771 7938 13790
rect 7350 13567 7351 13593
rect 7377 13567 7378 13593
rect 7350 13561 7378 13567
rect 2142 13537 2170 13543
rect 2142 13511 2143 13537
rect 2169 13511 2170 13537
rect 966 13113 994 13118
rect 2086 13482 2114 13487
rect 966 13033 994 13039
rect 966 13007 967 13033
rect 993 13007 994 13033
rect 966 12810 994 13007
rect 966 12777 994 12782
rect 966 11242 994 11247
rect 966 11195 994 11214
rect 966 10681 994 10687
rect 966 10655 967 10681
rect 993 10655 994 10681
rect 966 10458 994 10655
rect 2086 10514 2114 13454
rect 2142 13258 2170 13511
rect 7014 13537 7042 13543
rect 7014 13511 7015 13537
rect 7041 13511 7042 13537
rect 2142 13225 2170 13230
rect 5782 13258 5810 13263
rect 2142 13146 2170 13151
rect 2142 13099 2170 13118
rect 5782 13089 5810 13230
rect 5782 13063 5783 13089
rect 5809 13063 5810 13089
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 5782 12698 5810 13063
rect 5782 12665 5810 12670
rect 6062 13146 6090 13151
rect 7014 13146 7042 13511
rect 8246 13257 8274 13846
rect 8414 13593 8442 15946
rect 9310 13873 9338 13879
rect 9310 13847 9311 13873
rect 9337 13847 9338 13873
rect 9254 13818 9282 13823
rect 8414 13567 8415 13593
rect 8441 13567 8442 13593
rect 8414 13454 8442 13567
rect 8974 13817 9282 13818
rect 8974 13791 9255 13817
rect 9281 13791 9282 13817
rect 8974 13790 9282 13791
rect 8974 13593 9002 13790
rect 9254 13785 9282 13790
rect 8974 13567 8975 13593
rect 9001 13567 9002 13593
rect 8974 13561 9002 13567
rect 8246 13231 8247 13257
rect 8273 13231 8274 13257
rect 8246 13225 8274 13231
rect 8302 13426 8442 13454
rect 8638 13537 8666 13543
rect 8638 13511 8639 13537
rect 8665 13511 8666 13537
rect 8638 13454 8666 13511
rect 9310 13454 9338 13847
rect 9422 13594 9450 18607
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 10038 13594 10066 13599
rect 9422 13593 10066 13594
rect 9422 13567 10039 13593
rect 10065 13567 10066 13593
rect 9422 13566 10066 13567
rect 9422 13454 9450 13566
rect 10038 13561 10066 13566
rect 8638 13426 8778 13454
rect 8302 13257 8330 13426
rect 8302 13231 8303 13257
rect 8329 13231 8330 13257
rect 8302 13225 8330 13231
rect 7238 13146 7266 13151
rect 7462 13146 7490 13151
rect 7014 13145 7490 13146
rect 7014 13119 7239 13145
rect 7265 13119 7463 13145
rect 7489 13119 7490 13145
rect 7014 13118 7490 13119
rect 6062 12642 6090 13118
rect 7238 13113 7266 13118
rect 6846 13090 6874 13095
rect 7462 13090 7490 13118
rect 8134 13145 8162 13151
rect 8134 13119 8135 13145
rect 8161 13119 8162 13145
rect 7518 13090 7546 13095
rect 6846 13089 6930 13090
rect 6846 13063 6847 13089
rect 6873 13063 6930 13089
rect 6846 13062 6930 13063
rect 6846 13057 6874 13062
rect 6902 12753 6930 13062
rect 7462 13062 7518 13090
rect 6902 12727 6903 12753
rect 6929 12727 6930 12753
rect 6902 12721 6930 12727
rect 7014 12782 7154 12810
rect 7014 12697 7042 12782
rect 7126 12754 7154 12782
rect 7182 12754 7210 12759
rect 7126 12753 7210 12754
rect 7126 12727 7183 12753
rect 7209 12727 7210 12753
rect 7126 12726 7210 12727
rect 7182 12721 7210 12726
rect 7350 12754 7378 12759
rect 7350 12707 7378 12726
rect 7014 12671 7015 12697
rect 7041 12671 7042 12697
rect 7014 12665 7042 12671
rect 7070 12697 7098 12703
rect 7070 12671 7071 12697
rect 7097 12671 7098 12697
rect 6062 12305 6090 12614
rect 6062 12279 6063 12305
rect 6089 12279 6090 12305
rect 6062 12273 6090 12279
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 6790 11690 6818 11695
rect 6678 11466 6706 11471
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 2142 11186 2170 11191
rect 2142 11139 2170 11158
rect 5614 11186 5642 11191
rect 2142 10794 2170 10799
rect 2142 10747 2170 10766
rect 4998 10794 5026 10799
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 2086 10481 2114 10486
rect 966 10425 994 10430
rect 4998 10458 5026 10766
rect 5614 10737 5642 11158
rect 6678 10849 6706 11438
rect 6678 10823 6679 10849
rect 6705 10823 6706 10849
rect 6678 10817 6706 10823
rect 6790 11186 6818 11662
rect 6790 11185 7042 11186
rect 6790 11159 6791 11185
rect 6817 11159 7042 11185
rect 6790 11158 7042 11159
rect 5614 10711 5615 10737
rect 5641 10711 5642 10737
rect 5614 10705 5642 10711
rect 6062 10738 6090 10743
rect 4998 10411 5026 10430
rect 6062 10457 6090 10710
rect 6062 10431 6063 10457
rect 6089 10431 6090 10457
rect 6062 10425 6090 10431
rect 6790 10457 6818 11158
rect 7014 10793 7042 11158
rect 7070 10850 7098 12671
rect 7294 12698 7322 12703
rect 7294 12651 7322 12670
rect 7462 12362 7490 13062
rect 7518 13057 7546 13062
rect 8134 12810 8162 13119
rect 8134 12777 8162 12782
rect 8190 13145 8218 13151
rect 8190 13119 8191 13145
rect 8217 13119 8218 13145
rect 7518 12754 7546 12759
rect 7518 12707 7546 12726
rect 7798 12698 7826 12703
rect 7574 12642 7602 12647
rect 7574 12595 7602 12614
rect 7686 12641 7714 12647
rect 7686 12615 7687 12641
rect 7713 12615 7714 12641
rect 7462 12361 7658 12362
rect 7462 12335 7463 12361
rect 7489 12335 7658 12361
rect 7462 12334 7658 12335
rect 7462 12329 7490 12334
rect 7126 12306 7154 12311
rect 7126 12259 7154 12278
rect 7630 11857 7658 12334
rect 7686 12361 7714 12615
rect 7686 12335 7687 12361
rect 7713 12335 7714 12361
rect 7686 12329 7714 12335
rect 7630 11831 7631 11857
rect 7657 11831 7658 11857
rect 7630 11690 7658 11831
rect 7630 11657 7658 11662
rect 7182 11633 7210 11639
rect 7182 11607 7183 11633
rect 7209 11607 7210 11633
rect 7182 11578 7210 11607
rect 7574 11578 7602 11583
rect 7182 11545 7210 11550
rect 7546 11577 7602 11578
rect 7546 11551 7575 11577
rect 7601 11551 7602 11577
rect 7546 11545 7602 11551
rect 7686 11577 7714 11583
rect 7686 11551 7687 11577
rect 7713 11551 7714 11577
rect 7126 11466 7154 11471
rect 7126 11419 7154 11438
rect 7294 11466 7322 11471
rect 7294 11465 7490 11466
rect 7294 11439 7295 11465
rect 7321 11439 7490 11465
rect 7294 11438 7490 11439
rect 7294 11433 7322 11438
rect 7126 11129 7154 11135
rect 7126 11103 7127 11129
rect 7153 11103 7154 11129
rect 7126 10906 7154 11103
rect 7126 10873 7154 10878
rect 7350 11130 7378 11135
rect 7070 10817 7098 10822
rect 7014 10767 7015 10793
rect 7041 10767 7042 10793
rect 7014 10761 7042 10767
rect 7238 10793 7266 10799
rect 7238 10767 7239 10793
rect 7265 10767 7266 10793
rect 7238 10570 7266 10767
rect 7350 10793 7378 11102
rect 7350 10767 7351 10793
rect 7377 10767 7378 10793
rect 7350 10761 7378 10767
rect 7462 10793 7490 11438
rect 7546 11410 7574 11545
rect 7546 11382 7602 11410
rect 7574 11186 7602 11382
rect 7686 11242 7714 11551
rect 7742 11578 7770 11583
rect 7742 11531 7770 11550
rect 7798 11577 7826 12670
rect 8190 12698 8218 13119
rect 8414 13146 8442 13151
rect 8414 12754 8442 13118
rect 8750 13090 8778 13426
rect 9254 13426 9338 13454
rect 9366 13426 9450 13454
rect 10262 13481 10290 13487
rect 10262 13455 10263 13481
rect 10289 13455 10290 13481
rect 9254 13257 9282 13426
rect 9254 13231 9255 13257
rect 9281 13231 9282 13257
rect 9254 13225 9282 13231
rect 9310 13258 9338 13263
rect 9366 13258 9394 13426
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9310 13257 9394 13258
rect 9310 13231 9311 13257
rect 9337 13231 9394 13257
rect 9310 13230 9394 13231
rect 9310 13225 9338 13230
rect 8750 13043 8778 13062
rect 9142 13145 9170 13151
rect 9142 13119 9143 13145
rect 9169 13119 9170 13145
rect 9142 12810 9170 13119
rect 9142 12777 9170 12782
rect 9198 13145 9226 13151
rect 9198 13119 9199 13145
rect 9225 13119 9226 13145
rect 8414 12721 8442 12726
rect 8190 12665 8218 12670
rect 9198 12642 9226 13119
rect 9198 12609 9226 12614
rect 9366 13146 9394 13151
rect 9310 12474 9338 12479
rect 9366 12474 9394 13118
rect 9590 13145 9618 13151
rect 9590 13119 9591 13145
rect 9617 13119 9618 13145
rect 9590 13090 9618 13119
rect 9590 13057 9618 13062
rect 9982 13090 10010 13095
rect 10262 13090 10290 13455
rect 10878 13481 10906 18999
rect 12390 19025 12418 19031
rect 12390 18999 12391 19025
rect 12417 18999 12418 19025
rect 11382 18746 11410 18751
rect 11382 18699 11410 18718
rect 10990 18633 11018 18639
rect 10990 18607 10991 18633
rect 11017 18607 11018 18633
rect 10990 13538 11018 18607
rect 10990 13537 11074 13538
rect 10990 13511 10991 13537
rect 11017 13511 11074 13537
rect 10990 13510 11074 13511
rect 10990 13505 11018 13510
rect 10878 13455 10879 13481
rect 10905 13455 10906 13481
rect 10878 13449 10906 13455
rect 9982 13089 10066 13090
rect 9982 13063 9983 13089
rect 10009 13063 10066 13089
rect 9982 13062 10066 13063
rect 9982 13057 10010 13062
rect 9814 12810 9842 12815
rect 9814 12809 10010 12810
rect 9814 12783 9815 12809
rect 9841 12783 10010 12809
rect 9814 12782 10010 12783
rect 9814 12777 9842 12782
rect 9982 12753 10010 12782
rect 10038 12809 10066 13062
rect 10262 13057 10290 13062
rect 10934 13090 10962 13095
rect 10038 12783 10039 12809
rect 10065 12783 10066 12809
rect 10038 12777 10066 12783
rect 10654 12810 10682 12815
rect 9982 12727 9983 12753
rect 10009 12727 10010 12753
rect 9982 12721 10010 12727
rect 10318 12754 10346 12759
rect 10598 12754 10626 12759
rect 10318 12753 10626 12754
rect 10318 12727 10319 12753
rect 10345 12727 10599 12753
rect 10625 12727 10626 12753
rect 10318 12726 10626 12727
rect 10318 12721 10346 12726
rect 10598 12721 10626 12726
rect 9646 12698 9674 12703
rect 9646 12651 9674 12670
rect 9310 12473 9394 12474
rect 9310 12447 9311 12473
rect 9337 12447 9394 12473
rect 9310 12446 9394 12447
rect 9758 12642 9786 12647
rect 9310 12441 9338 12446
rect 7798 11551 7799 11577
rect 7825 11551 7826 11577
rect 7686 11209 7714 11214
rect 7574 11153 7602 11158
rect 7742 11074 7770 11079
rect 7686 11046 7742 11074
rect 7462 10767 7463 10793
rect 7489 10767 7490 10793
rect 7294 10738 7322 10743
rect 7294 10691 7322 10710
rect 7406 10738 7434 10743
rect 7014 10542 7266 10570
rect 7014 10513 7042 10542
rect 7014 10487 7015 10513
rect 7041 10487 7042 10513
rect 7014 10481 7042 10487
rect 6790 10431 6791 10457
rect 6817 10431 6818 10457
rect 6454 10402 6482 10407
rect 6454 10355 6482 10374
rect 6790 10402 6818 10431
rect 6958 10458 6986 10463
rect 6958 10411 6986 10430
rect 6790 10369 6818 10374
rect 7238 10402 7266 10407
rect 7238 10355 7266 10374
rect 7406 10346 7434 10710
rect 7462 10513 7490 10767
rect 7462 10487 7463 10513
rect 7489 10487 7490 10513
rect 7462 10481 7490 10487
rect 7518 10850 7546 10855
rect 7518 10401 7546 10822
rect 7518 10375 7519 10401
rect 7545 10375 7546 10401
rect 7518 10369 7546 10375
rect 7574 10793 7602 10799
rect 7574 10767 7575 10793
rect 7601 10767 7602 10793
rect 7462 10346 7490 10351
rect 7406 10345 7490 10346
rect 7406 10319 7463 10345
rect 7489 10319 7490 10345
rect 7406 10318 7490 10319
rect 7462 10313 7490 10318
rect 7574 10094 7602 10767
rect 7462 10066 7602 10094
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 966 9673 994 9679
rect 966 9647 967 9673
rect 993 9647 994 9673
rect 966 9450 994 9647
rect 7238 9674 7266 9679
rect 966 9417 994 9422
rect 2142 9617 2170 9623
rect 2142 9591 2143 9617
rect 2169 9591 2170 9617
rect 2142 9170 2170 9591
rect 7182 9617 7210 9623
rect 7182 9591 7183 9617
rect 7209 9591 7210 9617
rect 6678 9506 6706 9511
rect 6678 9225 6706 9478
rect 6678 9199 6679 9225
rect 6705 9199 6706 9225
rect 6678 9193 6706 9199
rect 7070 9225 7098 9231
rect 7070 9199 7071 9225
rect 7097 9199 7098 9225
rect 2142 9137 2170 9142
rect 5614 9170 5642 9175
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 5614 8778 5642 9142
rect 7070 8890 7098 9199
rect 7182 8945 7210 9591
rect 7238 9617 7266 9646
rect 7238 9591 7239 9617
rect 7265 9591 7266 9617
rect 7238 9585 7266 9591
rect 7462 9617 7490 10066
rect 7574 10028 7602 10038
rect 7462 9591 7463 9617
rect 7489 9591 7490 9617
rect 7462 9585 7490 9591
rect 7574 9954 7602 9959
rect 7294 9506 7322 9511
rect 7294 9459 7322 9478
rect 7350 9505 7378 9511
rect 7350 9479 7351 9505
rect 7377 9479 7378 9505
rect 7350 9282 7378 9479
rect 7294 9254 7378 9282
rect 7574 9338 7602 9926
rect 7686 9786 7714 11046
rect 7742 11041 7770 11046
rect 7742 10962 7770 10967
rect 7742 10793 7770 10934
rect 7742 10767 7743 10793
rect 7769 10767 7770 10793
rect 7742 9954 7770 10767
rect 7742 9921 7770 9926
rect 7798 9842 7826 11551
rect 7854 12362 7882 12367
rect 7854 10738 7882 12334
rect 7966 12361 7994 12367
rect 7966 12335 7967 12361
rect 7993 12335 7994 12361
rect 7910 12306 7938 12311
rect 7966 12306 7994 12335
rect 9422 12361 9450 12367
rect 9422 12335 9423 12361
rect 9449 12335 9450 12361
rect 8190 12306 8218 12311
rect 7966 12305 8218 12306
rect 7966 12279 8191 12305
rect 8217 12279 8218 12305
rect 7966 12278 8218 12279
rect 7910 12259 7938 12278
rect 7910 11578 7938 11583
rect 7910 11577 7994 11578
rect 7910 11551 7911 11577
rect 7937 11551 7994 11577
rect 7910 11550 7994 11551
rect 7910 11545 7938 11550
rect 7910 10850 7938 10855
rect 7910 10803 7938 10822
rect 7854 9954 7882 10710
rect 7966 10458 7994 11550
rect 8022 11074 8050 12278
rect 8190 12082 8218 12278
rect 8190 12049 8218 12054
rect 9422 12026 9450 12335
rect 9254 11998 9450 12026
rect 8806 11969 8834 11975
rect 8806 11943 8807 11969
rect 8833 11943 8834 11969
rect 8358 11914 8386 11919
rect 8302 11522 8330 11527
rect 8302 11475 8330 11494
rect 8022 11041 8050 11046
rect 8190 11241 8218 11247
rect 8190 11215 8191 11241
rect 8217 11215 8218 11241
rect 8190 11130 8218 11215
rect 8358 11185 8386 11886
rect 8694 11857 8722 11863
rect 8694 11831 8695 11857
rect 8721 11831 8722 11857
rect 8414 11242 8442 11247
rect 8414 11195 8442 11214
rect 8358 11159 8359 11185
rect 8385 11159 8386 11185
rect 8358 11153 8386 11159
rect 8638 11186 8666 11191
rect 8638 11139 8666 11158
rect 8022 10962 8050 10967
rect 8022 10905 8050 10934
rect 8022 10879 8023 10905
rect 8049 10879 8050 10905
rect 8022 10873 8050 10879
rect 8078 10906 8106 10911
rect 8078 10859 8106 10878
rect 7966 10065 7994 10430
rect 8134 10793 8162 10799
rect 8134 10767 8135 10793
rect 8161 10767 8162 10793
rect 8134 10094 8162 10767
rect 8190 10402 8218 11102
rect 8470 11074 8498 11079
rect 8470 11027 8498 11046
rect 8694 10962 8722 11831
rect 8694 10929 8722 10934
rect 8750 11521 8778 11527
rect 8750 11495 8751 11521
rect 8777 11495 8778 11521
rect 8750 10850 8778 11495
rect 8806 11242 8834 11943
rect 9198 11802 9226 11807
rect 9142 11774 9198 11802
rect 9086 11634 9114 11639
rect 9086 11587 9114 11606
rect 8862 11298 8890 11303
rect 8862 11251 8890 11270
rect 8806 11209 8834 11214
rect 9086 11185 9114 11191
rect 9086 11159 9087 11185
rect 9113 11159 9114 11185
rect 8806 11130 8834 11135
rect 8806 11083 8834 11102
rect 9086 11130 9114 11159
rect 9086 11097 9114 11102
rect 9086 10906 9114 10911
rect 9142 10906 9170 11774
rect 9198 11769 9226 11774
rect 9086 10905 9170 10906
rect 9086 10879 9087 10905
rect 9113 10879 9170 10905
rect 9086 10878 9170 10879
rect 9086 10873 9114 10878
rect 8750 10817 8778 10822
rect 8918 10849 8946 10855
rect 8918 10823 8919 10849
rect 8945 10823 8946 10849
rect 8246 10402 8274 10407
rect 8190 10401 8274 10402
rect 8190 10375 8247 10401
rect 8273 10375 8274 10401
rect 8190 10374 8274 10375
rect 8246 10369 8274 10374
rect 8414 10290 8442 10295
rect 8414 10289 8498 10290
rect 8414 10263 8415 10289
rect 8441 10263 8498 10289
rect 8414 10262 8498 10263
rect 8414 10257 8442 10262
rect 8414 10122 8442 10127
rect 7966 10039 7967 10065
rect 7993 10039 7994 10065
rect 7966 10033 7994 10039
rect 8078 10066 8106 10071
rect 8134 10066 8218 10094
rect 8078 10019 8106 10038
rect 7854 9921 7882 9926
rect 8022 10009 8050 10015
rect 8022 9983 8023 10009
rect 8049 9983 8050 10009
rect 7798 9814 7882 9842
rect 7686 9758 7826 9786
rect 7686 9674 7714 9679
rect 7686 9627 7714 9646
rect 7574 9281 7602 9310
rect 7574 9255 7575 9281
rect 7601 9255 7602 9281
rect 7182 8919 7183 8945
rect 7209 8919 7210 8945
rect 7182 8913 7210 8919
rect 7238 9170 7266 9175
rect 7070 8857 7098 8862
rect 7238 8833 7266 9142
rect 7238 8807 7239 8833
rect 7265 8807 7266 8833
rect 7238 8801 7266 8807
rect 5614 8745 5642 8750
rect 7182 8778 7210 8783
rect 7182 8731 7210 8750
rect 7238 8554 7266 8559
rect 7294 8554 7322 9254
rect 7574 9249 7602 9255
rect 7630 9394 7658 9399
rect 7630 9281 7658 9366
rect 7798 9338 7826 9758
rect 7854 9506 7882 9814
rect 8022 9618 8050 9983
rect 8134 10010 8162 10015
rect 8190 10010 8218 10066
rect 8246 10010 8274 10015
rect 8414 10010 8442 10094
rect 8190 10009 8442 10010
rect 8190 9983 8247 10009
rect 8273 9983 8442 10009
rect 8190 9982 8442 9983
rect 8134 9963 8162 9982
rect 8246 9977 8274 9982
rect 8302 9730 8330 9735
rect 8134 9729 8330 9730
rect 8134 9703 8303 9729
rect 8329 9703 8330 9729
rect 8134 9702 8330 9703
rect 8078 9618 8106 9623
rect 8134 9618 8162 9702
rect 8302 9697 8330 9702
rect 8022 9617 8162 9618
rect 8022 9591 8079 9617
rect 8105 9591 8162 9617
rect 8022 9590 8162 9591
rect 8414 9618 8442 9982
rect 8470 9730 8498 10262
rect 8918 10122 8946 10823
rect 9254 10346 9282 11998
rect 9478 11970 9506 11975
rect 9310 11969 9506 11970
rect 9310 11943 9479 11969
rect 9505 11943 9506 11969
rect 9310 11942 9506 11943
rect 9310 11633 9338 11942
rect 9478 11937 9506 11942
rect 9590 11970 9618 11975
rect 9590 11923 9618 11942
rect 9646 11913 9674 11919
rect 9646 11887 9647 11913
rect 9673 11887 9674 11913
rect 9310 11607 9311 11633
rect 9337 11607 9338 11633
rect 9310 11298 9338 11607
rect 9366 11802 9394 11807
rect 9366 11577 9394 11774
rect 9366 11551 9367 11577
rect 9393 11551 9394 11577
rect 9366 11545 9394 11551
rect 9422 11634 9450 11639
rect 9310 11185 9338 11270
rect 9310 11159 9311 11185
rect 9337 11159 9338 11185
rect 9310 11153 9338 11159
rect 9422 11186 9450 11606
rect 9646 11186 9674 11887
rect 9254 10094 9282 10318
rect 8918 10089 8946 10094
rect 8974 10066 9282 10094
rect 8974 10065 9002 10066
rect 8974 10039 8975 10065
rect 9001 10039 9002 10065
rect 8974 10033 9002 10039
rect 8694 10010 8722 10015
rect 8918 10010 8946 10015
rect 8694 10009 8890 10010
rect 8694 9983 8695 10009
rect 8721 9983 8890 10009
rect 8694 9982 8890 9983
rect 8694 9977 8722 9982
rect 8806 9897 8834 9903
rect 8806 9871 8807 9897
rect 8833 9871 8834 9897
rect 8806 9730 8834 9871
rect 8470 9729 8834 9730
rect 8470 9703 8471 9729
rect 8497 9703 8834 9729
rect 8470 9702 8834 9703
rect 8470 9697 8498 9702
rect 8414 9590 8498 9618
rect 8078 9585 8106 9590
rect 7966 9506 7994 9511
rect 7854 9505 7994 9506
rect 7854 9479 7967 9505
rect 7993 9479 7994 9505
rect 7854 9478 7994 9479
rect 7742 9337 7826 9338
rect 7742 9311 7799 9337
rect 7825 9311 7826 9337
rect 7742 9310 7826 9311
rect 7630 9255 7631 9281
rect 7657 9255 7658 9281
rect 7630 9249 7658 9255
rect 7686 9282 7714 9287
rect 7686 9235 7714 9254
rect 7406 9170 7434 9175
rect 7406 9169 7546 9170
rect 7406 9143 7407 9169
rect 7433 9143 7546 9169
rect 7406 9142 7546 9143
rect 7406 9137 7434 9142
rect 7350 8890 7378 8895
rect 7462 8890 7490 8895
rect 7378 8889 7490 8890
rect 7378 8863 7463 8889
rect 7489 8863 7490 8889
rect 7378 8862 7490 8863
rect 7350 8857 7378 8862
rect 7266 8526 7322 8554
rect 7238 8507 7266 8526
rect 2142 8442 2170 8447
rect 2142 8395 2170 8414
rect 5950 8442 5978 8447
rect 966 8329 994 8335
rect 966 8303 967 8329
rect 993 8303 994 8329
rect 966 8106 994 8303
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 966 8073 994 8078
rect 5950 7601 5978 8414
rect 7126 8441 7154 8447
rect 7126 8415 7127 8441
rect 7153 8415 7154 8441
rect 7126 8386 7154 8415
rect 7126 8353 7154 8358
rect 7182 8385 7210 8391
rect 7182 8359 7183 8385
rect 7209 8359 7210 8385
rect 7014 7714 7042 7719
rect 7182 7714 7210 8359
rect 7014 7713 7210 7714
rect 7014 7687 7015 7713
rect 7041 7687 7210 7713
rect 7014 7686 7210 7687
rect 7406 7714 7434 8862
rect 7462 8857 7490 8862
rect 7462 8442 7490 8447
rect 7518 8442 7546 9142
rect 7742 9058 7770 9310
rect 7798 9305 7826 9310
rect 7910 9394 7938 9399
rect 7910 9337 7938 9366
rect 7910 9311 7911 9337
rect 7937 9311 7938 9337
rect 7910 9305 7938 9311
rect 7742 9030 7938 9058
rect 7798 8890 7826 8895
rect 7910 8890 7938 9030
rect 7966 9002 7994 9478
rect 8358 9506 8386 9511
rect 8414 9506 8442 9511
rect 8358 9505 8414 9506
rect 8358 9479 8359 9505
rect 8385 9479 8414 9505
rect 8358 9478 8414 9479
rect 8078 9450 8106 9455
rect 8022 9281 8050 9287
rect 8022 9255 8023 9281
rect 8049 9255 8050 9281
rect 8022 9114 8050 9255
rect 8078 9281 8106 9422
rect 8078 9255 8079 9281
rect 8105 9255 8106 9281
rect 8078 9249 8106 9255
rect 8022 9081 8050 9086
rect 8246 9225 8274 9231
rect 8246 9199 8247 9225
rect 8273 9199 8274 9225
rect 8246 9170 8274 9199
rect 7966 8969 7994 8974
rect 7966 8890 7994 8895
rect 7910 8889 7994 8890
rect 7910 8863 7967 8889
rect 7993 8863 7994 8889
rect 7910 8862 7994 8863
rect 7742 8778 7770 8783
rect 7630 8498 7658 8503
rect 7742 8498 7770 8750
rect 7630 8451 7658 8470
rect 7686 8497 7770 8498
rect 7686 8471 7743 8497
rect 7769 8471 7770 8497
rect 7686 8470 7770 8471
rect 7462 8441 7546 8442
rect 7462 8415 7463 8441
rect 7489 8415 7546 8441
rect 7462 8414 7546 8415
rect 7462 8409 7490 8414
rect 7574 8386 7602 8391
rect 7574 8339 7602 8358
rect 7630 7714 7658 7719
rect 7406 7686 7630 7714
rect 7014 7681 7042 7686
rect 7406 7657 7434 7686
rect 7630 7667 7658 7686
rect 7406 7631 7407 7657
rect 7433 7631 7434 7657
rect 7406 7625 7434 7631
rect 5950 7575 5951 7601
rect 5977 7575 5978 7601
rect 5950 7569 5978 7575
rect 7462 7602 7490 7607
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 7462 7377 7490 7574
rect 7462 7351 7463 7377
rect 7489 7351 7490 7377
rect 7462 7345 7490 7351
rect 7630 7378 7658 7383
rect 7686 7378 7714 8470
rect 7742 8465 7770 8470
rect 7630 7377 7714 7378
rect 7630 7351 7631 7377
rect 7657 7351 7714 7377
rect 7630 7350 7714 7351
rect 7630 7345 7658 7350
rect 7798 7321 7826 8862
rect 7966 8857 7994 8862
rect 8246 8890 8274 9142
rect 8246 8857 8274 8862
rect 8358 8833 8386 9478
rect 8414 9473 8442 9478
rect 8414 9281 8442 9287
rect 8414 9255 8415 9281
rect 8441 9255 8442 9281
rect 8414 9226 8442 9255
rect 8414 9193 8442 9198
rect 8358 8807 8359 8833
rect 8385 8807 8386 8833
rect 8358 8801 8386 8807
rect 8246 8778 8274 8783
rect 8246 8731 8274 8750
rect 8022 8106 8050 8111
rect 8022 7657 8050 8078
rect 8470 8050 8498 9590
rect 8638 9617 8666 9702
rect 8638 9591 8639 9617
rect 8665 9591 8666 9617
rect 8638 9585 8666 9591
rect 8806 9225 8834 9702
rect 8806 9199 8807 9225
rect 8833 9199 8834 9225
rect 8806 9193 8834 9199
rect 8862 9618 8890 9982
rect 8918 9730 8946 9982
rect 9142 10009 9170 10015
rect 9142 9983 9143 10009
rect 9169 9983 9170 10009
rect 8974 9730 9002 9735
rect 8918 9702 8974 9730
rect 8974 9683 9002 9702
rect 9142 9618 9170 9983
rect 9254 9954 9282 9959
rect 9254 9729 9282 9926
rect 9422 9954 9450 11158
rect 9590 11158 9674 11186
rect 9702 11186 9730 11191
rect 9758 11186 9786 12614
rect 10094 12641 10122 12647
rect 10094 12615 10095 12641
rect 10121 12615 10122 12641
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 10094 12082 10122 12615
rect 10318 12417 10346 12423
rect 10318 12391 10319 12417
rect 10345 12391 10346 12417
rect 10150 12362 10178 12367
rect 10178 12334 10234 12362
rect 10150 12329 10178 12334
rect 10206 12305 10234 12334
rect 10206 12279 10207 12305
rect 10233 12279 10234 12305
rect 10206 12273 10234 12279
rect 10038 12054 10122 12082
rect 9982 11969 10010 11975
rect 9982 11943 9983 11969
rect 10009 11943 10010 11969
rect 9982 11914 10010 11943
rect 9982 11881 10010 11886
rect 9814 11857 9842 11863
rect 9814 11831 9815 11857
rect 9841 11831 9842 11857
rect 9814 11802 9842 11831
rect 10038 11858 10066 12054
rect 10318 12026 10346 12391
rect 10374 12306 10402 12311
rect 10374 12259 10402 12278
rect 10374 12026 10402 12031
rect 10318 11998 10374 12026
rect 10374 11993 10402 11998
rect 10094 11970 10122 11975
rect 10094 11969 10290 11970
rect 10094 11943 10095 11969
rect 10121 11943 10290 11969
rect 10094 11942 10290 11943
rect 10094 11937 10122 11942
rect 10206 11858 10234 11863
rect 10038 11830 10206 11858
rect 10262 11858 10290 11942
rect 10374 11914 10402 11919
rect 10318 11858 10346 11863
rect 10262 11857 10346 11858
rect 10262 11831 10319 11857
rect 10345 11831 10346 11857
rect 10262 11830 10346 11831
rect 10206 11811 10234 11830
rect 9814 11769 9842 11774
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 10094 11522 10122 11527
rect 9814 11186 9842 11191
rect 9758 11158 9814 11186
rect 9590 10850 9618 11158
rect 9702 11139 9730 11158
rect 9814 11153 9842 11158
rect 9926 11185 9954 11191
rect 9926 11159 9927 11185
rect 9953 11159 9954 11185
rect 9926 11130 9954 11159
rect 9982 11186 10010 11191
rect 9982 11139 10010 11158
rect 9926 11097 9954 11102
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 9926 10906 9954 10911
rect 9590 10822 9674 10850
rect 9590 10738 9618 10743
rect 9590 10691 9618 10710
rect 9422 9907 9450 9926
rect 9254 9703 9255 9729
rect 9281 9703 9282 9729
rect 9254 9697 9282 9703
rect 8862 9617 9170 9618
rect 8862 9591 8863 9617
rect 8889 9591 9170 9617
rect 8862 9590 9170 9591
rect 9310 9674 9338 9679
rect 9310 9617 9338 9646
rect 9310 9591 9311 9617
rect 9337 9591 9338 9617
rect 8862 9226 8890 9590
rect 8862 8834 8890 9198
rect 8918 9338 8946 9343
rect 9142 9338 9170 9343
rect 8918 8889 8946 9310
rect 9086 9310 9142 9338
rect 9030 9226 9058 9231
rect 9030 9179 9058 9198
rect 9030 8946 9058 8951
rect 9086 8946 9114 9310
rect 9142 9305 9170 9310
rect 9310 9282 9338 9591
rect 9646 9618 9674 10822
rect 9870 10794 9898 10799
rect 9870 10747 9898 10766
rect 9702 10514 9730 10519
rect 9730 10486 9786 10514
rect 9702 10481 9730 10486
rect 9758 10066 9786 10486
rect 9926 10513 9954 10878
rect 9926 10487 9927 10513
rect 9953 10487 9954 10513
rect 9926 10481 9954 10487
rect 9870 10458 9898 10463
rect 9870 10411 9898 10430
rect 9814 10402 9842 10407
rect 9814 10345 9842 10374
rect 9814 10319 9815 10345
rect 9841 10319 9842 10345
rect 9814 10313 9842 10319
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9870 10066 9898 10071
rect 9758 10065 9898 10066
rect 9758 10039 9871 10065
rect 9897 10039 9898 10065
rect 9758 10038 9898 10039
rect 9870 10033 9898 10038
rect 10038 10010 10066 10015
rect 10094 10010 10122 11494
rect 10318 11242 10346 11830
rect 10150 11214 10346 11242
rect 10150 10962 10178 11214
rect 10374 11186 10402 11886
rect 10150 10929 10178 10934
rect 10206 11158 10402 11186
rect 10206 11129 10234 11158
rect 10206 11103 10207 11129
rect 10233 11103 10234 11129
rect 10066 9982 10122 10010
rect 10150 10850 10178 10855
rect 10150 10457 10178 10822
rect 10206 10794 10234 11103
rect 10430 11130 10458 11135
rect 10262 11074 10290 11079
rect 10262 11073 10402 11074
rect 10262 11047 10263 11073
rect 10289 11047 10402 11073
rect 10262 11046 10402 11047
rect 10262 11041 10290 11046
rect 10206 10761 10234 10766
rect 10262 10962 10290 10967
rect 10150 10431 10151 10457
rect 10177 10431 10178 10457
rect 10150 10402 10178 10431
rect 10038 9963 10066 9982
rect 9366 9562 9394 9567
rect 9366 9515 9394 9534
rect 9310 9249 9338 9254
rect 9646 9338 9674 9590
rect 9814 9730 9842 9735
rect 10150 9730 10178 10374
rect 10206 10122 10234 10127
rect 10262 10122 10290 10934
rect 10374 10906 10402 11046
rect 10374 10873 10402 10878
rect 10430 10849 10458 11102
rect 10654 11129 10682 12782
rect 10934 12753 10962 13062
rect 10934 12727 10935 12753
rect 10961 12727 10962 12753
rect 10934 12721 10962 12727
rect 11046 13089 11074 13510
rect 11046 13063 11047 13089
rect 11073 13063 11074 13089
rect 10710 12698 10738 12703
rect 10710 12651 10738 12670
rect 10766 12697 10794 12703
rect 10766 12671 10767 12697
rect 10793 12671 10794 12697
rect 10654 11103 10655 11129
rect 10681 11103 10682 11129
rect 10430 10823 10431 10849
rect 10457 10823 10458 10849
rect 10430 10817 10458 10823
rect 10598 11074 10626 11079
rect 10542 10794 10570 10799
rect 10206 10121 10290 10122
rect 10206 10095 10207 10121
rect 10233 10095 10290 10121
rect 10206 10094 10290 10095
rect 10318 10401 10346 10407
rect 10318 10375 10319 10401
rect 10345 10375 10346 10401
rect 10206 10089 10234 10094
rect 10318 10009 10346 10375
rect 10542 10121 10570 10766
rect 10598 10738 10626 11046
rect 10654 11018 10682 11103
rect 10654 10985 10682 10990
rect 10766 12306 10794 12671
rect 11046 12698 11074 13063
rect 11270 13090 11298 13095
rect 11270 13043 11298 13062
rect 11494 13090 11522 13095
rect 11494 13043 11522 13062
rect 12390 12809 12418 18999
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 13062 13202 13090 13207
rect 13062 13155 13090 13174
rect 13118 13146 13146 13151
rect 14014 13146 14042 13151
rect 13118 13145 13202 13146
rect 13118 13119 13119 13145
rect 13145 13119 13202 13145
rect 13118 13118 13202 13119
rect 13118 13113 13146 13118
rect 12390 12783 12391 12809
rect 12417 12783 12418 12809
rect 11326 12698 11354 12703
rect 11046 12665 11074 12670
rect 11270 12697 11354 12698
rect 11270 12671 11327 12697
rect 11353 12671 11354 12697
rect 11270 12670 11354 12671
rect 11270 12473 11298 12670
rect 11326 12665 11354 12670
rect 11774 12474 11802 12479
rect 11270 12447 11271 12473
rect 11297 12447 11298 12473
rect 11270 12441 11298 12447
rect 11438 12473 11802 12474
rect 11438 12447 11775 12473
rect 11801 12447 11802 12473
rect 11438 12446 11802 12447
rect 11438 12417 11466 12446
rect 11774 12441 11802 12446
rect 11438 12391 11439 12417
rect 11465 12391 11466 12417
rect 11438 12385 11466 12391
rect 11942 12418 11970 12423
rect 12390 12418 12418 12783
rect 12614 13090 12642 13095
rect 12670 13090 12698 13095
rect 12642 13089 12698 13090
rect 12642 13063 12671 13089
rect 12697 13063 12698 13089
rect 12642 13062 12698 13063
rect 12614 12754 12642 13062
rect 12670 13057 12698 13062
rect 13174 13090 13202 13118
rect 13342 13090 13370 13095
rect 13174 13089 13370 13090
rect 13174 13063 13343 13089
rect 13369 13063 13370 13089
rect 13174 13062 13370 13063
rect 13062 13033 13090 13039
rect 13062 13007 13063 13033
rect 13089 13007 13090 13033
rect 12614 12753 12698 12754
rect 12614 12727 12615 12753
rect 12641 12727 12698 12753
rect 12614 12726 12698 12727
rect 12614 12721 12642 12726
rect 11942 12417 12418 12418
rect 11942 12391 11943 12417
rect 11969 12391 12418 12417
rect 11942 12390 12418 12391
rect 12670 12642 12698 12726
rect 12950 12698 12978 12703
rect 12670 12473 12698 12614
rect 12670 12447 12671 12473
rect 12697 12447 12698 12473
rect 11942 12385 11970 12390
rect 11102 12361 11130 12367
rect 11102 12335 11103 12361
rect 11129 12335 11130 12361
rect 10878 12306 10906 12311
rect 10766 12305 10906 12306
rect 10766 12279 10879 12305
rect 10905 12279 10906 12305
rect 10766 12278 10906 12279
rect 10766 11858 10794 12278
rect 10878 12273 10906 12278
rect 11102 12306 11130 12335
rect 11102 12273 11130 12278
rect 11270 12361 11298 12367
rect 11270 12335 11271 12361
rect 11297 12335 11298 12361
rect 11214 12082 11242 12087
rect 11214 12035 11242 12054
rect 10598 10705 10626 10710
rect 10654 10793 10682 10799
rect 10654 10767 10655 10793
rect 10681 10767 10682 10793
rect 10542 10095 10543 10121
rect 10569 10095 10570 10121
rect 10542 10089 10570 10095
rect 10318 9983 10319 10009
rect 10345 9983 10346 10009
rect 10206 9898 10234 9903
rect 10234 9870 10290 9898
rect 10206 9865 10234 9870
rect 10150 9702 10234 9730
rect 9702 9562 9730 9567
rect 9702 9515 9730 9534
rect 9758 9561 9786 9567
rect 9758 9535 9759 9561
rect 9785 9535 9786 9561
rect 9758 9394 9786 9535
rect 9254 9225 9282 9231
rect 9254 9199 9255 9225
rect 9281 9199 9282 9225
rect 9254 9170 9282 9199
rect 9254 9137 9282 9142
rect 9590 9225 9618 9231
rect 9590 9199 9591 9225
rect 9617 9199 9618 9225
rect 9590 9170 9618 9199
rect 9590 9137 9618 9142
rect 9646 9169 9674 9310
rect 9702 9366 9786 9394
rect 9702 9226 9730 9366
rect 9758 9282 9786 9287
rect 9758 9235 9786 9254
rect 9702 9193 9730 9198
rect 9646 9143 9647 9169
rect 9673 9143 9674 9169
rect 9646 9137 9674 9143
rect 9030 8945 9114 8946
rect 9030 8919 9031 8945
rect 9057 8919 9114 8945
rect 9030 8918 9114 8919
rect 9534 9114 9562 9119
rect 9030 8913 9058 8918
rect 8918 8863 8919 8889
rect 8945 8863 8946 8889
rect 8918 8857 8946 8863
rect 8862 8801 8890 8806
rect 9366 8834 9394 8839
rect 9366 8787 9394 8806
rect 9534 8777 9562 9086
rect 9814 8833 9842 9702
rect 9926 9674 9954 9679
rect 10094 9674 10122 9679
rect 9926 9506 9954 9646
rect 10038 9646 10094 9674
rect 9982 9618 10010 9623
rect 9982 9571 10010 9590
rect 10038 9617 10066 9646
rect 10094 9641 10122 9646
rect 10038 9591 10039 9617
rect 10065 9591 10066 9617
rect 10038 9585 10066 9591
rect 10206 9562 10234 9702
rect 10262 9617 10290 9870
rect 10262 9591 10263 9617
rect 10289 9591 10290 9617
rect 10262 9585 10290 9591
rect 10318 9618 10346 9983
rect 10654 9954 10682 10767
rect 10150 9534 10234 9562
rect 10094 9506 10122 9511
rect 9926 9478 10094 9506
rect 10094 9459 10122 9478
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 10150 9338 10178 9534
rect 10094 9310 10178 9338
rect 9982 9282 10010 9287
rect 10094 9282 10122 9310
rect 9982 9281 10122 9282
rect 9982 9255 9983 9281
rect 10009 9255 10122 9281
rect 9982 9254 10122 9255
rect 10318 9282 10346 9590
rect 9982 9249 10010 9254
rect 10318 9249 10346 9254
rect 10430 9674 10458 9679
rect 10430 9226 10458 9646
rect 10654 9673 10682 9926
rect 10654 9647 10655 9673
rect 10681 9647 10682 9673
rect 10654 9641 10682 9647
rect 10710 10009 10738 10015
rect 10710 9983 10711 10009
rect 10737 9983 10738 10009
rect 10710 9674 10738 9983
rect 10766 9786 10794 11830
rect 10878 12026 10906 12031
rect 10878 11914 10906 11998
rect 10990 11970 11018 11975
rect 10934 11969 11018 11970
rect 10934 11943 10991 11969
rect 11017 11943 11018 11969
rect 10934 11942 11018 11943
rect 10934 11914 10962 11942
rect 10990 11937 11018 11942
rect 10878 11886 10962 11914
rect 11270 11914 11298 12335
rect 11662 12361 11690 12367
rect 11662 12335 11663 12361
rect 11689 12335 11690 12361
rect 11550 11970 11578 11975
rect 11550 11923 11578 11942
rect 11298 11886 11410 11914
rect 10822 11185 10850 11191
rect 10822 11159 10823 11185
rect 10849 11159 10850 11185
rect 10822 10962 10850 11159
rect 10822 10929 10850 10934
rect 10878 10906 10906 11886
rect 11270 11867 11298 11886
rect 11046 11185 11074 11191
rect 11046 11159 11047 11185
rect 11073 11159 11074 11185
rect 11046 11074 11074 11159
rect 11382 11129 11410 11886
rect 11438 11858 11466 11863
rect 11438 11811 11466 11830
rect 11662 11186 11690 12335
rect 11662 11153 11690 11158
rect 11718 12361 11746 12367
rect 11718 12335 11719 12361
rect 11745 12335 11746 12361
rect 11382 11103 11383 11129
rect 11409 11103 11410 11129
rect 11382 11097 11410 11103
rect 11046 11041 11074 11046
rect 11214 11073 11242 11079
rect 11214 11047 11215 11073
rect 11241 11047 11242 11073
rect 11214 10962 11242 11047
rect 11214 10929 11242 10934
rect 11550 11074 11578 11079
rect 11718 11074 11746 12335
rect 11830 12361 11858 12367
rect 11830 12335 11831 12361
rect 11857 12335 11858 12361
rect 11830 11970 11858 12335
rect 12670 12362 12698 12447
rect 12894 12697 12978 12698
rect 12894 12671 12951 12697
rect 12977 12671 12978 12697
rect 12894 12670 12978 12671
rect 12838 12362 12866 12367
rect 12670 12361 12866 12362
rect 12670 12335 12839 12361
rect 12865 12335 12866 12361
rect 12670 12334 12866 12335
rect 12838 12329 12866 12334
rect 11830 11937 11858 11942
rect 12726 12194 12754 12199
rect 12726 11969 12754 12166
rect 12894 12025 12922 12670
rect 12950 12665 12978 12670
rect 12894 11999 12895 12025
rect 12921 11999 12922 12025
rect 12894 11993 12922 11999
rect 12950 12250 12978 12255
rect 12726 11943 12727 11969
rect 12753 11943 12754 11969
rect 12726 11937 12754 11943
rect 12950 11970 12978 12222
rect 13062 12194 13090 13007
rect 13062 12161 13090 12166
rect 13062 11970 13090 11975
rect 12950 11969 13090 11970
rect 12950 11943 12951 11969
rect 12977 11943 13063 11969
rect 13089 11943 13090 11969
rect 12950 11942 13090 11943
rect 12950 11937 12978 11942
rect 13062 11937 13090 11942
rect 12614 11913 12642 11919
rect 12614 11887 12615 11913
rect 12641 11887 12642 11913
rect 10822 10850 10850 10855
rect 10822 10803 10850 10822
rect 10878 10793 10906 10878
rect 10878 10767 10879 10793
rect 10905 10767 10906 10793
rect 10878 10761 10906 10767
rect 11158 10850 11186 10855
rect 10934 10514 10962 10519
rect 10934 10401 10962 10486
rect 10934 10375 10935 10401
rect 10961 10375 10962 10401
rect 10934 10369 10962 10375
rect 10878 10010 10906 10015
rect 10878 9963 10906 9982
rect 10766 9753 10794 9758
rect 10934 9898 10962 9903
rect 10934 9729 10962 9870
rect 10934 9703 10935 9729
rect 10961 9703 10962 9729
rect 10934 9697 10962 9703
rect 10710 9641 10738 9646
rect 11102 9674 11130 9679
rect 10766 9617 10794 9623
rect 10766 9591 10767 9617
rect 10793 9591 10794 9617
rect 10710 9506 10738 9511
rect 10766 9506 10794 9591
rect 10738 9478 10794 9506
rect 10430 9193 10458 9198
rect 10486 9282 10514 9287
rect 10486 9225 10514 9254
rect 10486 9199 10487 9225
rect 10513 9199 10514 9225
rect 10486 9193 10514 9199
rect 10710 9225 10738 9478
rect 11046 9226 11074 9231
rect 10710 9199 10711 9225
rect 10737 9199 10738 9225
rect 10710 9193 10738 9199
rect 10990 9198 11046 9226
rect 10038 9114 10066 9119
rect 10038 9067 10066 9086
rect 10766 9113 10794 9119
rect 10766 9087 10767 9113
rect 10793 9087 10794 9113
rect 9814 8807 9815 8833
rect 9841 8807 9842 8833
rect 9814 8801 9842 8807
rect 10038 9002 10066 9007
rect 10038 8833 10066 8974
rect 10318 8890 10346 8895
rect 10318 8889 10626 8890
rect 10318 8863 10319 8889
rect 10345 8863 10626 8889
rect 10318 8862 10626 8863
rect 10318 8857 10346 8862
rect 10038 8807 10039 8833
rect 10065 8807 10066 8833
rect 10038 8801 10066 8807
rect 10262 8834 10290 8839
rect 10262 8787 10290 8806
rect 9534 8751 9535 8777
rect 9561 8751 9562 8777
rect 9534 8745 9562 8751
rect 9198 8722 9226 8727
rect 9310 8722 9338 8727
rect 9142 8721 9226 8722
rect 9142 8695 9199 8721
rect 9225 8695 9226 8721
rect 9142 8694 9226 8695
rect 9142 8106 9170 8694
rect 9198 8689 9226 8694
rect 9254 8694 9310 8722
rect 9254 8442 9282 8694
rect 9310 8689 9338 8694
rect 9702 8722 9730 8727
rect 9702 8675 9730 8694
rect 10150 8721 10178 8727
rect 10150 8695 10151 8721
rect 10177 8695 10178 8721
rect 10150 8666 10178 8695
rect 10318 8722 10346 8727
rect 10346 8694 10402 8722
rect 10318 8675 10346 8694
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10150 8633 10178 8638
rect 9918 8605 10050 8610
rect 9142 8073 9170 8078
rect 9198 8414 9282 8442
rect 8470 8022 9114 8050
rect 8694 7769 8722 8022
rect 9086 7994 9114 8022
rect 9198 8049 9226 8414
rect 9198 8023 9199 8049
rect 9225 8023 9226 8049
rect 9198 8017 9226 8023
rect 10374 8050 10402 8694
rect 10374 8017 10402 8022
rect 9142 7994 9170 7999
rect 9086 7993 9170 7994
rect 9086 7967 9143 7993
rect 9169 7967 9170 7993
rect 9086 7966 9170 7967
rect 9142 7961 9170 7966
rect 9030 7937 9058 7943
rect 9030 7911 9031 7937
rect 9057 7911 9058 7937
rect 8694 7743 8695 7769
rect 8721 7743 8722 7769
rect 8694 7737 8722 7743
rect 8806 7770 8834 7775
rect 8806 7723 8834 7742
rect 8022 7631 8023 7657
rect 8049 7631 8050 7657
rect 8022 7625 8050 7631
rect 8078 7714 8106 7719
rect 7854 7602 7882 7621
rect 7854 7569 7882 7574
rect 7910 7601 7938 7607
rect 7910 7575 7911 7601
rect 7937 7575 7938 7601
rect 7798 7295 7799 7321
rect 7825 7295 7826 7321
rect 7798 7289 7826 7295
rect 6678 7154 6706 7159
rect 6678 6817 6706 7126
rect 7518 7154 7546 7159
rect 7910 7154 7938 7575
rect 7518 7107 7546 7126
rect 7742 7126 7938 7154
rect 7742 6929 7770 7126
rect 7742 6903 7743 6929
rect 7769 6903 7770 6929
rect 7742 6897 7770 6903
rect 8078 6986 8106 7686
rect 9030 7657 9058 7911
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 10150 7714 10178 7719
rect 10262 7714 10290 7719
rect 10150 7713 10262 7714
rect 10150 7687 10151 7713
rect 10177 7687 10262 7713
rect 10150 7686 10262 7687
rect 10150 7681 10178 7686
rect 10262 7681 10290 7686
rect 9030 7631 9031 7657
rect 9057 7631 9058 7657
rect 8750 7601 8778 7607
rect 8750 7575 8751 7601
rect 8777 7575 8778 7601
rect 8750 7378 8778 7575
rect 8750 7350 8890 7378
rect 8862 7321 8890 7350
rect 8862 7295 8863 7321
rect 8889 7295 8890 7321
rect 8862 7289 8890 7295
rect 8470 7154 8498 7159
rect 8358 6986 8386 6991
rect 8414 6986 8442 6991
rect 8078 6985 8414 6986
rect 8078 6959 8359 6985
rect 8385 6959 8414 6985
rect 8078 6958 8414 6959
rect 8078 6873 8106 6958
rect 8358 6953 8386 6958
rect 8414 6953 8442 6958
rect 8078 6847 8079 6873
rect 8105 6847 8106 6873
rect 8078 6841 8106 6847
rect 6678 6791 6679 6817
rect 6705 6791 6706 6817
rect 6678 6785 6706 6791
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8470 1777 8498 7126
rect 9030 7098 9058 7631
rect 9478 7658 9506 7663
rect 9254 7266 9282 7271
rect 9478 7266 9506 7630
rect 9758 7658 9786 7663
rect 9758 7611 9786 7630
rect 10094 7658 10122 7663
rect 10094 7490 10122 7630
rect 10094 7462 10178 7490
rect 9030 7065 9058 7070
rect 9198 7265 9506 7266
rect 9198 7239 9255 7265
rect 9281 7239 9479 7265
rect 9505 7239 9506 7265
rect 9198 7238 9506 7239
rect 8862 6986 8890 6991
rect 8862 6481 8890 6958
rect 9198 6986 9226 7238
rect 9254 7233 9282 7238
rect 9478 7233 9506 7238
rect 9422 7154 9450 7159
rect 9198 6953 9226 6958
rect 9366 7098 9394 7103
rect 9366 6985 9394 7070
rect 9366 6959 9367 6985
rect 9393 6959 9394 6985
rect 9366 6953 9394 6959
rect 9422 6929 9450 7126
rect 10094 7154 10122 7159
rect 10094 7107 10122 7126
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 10150 6986 10178 7462
rect 10262 7266 10290 7271
rect 10598 7266 10626 8862
rect 10654 8666 10682 8671
rect 10654 8049 10682 8638
rect 10710 8554 10738 8559
rect 10766 8554 10794 9087
rect 10738 8526 10794 8554
rect 10710 8521 10738 8526
rect 10654 8023 10655 8049
rect 10681 8023 10682 8049
rect 10654 8017 10682 8023
rect 10710 7937 10738 7943
rect 10710 7911 10711 7937
rect 10737 7911 10738 7937
rect 10710 7714 10738 7911
rect 10710 7681 10738 7686
rect 10766 7574 10794 8526
rect 10934 8721 10962 8727
rect 10934 8695 10935 8721
rect 10961 8695 10962 8721
rect 10934 8498 10962 8695
rect 10934 8451 10962 8470
rect 10934 8162 10962 8167
rect 10990 8162 11018 9198
rect 11046 9193 11074 9198
rect 11102 9170 11130 9646
rect 11158 9673 11186 10822
rect 11270 9953 11298 9959
rect 11270 9927 11271 9953
rect 11297 9927 11298 9953
rect 11214 9730 11242 9735
rect 11270 9730 11298 9927
rect 11214 9729 11466 9730
rect 11214 9703 11215 9729
rect 11241 9703 11466 9729
rect 11214 9702 11466 9703
rect 11214 9697 11242 9702
rect 11158 9647 11159 9673
rect 11185 9647 11186 9673
rect 11158 9641 11186 9647
rect 11102 8889 11130 9142
rect 11102 8863 11103 8889
rect 11129 8863 11130 8889
rect 11102 8857 11130 8863
rect 11214 9562 11242 9567
rect 10934 8161 11018 8162
rect 10934 8135 10935 8161
rect 10961 8135 11018 8161
rect 10934 8134 11018 8135
rect 10934 8129 10962 8134
rect 10822 8050 10850 8055
rect 10822 8003 10850 8022
rect 11046 8049 11074 8055
rect 11046 8023 11047 8049
rect 11073 8023 11074 8049
rect 11046 7882 11074 8023
rect 11214 7993 11242 9534
rect 11438 9561 11466 9702
rect 11438 9535 11439 9561
rect 11465 9535 11466 9561
rect 11438 9529 11466 9535
rect 11550 9505 11578 11046
rect 11662 11046 11718 11074
rect 11662 10682 11690 11046
rect 11718 11027 11746 11046
rect 11886 11577 11914 11583
rect 11886 11551 11887 11577
rect 11913 11551 11914 11577
rect 11718 10794 11746 10799
rect 11718 10747 11746 10766
rect 11662 10654 11746 10682
rect 11662 9730 11690 9735
rect 11550 9479 11551 9505
rect 11577 9479 11578 9505
rect 11382 9282 11410 9287
rect 11550 9282 11578 9479
rect 11606 9673 11634 9679
rect 11606 9647 11607 9673
rect 11633 9647 11634 9673
rect 11606 9450 11634 9647
rect 11662 9617 11690 9702
rect 11662 9591 11663 9617
rect 11689 9591 11690 9617
rect 11662 9585 11690 9591
rect 11606 9417 11634 9422
rect 11410 9254 11578 9282
rect 11382 9249 11410 9254
rect 11718 8834 11746 10654
rect 11886 10345 11914 11551
rect 12614 11241 12642 11887
rect 12838 11914 12866 11919
rect 12838 11867 12866 11886
rect 13174 11858 13202 13062
rect 13342 13057 13370 13062
rect 14014 12809 14042 13118
rect 18830 13146 18858 13151
rect 18830 13099 18858 13118
rect 20006 13033 20034 13039
rect 20006 13007 20007 13033
rect 20033 13007 20034 13033
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 14014 12783 14015 12809
rect 14041 12783 14042 12809
rect 14014 12777 14042 12783
rect 20006 12810 20034 13007
rect 20006 12777 20034 12782
rect 13342 12642 13370 12647
rect 13174 11825 13202 11830
rect 13230 12305 13258 12311
rect 13230 12279 13231 12305
rect 13257 12279 13258 12305
rect 13230 11857 13258 12279
rect 13286 11914 13314 11919
rect 13286 11867 13314 11886
rect 13230 11831 13231 11857
rect 13257 11831 13258 11857
rect 13230 11825 13258 11831
rect 13006 11802 13034 11807
rect 12614 11215 12615 11241
rect 12641 11215 12642 11241
rect 12614 11209 12642 11215
rect 12950 11774 13006 11802
rect 12894 11186 12922 11191
rect 12950 11186 12978 11774
rect 13006 11769 13034 11774
rect 13342 11241 13370 12614
rect 14182 12362 14210 12367
rect 13734 12082 13762 12087
rect 13762 12054 13818 12082
rect 13734 12049 13762 12054
rect 13454 11998 13650 12026
rect 13398 11970 13426 11975
rect 13454 11970 13482 11998
rect 13398 11969 13482 11970
rect 13398 11943 13399 11969
rect 13425 11943 13482 11969
rect 13398 11942 13482 11943
rect 13622 11969 13650 11998
rect 13622 11943 13623 11969
rect 13649 11943 13650 11969
rect 13398 11937 13426 11942
rect 13622 11937 13650 11943
rect 13734 11970 13762 11975
rect 13734 11923 13762 11942
rect 13566 11914 13594 11919
rect 13454 11913 13594 11914
rect 13454 11887 13567 11913
rect 13593 11887 13594 11913
rect 13454 11886 13594 11887
rect 13398 11858 13426 11863
rect 13454 11858 13482 11886
rect 13566 11881 13594 11886
rect 13426 11830 13482 11858
rect 13398 11689 13426 11830
rect 13398 11663 13399 11689
rect 13425 11663 13426 11689
rect 13398 11657 13426 11663
rect 13342 11215 13343 11241
rect 13369 11215 13370 11241
rect 12894 11185 12978 11186
rect 12894 11159 12895 11185
rect 12921 11159 12978 11185
rect 12894 11158 12978 11159
rect 13006 11186 13034 11191
rect 11886 10319 11887 10345
rect 11913 10319 11914 10345
rect 11830 9730 11858 9735
rect 11830 9337 11858 9702
rect 11830 9311 11831 9337
rect 11857 9311 11858 9337
rect 11830 9305 11858 9311
rect 11718 8801 11746 8806
rect 11774 9225 11802 9231
rect 11774 9199 11775 9225
rect 11801 9199 11802 9225
rect 11774 8666 11802 9199
rect 11774 8633 11802 8638
rect 11438 8498 11466 8503
rect 11326 8050 11354 8055
rect 11326 8003 11354 8022
rect 11214 7967 11215 7993
rect 11241 7967 11242 7993
rect 11214 7961 11242 7967
rect 11270 7937 11298 7943
rect 11270 7911 11271 7937
rect 11297 7911 11298 7937
rect 11270 7882 11298 7911
rect 11046 7854 11298 7882
rect 11438 7769 11466 8470
rect 11886 8441 11914 10319
rect 12614 11073 12642 11079
rect 12726 11074 12754 11079
rect 12614 11047 12615 11073
rect 12641 11047 12642 11073
rect 12614 10794 12642 11047
rect 12334 9954 12362 9959
rect 12278 9953 12362 9954
rect 12278 9927 12335 9953
rect 12361 9927 12362 9953
rect 12278 9926 12362 9927
rect 11942 9786 11970 9791
rect 11942 9225 11970 9758
rect 12166 9618 12194 9623
rect 12278 9618 12306 9926
rect 12334 9921 12362 9926
rect 12390 9786 12418 9791
rect 12194 9590 12306 9618
rect 12334 9730 12362 9735
rect 12166 9571 12194 9590
rect 12166 9282 12194 9287
rect 12334 9282 12362 9702
rect 12166 9281 12362 9282
rect 12166 9255 12167 9281
rect 12193 9255 12362 9281
rect 12166 9254 12362 9255
rect 12166 9249 12194 9254
rect 11942 9199 11943 9225
rect 11969 9199 11970 9225
rect 11942 9193 11970 9199
rect 12110 9113 12138 9119
rect 12110 9087 12111 9113
rect 12137 9087 12138 9113
rect 12110 8778 12138 9087
rect 12166 8778 12194 8783
rect 12110 8777 12194 8778
rect 12110 8751 12167 8777
rect 12193 8751 12194 8777
rect 12110 8750 12194 8751
rect 12166 8666 12194 8750
rect 12166 8633 12194 8638
rect 11886 8415 11887 8441
rect 11913 8415 11914 8441
rect 11886 8409 11914 8415
rect 12390 8161 12418 9758
rect 12446 9674 12474 9679
rect 12446 9627 12474 9646
rect 12614 9394 12642 10766
rect 12670 11073 12754 11074
rect 12670 11047 12727 11073
rect 12753 11047 12754 11073
rect 12670 11046 12754 11047
rect 12670 9786 12698 11046
rect 12726 11041 12754 11046
rect 12726 10794 12754 10799
rect 12838 10794 12866 10799
rect 12726 10747 12754 10766
rect 12782 10793 12866 10794
rect 12782 10767 12839 10793
rect 12865 10767 12866 10793
rect 12782 10766 12866 10767
rect 12670 9753 12698 9758
rect 12726 10009 12754 10015
rect 12726 9983 12727 10009
rect 12753 9983 12754 10009
rect 12726 9730 12754 9983
rect 12782 9786 12810 10766
rect 12838 10761 12866 10766
rect 12838 10122 12866 10127
rect 12894 10122 12922 11158
rect 13006 11139 13034 11158
rect 13062 11074 13090 11079
rect 13174 11074 13202 11079
rect 13062 11027 13090 11046
rect 13118 11073 13202 11074
rect 13118 11047 13175 11073
rect 13201 11047 13202 11073
rect 13118 11046 13202 11047
rect 13062 10850 13090 10855
rect 13118 10850 13146 11046
rect 13174 11041 13202 11046
rect 13230 11074 13258 11079
rect 13062 10849 13146 10850
rect 13062 10823 13063 10849
rect 13089 10823 13146 10849
rect 13062 10822 13146 10823
rect 13062 10817 13090 10822
rect 12950 10794 12978 10799
rect 12950 10747 12978 10766
rect 13006 10682 13034 10687
rect 13006 10635 13034 10654
rect 12838 10121 12922 10122
rect 12838 10095 12839 10121
rect 12865 10095 12922 10121
rect 12838 10094 12922 10095
rect 12838 10089 12866 10094
rect 13230 10066 13258 11046
rect 13286 10794 13314 10799
rect 13342 10794 13370 11215
rect 13286 10793 13370 10794
rect 13286 10767 13287 10793
rect 13313 10767 13370 10793
rect 13286 10766 13370 10767
rect 13734 10794 13762 10799
rect 13286 10761 13314 10766
rect 13622 10738 13650 10743
rect 13622 10691 13650 10710
rect 13734 10401 13762 10766
rect 13734 10375 13735 10401
rect 13761 10375 13762 10401
rect 13734 10369 13762 10375
rect 13454 10346 13482 10351
rect 13454 10299 13482 10318
rect 13622 10289 13650 10295
rect 13622 10263 13623 10289
rect 13649 10263 13650 10289
rect 13286 10066 13314 10071
rect 13230 10065 13314 10066
rect 13230 10039 13287 10065
rect 13313 10039 13314 10065
rect 13230 10038 13314 10039
rect 13286 10033 13314 10038
rect 12838 10009 12866 10015
rect 12838 9983 12839 10009
rect 12865 9983 12866 10009
rect 12838 9898 12866 9983
rect 13006 10010 13034 10015
rect 13118 10010 13146 10015
rect 13006 10009 13118 10010
rect 13006 9983 13007 10009
rect 13033 9983 13118 10009
rect 13006 9982 13118 9983
rect 13006 9977 13034 9982
rect 12838 9865 12866 9870
rect 12782 9758 12922 9786
rect 12726 9697 12754 9702
rect 12838 9618 12866 9623
rect 12390 8135 12391 8161
rect 12417 8135 12418 8161
rect 12390 8129 12418 8135
rect 12502 9366 12642 9394
rect 12670 9617 12866 9618
rect 12670 9591 12839 9617
rect 12865 9591 12866 9617
rect 12670 9590 12866 9591
rect 12446 8106 12474 8111
rect 11438 7743 11439 7769
rect 11465 7743 11466 7769
rect 11214 7602 11242 7621
rect 10766 7546 10850 7574
rect 11214 7569 11242 7574
rect 11438 7574 11466 7743
rect 11494 7993 11522 7999
rect 11494 7967 11495 7993
rect 11521 7967 11522 7993
rect 11494 7658 11522 7967
rect 11494 7625 11522 7630
rect 12222 7937 12250 7943
rect 12222 7911 12223 7937
rect 12249 7911 12250 7937
rect 11886 7602 11914 7607
rect 11438 7546 11802 7574
rect 10654 7266 10682 7271
rect 10598 7265 10682 7266
rect 10598 7239 10655 7265
rect 10681 7239 10682 7265
rect 10598 7238 10682 7239
rect 10262 7219 10290 7238
rect 10654 7233 10682 7238
rect 10766 7266 10794 7271
rect 10822 7266 10850 7546
rect 10766 7265 10850 7266
rect 10766 7239 10767 7265
rect 10793 7239 10850 7265
rect 10766 7238 10850 7239
rect 10934 7266 10962 7271
rect 10766 7233 10794 7238
rect 10934 7219 10962 7238
rect 11214 7209 11242 7215
rect 11214 7183 11215 7209
rect 11241 7183 11242 7209
rect 10206 7153 10234 7159
rect 10206 7127 10207 7153
rect 10233 7127 10234 7153
rect 10206 7098 10234 7127
rect 10822 7153 10850 7159
rect 10822 7127 10823 7153
rect 10849 7127 10850 7153
rect 10822 7098 10850 7127
rect 10878 7154 10906 7159
rect 10878 7107 10906 7126
rect 11158 7154 11186 7159
rect 11158 7107 11186 7126
rect 10206 7070 10346 7098
rect 10206 6986 10234 6991
rect 10150 6958 10206 6986
rect 9422 6903 9423 6929
rect 9449 6903 9450 6929
rect 9422 6897 9450 6903
rect 9254 6873 9282 6879
rect 9254 6847 9255 6873
rect 9281 6847 9282 6873
rect 9254 6537 9282 6847
rect 10206 6873 10234 6958
rect 10206 6847 10207 6873
rect 10233 6847 10234 6873
rect 10206 6841 10234 6847
rect 9254 6511 9255 6537
rect 9281 6511 9282 6537
rect 9254 6505 9282 6511
rect 10318 6537 10346 7070
rect 10542 7070 10850 7098
rect 10542 6929 10570 7070
rect 10542 6903 10543 6929
rect 10569 6903 10570 6929
rect 10542 6897 10570 6903
rect 10766 6986 10794 6991
rect 10318 6511 10319 6537
rect 10345 6511 10346 6537
rect 8862 6455 8863 6481
rect 8889 6455 8890 6481
rect 8862 6449 8890 6455
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 10318 4214 10346 6511
rect 10766 6537 10794 6958
rect 11214 6762 11242 7183
rect 11774 6986 11802 7546
rect 11830 6986 11858 6991
rect 11774 6958 11830 6986
rect 11830 6939 11858 6958
rect 11214 6729 11242 6734
rect 11606 6817 11634 6823
rect 11606 6791 11607 6817
rect 11633 6791 11634 6817
rect 11606 6762 11634 6791
rect 11606 6729 11634 6734
rect 10766 6511 10767 6537
rect 10793 6511 10794 6537
rect 10766 6505 10794 6511
rect 11886 4214 11914 7574
rect 12222 7574 12250 7911
rect 12222 7546 12362 7574
rect 12334 7265 12362 7546
rect 12334 7239 12335 7265
rect 12361 7239 12362 7265
rect 12334 7233 12362 7239
rect 12446 7265 12474 8078
rect 12502 8105 12530 9366
rect 12670 9338 12698 9590
rect 12838 9585 12866 9590
rect 12894 9450 12922 9758
rect 12894 9417 12922 9422
rect 12614 9337 12698 9338
rect 12614 9311 12671 9337
rect 12697 9311 12698 9337
rect 12614 9310 12698 9311
rect 12558 8834 12586 8839
rect 12614 8834 12642 9310
rect 12670 9305 12698 9310
rect 13118 9282 13146 9982
rect 13174 10009 13202 10015
rect 13174 9983 13175 10009
rect 13201 9983 13202 10009
rect 13174 9898 13202 9983
rect 13510 10009 13538 10015
rect 13510 9983 13511 10009
rect 13537 9983 13538 10009
rect 13230 9954 13258 9959
rect 13230 9953 13426 9954
rect 13230 9927 13231 9953
rect 13257 9927 13426 9953
rect 13230 9926 13426 9927
rect 13230 9921 13258 9926
rect 13174 9865 13202 9870
rect 13230 9562 13258 9567
rect 13230 9561 13370 9562
rect 13230 9535 13231 9561
rect 13257 9535 13370 9561
rect 13230 9534 13370 9535
rect 13230 9529 13258 9534
rect 13118 9249 13146 9254
rect 13286 9450 13314 9455
rect 13286 9281 13314 9422
rect 13342 9337 13370 9534
rect 13342 9311 13343 9337
rect 13369 9311 13370 9337
rect 13342 9305 13370 9311
rect 13286 9255 13287 9281
rect 13313 9255 13314 9281
rect 13286 9249 13314 9255
rect 13398 9282 13426 9926
rect 13510 9618 13538 9983
rect 13622 10010 13650 10263
rect 13622 9977 13650 9982
rect 13510 9585 13538 9590
rect 13622 9898 13650 9903
rect 13398 9254 13482 9282
rect 13174 9226 13202 9231
rect 13174 9179 13202 9198
rect 13342 9226 13370 9231
rect 12558 8833 12642 8834
rect 12558 8807 12559 8833
rect 12585 8807 12642 8833
rect 12558 8806 12642 8807
rect 12558 8801 12586 8806
rect 12502 8079 12503 8105
rect 12529 8079 12530 8105
rect 12502 7770 12530 8079
rect 12614 8554 12642 8806
rect 12614 7770 12642 8526
rect 13118 8554 13146 8559
rect 13146 8526 13314 8554
rect 13118 8507 13146 8526
rect 13286 8441 13314 8526
rect 13286 8415 13287 8441
rect 13313 8415 13314 8441
rect 13286 8409 13314 8415
rect 13286 8050 13314 8055
rect 13342 8050 13370 9198
rect 13454 9225 13482 9254
rect 13622 9281 13650 9870
rect 13734 9338 13762 9343
rect 13790 9338 13818 12054
rect 14070 11970 14098 11975
rect 14070 11923 14098 11942
rect 13846 11914 13874 11919
rect 13846 11867 13874 11886
rect 14182 11913 14210 12334
rect 18830 12362 18858 12367
rect 18830 12315 18858 12334
rect 14294 12305 14322 12311
rect 14294 12279 14295 12305
rect 14321 12279 14322 12305
rect 14294 11970 14322 12279
rect 20006 12249 20034 12255
rect 20006 12223 20007 12249
rect 20033 12223 20034 12249
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 20006 12138 20034 12223
rect 20006 12105 20034 12110
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 14294 11937 14322 11942
rect 18830 11970 18858 11975
rect 18830 11923 18858 11942
rect 14182 11887 14183 11913
rect 14209 11887 14210 11913
rect 14182 11881 14210 11887
rect 20006 11802 20034 11999
rect 20006 11769 20034 11774
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 20118 11073 20146 11079
rect 20118 11047 20119 11073
rect 20145 11047 20146 11073
rect 13846 10794 13874 10799
rect 13846 10345 13874 10766
rect 14686 10794 14714 10799
rect 14686 10737 14714 10766
rect 18830 10794 18858 10799
rect 18830 10747 18858 10766
rect 20118 10794 20146 11047
rect 20118 10761 20146 10766
rect 14686 10711 14687 10737
rect 14713 10711 14714 10737
rect 14686 10705 14714 10711
rect 20006 10681 20034 10687
rect 20006 10655 20007 10681
rect 20033 10655 20034 10681
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 20006 10458 20034 10655
rect 20006 10425 20034 10430
rect 13846 10319 13847 10345
rect 13873 10319 13874 10345
rect 13846 10313 13874 10319
rect 13902 10345 13930 10351
rect 13902 10319 13903 10345
rect 13929 10319 13930 10345
rect 13902 10010 13930 10319
rect 13902 9977 13930 9982
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 14294 9673 14322 9679
rect 14294 9647 14295 9673
rect 14321 9647 14322 9673
rect 14294 9618 14322 9647
rect 20006 9673 20034 9679
rect 20006 9647 20007 9673
rect 20033 9647 20034 9673
rect 14294 9585 14322 9590
rect 18830 9618 18858 9623
rect 18830 9571 18858 9590
rect 20006 9450 20034 9647
rect 20006 9417 20034 9422
rect 13734 9337 13818 9338
rect 13734 9311 13735 9337
rect 13761 9311 13818 9337
rect 13734 9310 13818 9311
rect 13734 9305 13762 9310
rect 13622 9255 13623 9281
rect 13649 9255 13650 9281
rect 13622 9249 13650 9255
rect 13454 9199 13455 9225
rect 13481 9199 13482 9225
rect 13454 9193 13482 9199
rect 13678 9226 13706 9231
rect 13678 9179 13706 9198
rect 13790 9058 13818 9310
rect 14126 9338 14154 9343
rect 14126 9291 14154 9310
rect 14742 9338 14770 9343
rect 14070 9282 14098 9287
rect 14070 9235 14098 9254
rect 13958 9225 13986 9231
rect 13958 9199 13959 9225
rect 13985 9199 13986 9225
rect 13958 9114 13986 9199
rect 14126 9114 14154 9119
rect 13958 9113 14154 9114
rect 13958 9087 14127 9113
rect 14153 9087 14154 9113
rect 13958 9086 14154 9087
rect 14126 9081 14154 9086
rect 13510 9030 13818 9058
rect 13510 8889 13538 9030
rect 13510 8863 13511 8889
rect 13537 8863 13538 8889
rect 13510 8857 13538 8863
rect 14742 8834 14770 9310
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 13678 8498 13706 8503
rect 13678 8451 13706 8470
rect 14742 8385 14770 8806
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 14742 8359 14743 8385
rect 14769 8359 14770 8385
rect 14742 8353 14770 8359
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 13286 8049 13370 8050
rect 13286 8023 13287 8049
rect 13313 8023 13370 8049
rect 13286 8022 13370 8023
rect 13286 8017 13314 8022
rect 13118 7938 13146 7943
rect 13006 7937 13146 7938
rect 13006 7911 13119 7937
rect 13145 7911 13146 7937
rect 13006 7910 13146 7911
rect 12670 7770 12698 7775
rect 12614 7769 12698 7770
rect 12614 7743 12671 7769
rect 12697 7743 12698 7769
rect 12614 7742 12698 7743
rect 12502 7737 12530 7742
rect 12446 7239 12447 7265
rect 12473 7239 12474 7265
rect 12446 7233 12474 7239
rect 12558 7658 12586 7663
rect 12558 7265 12586 7630
rect 12670 7574 12698 7742
rect 13006 7714 13034 7910
rect 13118 7905 13146 7910
rect 13342 7770 13370 7775
rect 13342 7723 13370 7742
rect 13622 7769 13650 7775
rect 13622 7743 13623 7769
rect 13649 7743 13650 7769
rect 12670 7546 12866 7574
rect 12558 7239 12559 7265
rect 12585 7239 12586 7265
rect 12558 7233 12586 7239
rect 12614 7266 12642 7271
rect 12614 7219 12642 7238
rect 12502 7154 12530 7159
rect 12502 7107 12530 7126
rect 12334 6986 12362 6991
rect 12334 6939 12362 6958
rect 12670 6986 12698 7546
rect 12838 7265 12866 7546
rect 12838 7239 12839 7265
rect 12865 7239 12866 7265
rect 12838 7233 12866 7239
rect 13006 7266 13034 7686
rect 13566 7714 13594 7719
rect 13622 7714 13650 7743
rect 13678 7714 13706 7719
rect 13622 7686 13678 7714
rect 13566 7667 13594 7686
rect 13678 7681 13706 7686
rect 13062 7658 13090 7663
rect 13062 7601 13090 7630
rect 13230 7657 13258 7663
rect 13230 7631 13231 7657
rect 13257 7631 13258 7657
rect 13062 7575 13063 7601
rect 13089 7575 13090 7601
rect 13062 7569 13090 7575
rect 13118 7602 13146 7621
rect 13118 7569 13146 7574
rect 13230 7321 13258 7631
rect 13398 7658 13426 7663
rect 13398 7611 13426 7630
rect 13734 7658 13762 7663
rect 13734 7611 13762 7630
rect 14294 7658 14322 7663
rect 13230 7295 13231 7321
rect 13257 7295 13258 7321
rect 13230 7289 13258 7295
rect 14070 7602 14098 7607
rect 13006 7233 13034 7238
rect 12670 6873 12698 6958
rect 13006 7154 13034 7159
rect 13006 6929 13034 7126
rect 13006 6903 13007 6929
rect 13033 6903 13034 6929
rect 13006 6897 13034 6903
rect 12670 6847 12671 6873
rect 12697 6847 12698 6873
rect 12670 6841 12698 6847
rect 14070 6817 14098 7574
rect 14294 7321 14322 7630
rect 18830 7658 18858 7663
rect 18830 7611 18858 7630
rect 20006 7601 20034 7607
rect 20006 7575 20007 7601
rect 20033 7575 20034 7601
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 20006 7434 20034 7575
rect 20006 7401 20034 7406
rect 14294 7295 14295 7321
rect 14321 7295 14322 7321
rect 14294 7289 14322 7295
rect 14070 6791 14071 6817
rect 14097 6791 14098 6817
rect 10318 4186 10570 4214
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 10542 2169 10570 4186
rect 10542 2143 10543 2169
rect 10569 2143 10570 2169
rect 10542 2137 10570 2143
rect 11774 4186 11914 4214
rect 12278 6762 12306 6767
rect 14070 6762 14098 6791
rect 14070 6734 14322 6762
rect 8470 1751 8471 1777
rect 8497 1751 8498 1777
rect 8470 1745 8498 1751
rect 10430 2058 10458 2063
rect 8078 1722 8106 1727
rect 7182 1666 7210 1671
rect 7070 1665 7210 1666
rect 7070 1639 7183 1665
rect 7209 1639 7210 1665
rect 7070 1638 7210 1639
rect 7070 400 7098 1638
rect 7182 1633 7210 1638
rect 8078 400 8106 1694
rect 9254 1722 9282 1727
rect 9254 1675 9282 1694
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10430 400 10458 2030
rect 11046 2058 11074 2063
rect 11046 2011 11074 2030
rect 10822 1834 10850 1839
rect 10766 1833 10850 1834
rect 10766 1807 10823 1833
rect 10849 1807 10850 1833
rect 10766 1806 10850 1807
rect 10766 400 10794 1806
rect 10822 1801 10850 1806
rect 11438 1834 11466 1839
rect 11438 400 11466 1806
rect 11774 1777 11802 4186
rect 11774 1751 11775 1777
rect 11801 1751 11802 1777
rect 11774 1745 11802 1751
rect 12278 1777 12306 6734
rect 14294 2169 14322 6734
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 14294 2143 14295 2169
rect 14321 2143 14322 2169
rect 14294 2137 14322 2143
rect 13342 2058 13370 2063
rect 13118 2057 13370 2058
rect 13118 2031 13343 2057
rect 13369 2031 13370 2057
rect 13118 2030 13370 2031
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1745 12306 1751
rect 13118 400 13146 2030
rect 13342 2025 13370 2030
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 14238 1666 14266 1671
rect 14126 1665 14266 1666
rect 14126 1639 14239 1665
rect 14265 1639 14266 1665
rect 14126 1638 14266 1639
rect 14126 400 14154 1638
rect 14238 1633 14266 1638
rect 7056 0 7112 400
rect 8064 0 8120 400
rect 10416 0 10472 400
rect 10752 0 10808 400
rect 11424 0 11480 400
rect 13104 0 13160 400
rect 14112 0 14168 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 8414 19110 8442 19138
rect 9030 19137 9058 19138
rect 9030 19111 9031 19137
rect 9031 19111 9057 19137
rect 9057 19111 9058 19137
rect 9030 19110 9058 19111
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 12110 19110 12138 19138
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 10766 18718 10794 18746
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 7350 13790 7378 13818
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 7910 13817 7938 13818
rect 7910 13791 7911 13817
rect 7911 13791 7937 13817
rect 7937 13791 7938 13817
rect 7910 13790 7938 13791
rect 966 13118 994 13146
rect 2086 13454 2114 13482
rect 966 12782 994 12810
rect 966 11241 994 11242
rect 966 11215 967 11241
rect 967 11215 993 11241
rect 993 11215 994 11241
rect 966 11214 994 11215
rect 2142 13230 2170 13258
rect 5782 13230 5810 13258
rect 2142 13145 2170 13146
rect 2142 13119 2143 13145
rect 2143 13119 2169 13145
rect 2169 13119 2170 13145
rect 2142 13118 2170 13119
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 5782 12670 5810 12698
rect 6062 13118 6090 13146
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 7518 13062 7546 13090
rect 7350 12753 7378 12754
rect 7350 12727 7351 12753
rect 7351 12727 7377 12753
rect 7377 12727 7378 12753
rect 7350 12726 7378 12727
rect 6062 12614 6090 12642
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 6790 11662 6818 11690
rect 6678 11438 6706 11466
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 2142 11185 2170 11186
rect 2142 11159 2143 11185
rect 2143 11159 2169 11185
rect 2169 11159 2170 11185
rect 2142 11158 2170 11159
rect 5614 11158 5642 11186
rect 2142 10793 2170 10794
rect 2142 10767 2143 10793
rect 2143 10767 2169 10793
rect 2169 10767 2170 10793
rect 2142 10766 2170 10767
rect 4998 10766 5026 10794
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 2086 10486 2114 10514
rect 966 10430 994 10458
rect 6062 10710 6090 10738
rect 4998 10457 5026 10458
rect 4998 10431 4999 10457
rect 4999 10431 5025 10457
rect 5025 10431 5026 10457
rect 4998 10430 5026 10431
rect 7294 12697 7322 12698
rect 7294 12671 7295 12697
rect 7295 12671 7321 12697
rect 7321 12671 7322 12697
rect 7294 12670 7322 12671
rect 8134 12782 8162 12810
rect 7518 12753 7546 12754
rect 7518 12727 7519 12753
rect 7519 12727 7545 12753
rect 7545 12727 7546 12753
rect 7518 12726 7546 12727
rect 7798 12670 7826 12698
rect 7574 12641 7602 12642
rect 7574 12615 7575 12641
rect 7575 12615 7601 12641
rect 7601 12615 7602 12641
rect 7574 12614 7602 12615
rect 7126 12305 7154 12306
rect 7126 12279 7127 12305
rect 7127 12279 7153 12305
rect 7153 12279 7154 12305
rect 7126 12278 7154 12279
rect 7630 11662 7658 11690
rect 7182 11550 7210 11578
rect 7126 11465 7154 11466
rect 7126 11439 7127 11465
rect 7127 11439 7153 11465
rect 7153 11439 7154 11465
rect 7126 11438 7154 11439
rect 7126 10878 7154 10906
rect 7350 11102 7378 11130
rect 7070 10822 7098 10850
rect 7742 11577 7770 11578
rect 7742 11551 7743 11577
rect 7743 11551 7769 11577
rect 7769 11551 7770 11577
rect 7742 11550 7770 11551
rect 8414 13145 8442 13146
rect 8414 13119 8415 13145
rect 8415 13119 8441 13145
rect 8441 13119 8442 13145
rect 8414 13118 8442 13119
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 8750 13089 8778 13090
rect 8750 13063 8751 13089
rect 8751 13063 8777 13089
rect 8777 13063 8778 13089
rect 8750 13062 8778 13063
rect 9142 12782 9170 12810
rect 8414 12726 8442 12754
rect 8190 12670 8218 12698
rect 9198 12614 9226 12642
rect 9366 13145 9394 13146
rect 9366 13119 9367 13145
rect 9367 13119 9393 13145
rect 9393 13119 9394 13145
rect 9366 13118 9394 13119
rect 9590 13062 9618 13090
rect 11382 18745 11410 18746
rect 11382 18719 11383 18745
rect 11383 18719 11409 18745
rect 11409 18719 11410 18745
rect 11382 18718 11410 18719
rect 10262 13062 10290 13090
rect 10934 13062 10962 13090
rect 10654 12782 10682 12810
rect 9646 12697 9674 12698
rect 9646 12671 9647 12697
rect 9647 12671 9673 12697
rect 9673 12671 9674 12697
rect 9646 12670 9674 12671
rect 9758 12641 9786 12642
rect 9758 12615 9759 12641
rect 9759 12615 9785 12641
rect 9785 12615 9786 12641
rect 9758 12614 9786 12615
rect 7686 11214 7714 11242
rect 7574 11158 7602 11186
rect 7742 11046 7770 11074
rect 7294 10737 7322 10738
rect 7294 10711 7295 10737
rect 7295 10711 7321 10737
rect 7321 10711 7322 10737
rect 7294 10710 7322 10711
rect 7406 10710 7434 10738
rect 6454 10401 6482 10402
rect 6454 10375 6455 10401
rect 6455 10375 6481 10401
rect 6481 10375 6482 10401
rect 6454 10374 6482 10375
rect 6958 10457 6986 10458
rect 6958 10431 6959 10457
rect 6959 10431 6985 10457
rect 6985 10431 6986 10457
rect 6958 10430 6986 10431
rect 6790 10374 6818 10402
rect 7238 10401 7266 10402
rect 7238 10375 7239 10401
rect 7239 10375 7265 10401
rect 7265 10375 7266 10401
rect 7238 10374 7266 10375
rect 7518 10822 7546 10850
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 7238 9646 7266 9674
rect 966 9422 994 9450
rect 6678 9478 6706 9506
rect 2142 9142 2170 9170
rect 5614 9169 5642 9170
rect 5614 9143 5615 9169
rect 5615 9143 5641 9169
rect 5641 9143 5642 9169
rect 5614 9142 5642 9143
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 7574 10038 7602 10066
rect 7574 9926 7602 9954
rect 7294 9505 7322 9506
rect 7294 9479 7295 9505
rect 7295 9479 7321 9505
rect 7321 9479 7322 9505
rect 7294 9478 7322 9479
rect 7742 10934 7770 10962
rect 7742 9926 7770 9954
rect 7854 12361 7882 12362
rect 7854 12335 7855 12361
rect 7855 12335 7881 12361
rect 7881 12335 7882 12361
rect 7854 12334 7882 12335
rect 7910 12305 7938 12306
rect 7910 12279 7911 12305
rect 7911 12279 7937 12305
rect 7937 12279 7938 12305
rect 7910 12278 7938 12279
rect 7910 10849 7938 10850
rect 7910 10823 7911 10849
rect 7911 10823 7937 10849
rect 7937 10823 7938 10849
rect 7910 10822 7938 10823
rect 7854 10710 7882 10738
rect 8190 12054 8218 12082
rect 8358 11886 8386 11914
rect 8302 11521 8330 11522
rect 8302 11495 8303 11521
rect 8303 11495 8329 11521
rect 8329 11495 8330 11521
rect 8302 11494 8330 11495
rect 8022 11046 8050 11074
rect 8414 11241 8442 11242
rect 8414 11215 8415 11241
rect 8415 11215 8441 11241
rect 8441 11215 8442 11241
rect 8414 11214 8442 11215
rect 8638 11185 8666 11186
rect 8638 11159 8639 11185
rect 8639 11159 8665 11185
rect 8665 11159 8666 11185
rect 8638 11158 8666 11159
rect 8190 11102 8218 11130
rect 8022 10934 8050 10962
rect 8078 10905 8106 10906
rect 8078 10879 8079 10905
rect 8079 10879 8105 10905
rect 8105 10879 8106 10905
rect 8078 10878 8106 10879
rect 7966 10430 7994 10458
rect 8470 11073 8498 11074
rect 8470 11047 8471 11073
rect 8471 11047 8497 11073
rect 8497 11047 8498 11073
rect 8470 11046 8498 11047
rect 8694 10934 8722 10962
rect 9198 11774 9226 11802
rect 9086 11633 9114 11634
rect 9086 11607 9087 11633
rect 9087 11607 9113 11633
rect 9113 11607 9114 11633
rect 9086 11606 9114 11607
rect 8862 11297 8890 11298
rect 8862 11271 8863 11297
rect 8863 11271 8889 11297
rect 8889 11271 8890 11297
rect 8862 11270 8890 11271
rect 8806 11214 8834 11242
rect 8806 11129 8834 11130
rect 8806 11103 8807 11129
rect 8807 11103 8833 11129
rect 8833 11103 8834 11129
rect 8806 11102 8834 11103
rect 9086 11102 9114 11130
rect 8750 10822 8778 10850
rect 8414 10094 8442 10122
rect 8078 10065 8106 10066
rect 8078 10039 8079 10065
rect 8079 10039 8105 10065
rect 8105 10039 8106 10065
rect 8078 10038 8106 10039
rect 7854 9926 7882 9954
rect 7686 9673 7714 9674
rect 7686 9647 7687 9673
rect 7687 9647 7713 9673
rect 7713 9647 7714 9673
rect 7686 9646 7714 9647
rect 7574 9310 7602 9338
rect 7238 9142 7266 9170
rect 7070 8862 7098 8890
rect 5614 8750 5642 8778
rect 7182 8777 7210 8778
rect 7182 8751 7183 8777
rect 7183 8751 7209 8777
rect 7209 8751 7210 8777
rect 7182 8750 7210 8751
rect 7630 9366 7658 9394
rect 8134 10009 8162 10010
rect 8134 9983 8135 10009
rect 8135 9983 8161 10009
rect 8161 9983 8162 10009
rect 8134 9982 8162 9983
rect 8918 10094 8946 10122
rect 9590 11969 9618 11970
rect 9590 11943 9591 11969
rect 9591 11943 9617 11969
rect 9617 11943 9618 11969
rect 9590 11942 9618 11943
rect 9366 11774 9394 11802
rect 9422 11606 9450 11634
rect 9310 11270 9338 11298
rect 9422 11158 9450 11186
rect 9254 10318 9282 10346
rect 7686 9281 7714 9282
rect 7686 9255 7687 9281
rect 7687 9255 7713 9281
rect 7713 9255 7714 9281
rect 7686 9254 7714 9255
rect 7350 8862 7378 8890
rect 7238 8553 7266 8554
rect 7238 8527 7239 8553
rect 7239 8527 7265 8553
rect 7265 8527 7266 8553
rect 7238 8526 7266 8527
rect 2142 8441 2170 8442
rect 2142 8415 2143 8441
rect 2143 8415 2169 8441
rect 2169 8415 2170 8441
rect 2142 8414 2170 8415
rect 5950 8414 5978 8442
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 966 8078 994 8106
rect 7126 8358 7154 8386
rect 7910 9366 7938 9394
rect 7798 8862 7826 8890
rect 8414 9478 8442 9506
rect 8078 9422 8106 9450
rect 8022 9086 8050 9114
rect 8246 9142 8274 9170
rect 7966 8974 7994 9002
rect 7742 8750 7770 8778
rect 7630 8497 7658 8498
rect 7630 8471 7631 8497
rect 7631 8471 7657 8497
rect 7657 8471 7658 8497
rect 7630 8470 7658 8471
rect 7574 8385 7602 8386
rect 7574 8359 7575 8385
rect 7575 8359 7601 8385
rect 7601 8359 7602 8385
rect 7574 8358 7602 8359
rect 7630 7713 7658 7714
rect 7630 7687 7631 7713
rect 7631 7687 7657 7713
rect 7657 7687 7658 7713
rect 7630 7686 7658 7687
rect 7462 7574 7490 7602
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 8246 8862 8274 8890
rect 8414 9198 8442 9226
rect 8246 8777 8274 8778
rect 8246 8751 8247 8777
rect 8247 8751 8273 8777
rect 8273 8751 8274 8777
rect 8246 8750 8274 8751
rect 8022 8078 8050 8106
rect 8918 9982 8946 10010
rect 8974 9729 9002 9730
rect 8974 9703 8975 9729
rect 8975 9703 9001 9729
rect 9001 9703 9002 9729
rect 8974 9702 9002 9703
rect 9254 9926 9282 9954
rect 9702 11185 9730 11186
rect 9702 11159 9703 11185
rect 9703 11159 9729 11185
rect 9729 11159 9730 11185
rect 9702 11158 9730 11159
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 10150 12334 10178 12362
rect 9982 11886 10010 11914
rect 10374 12305 10402 12306
rect 10374 12279 10375 12305
rect 10375 12279 10401 12305
rect 10401 12279 10402 12305
rect 10374 12278 10402 12279
rect 10374 11998 10402 12026
rect 10206 11857 10234 11858
rect 10206 11831 10207 11857
rect 10207 11831 10233 11857
rect 10233 11831 10234 11857
rect 10206 11830 10234 11831
rect 10374 11913 10402 11914
rect 10374 11887 10375 11913
rect 10375 11887 10401 11913
rect 10401 11887 10402 11913
rect 10374 11886 10402 11887
rect 9814 11774 9842 11802
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 10094 11521 10122 11522
rect 10094 11495 10095 11521
rect 10095 11495 10121 11521
rect 10121 11495 10122 11521
rect 10094 11494 10122 11495
rect 9814 11158 9842 11186
rect 9982 11185 10010 11186
rect 9982 11159 9983 11185
rect 9983 11159 10009 11185
rect 10009 11159 10010 11185
rect 9982 11158 10010 11159
rect 9926 11102 9954 11130
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 9926 10878 9954 10906
rect 9590 10737 9618 10738
rect 9590 10711 9591 10737
rect 9591 10711 9617 10737
rect 9617 10711 9618 10737
rect 9590 10710 9618 10711
rect 9422 9953 9450 9954
rect 9422 9927 9423 9953
rect 9423 9927 9449 9953
rect 9449 9927 9450 9953
rect 9422 9926 9450 9927
rect 9310 9646 9338 9674
rect 8862 9198 8890 9226
rect 8918 9310 8946 9338
rect 9142 9310 9170 9338
rect 9030 9225 9058 9226
rect 9030 9199 9031 9225
rect 9031 9199 9057 9225
rect 9057 9199 9058 9225
rect 9030 9198 9058 9199
rect 9870 10793 9898 10794
rect 9870 10767 9871 10793
rect 9871 10767 9897 10793
rect 9897 10767 9898 10793
rect 9870 10766 9898 10767
rect 9702 10486 9730 10514
rect 9870 10457 9898 10458
rect 9870 10431 9871 10457
rect 9871 10431 9897 10457
rect 9897 10431 9898 10457
rect 9870 10430 9898 10431
rect 9814 10374 9842 10402
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 10150 10934 10178 10962
rect 10038 10009 10066 10010
rect 10038 9983 10039 10009
rect 10039 9983 10065 10009
rect 10065 9983 10066 10009
rect 10038 9982 10066 9983
rect 10150 10822 10178 10850
rect 10430 11102 10458 11130
rect 10206 10766 10234 10794
rect 10262 10934 10290 10962
rect 10150 10374 10178 10402
rect 9646 9590 9674 9618
rect 9366 9561 9394 9562
rect 9366 9535 9367 9561
rect 9367 9535 9393 9561
rect 9393 9535 9394 9561
rect 9366 9534 9394 9535
rect 9310 9254 9338 9282
rect 9814 9702 9842 9730
rect 10374 10878 10402 10906
rect 10710 12697 10738 12698
rect 10710 12671 10711 12697
rect 10711 12671 10737 12697
rect 10737 12671 10738 12697
rect 10710 12670 10738 12671
rect 10598 11046 10626 11074
rect 10542 10766 10570 10794
rect 10654 10990 10682 11018
rect 11270 13089 11298 13090
rect 11270 13063 11271 13089
rect 11271 13063 11297 13089
rect 11297 13063 11298 13089
rect 11270 13062 11298 13063
rect 11494 13089 11522 13090
rect 11494 13063 11495 13089
rect 11495 13063 11521 13089
rect 11521 13063 11522 13089
rect 11494 13062 11522 13063
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 13062 13201 13090 13202
rect 13062 13175 13063 13201
rect 13063 13175 13089 13201
rect 13089 13175 13090 13201
rect 13062 13174 13090 13175
rect 11046 12670 11074 12698
rect 12614 13062 12642 13090
rect 14014 13118 14042 13146
rect 12670 12614 12698 12642
rect 11102 12278 11130 12306
rect 11214 12081 11242 12082
rect 11214 12055 11215 12081
rect 11215 12055 11241 12081
rect 11241 12055 11242 12081
rect 11214 12054 11242 12055
rect 10766 11830 10794 11858
rect 10598 10710 10626 10738
rect 10206 9870 10234 9898
rect 9702 9561 9730 9562
rect 9702 9535 9703 9561
rect 9703 9535 9729 9561
rect 9729 9535 9730 9561
rect 9702 9534 9730 9535
rect 9646 9310 9674 9338
rect 9254 9142 9282 9170
rect 9590 9142 9618 9170
rect 9758 9281 9786 9282
rect 9758 9255 9759 9281
rect 9759 9255 9785 9281
rect 9785 9255 9786 9281
rect 9758 9254 9786 9255
rect 9702 9198 9730 9226
rect 9534 9086 9562 9114
rect 8862 8806 8890 8834
rect 9366 8833 9394 8834
rect 9366 8807 9367 8833
rect 9367 8807 9393 8833
rect 9393 8807 9394 8833
rect 9366 8806 9394 8807
rect 9926 9646 9954 9674
rect 10094 9646 10122 9674
rect 9982 9617 10010 9618
rect 9982 9591 9983 9617
rect 9983 9591 10009 9617
rect 10009 9591 10010 9617
rect 9982 9590 10010 9591
rect 10654 9926 10682 9954
rect 10318 9590 10346 9618
rect 10094 9505 10122 9506
rect 10094 9479 10095 9505
rect 10095 9479 10121 9505
rect 10121 9479 10122 9505
rect 10094 9478 10122 9479
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 10318 9254 10346 9282
rect 10430 9646 10458 9674
rect 10878 11998 10906 12026
rect 11550 11969 11578 11970
rect 11550 11943 11551 11969
rect 11551 11943 11577 11969
rect 11577 11943 11578 11969
rect 11550 11942 11578 11943
rect 11270 11913 11298 11914
rect 11270 11887 11271 11913
rect 11271 11887 11297 11913
rect 11297 11887 11298 11913
rect 11270 11886 11298 11887
rect 10822 10934 10850 10962
rect 11438 11857 11466 11858
rect 11438 11831 11439 11857
rect 11439 11831 11465 11857
rect 11465 11831 11466 11857
rect 11438 11830 11466 11831
rect 11662 11158 11690 11186
rect 11046 11046 11074 11074
rect 11214 10934 11242 10962
rect 11830 11942 11858 11970
rect 12726 12166 12754 12194
rect 12950 12222 12978 12250
rect 13062 12166 13090 12194
rect 11550 11073 11578 11074
rect 11550 11047 11551 11073
rect 11551 11047 11577 11073
rect 11577 11047 11578 11073
rect 11550 11046 11578 11047
rect 10878 10878 10906 10906
rect 10822 10849 10850 10850
rect 10822 10823 10823 10849
rect 10823 10823 10849 10849
rect 10849 10823 10850 10849
rect 10822 10822 10850 10823
rect 11158 10822 11186 10850
rect 10934 10486 10962 10514
rect 10878 10009 10906 10010
rect 10878 9983 10879 10009
rect 10879 9983 10905 10009
rect 10905 9983 10906 10009
rect 10878 9982 10906 9983
rect 10766 9758 10794 9786
rect 10934 9870 10962 9898
rect 10710 9646 10738 9674
rect 11102 9646 11130 9674
rect 10710 9478 10738 9506
rect 10430 9198 10458 9226
rect 10486 9254 10514 9282
rect 11046 9198 11074 9226
rect 10038 9113 10066 9114
rect 10038 9087 10039 9113
rect 10039 9087 10065 9113
rect 10065 9087 10066 9113
rect 10038 9086 10066 9087
rect 10038 8974 10066 9002
rect 10262 8833 10290 8834
rect 10262 8807 10263 8833
rect 10263 8807 10289 8833
rect 10289 8807 10290 8833
rect 10262 8806 10290 8807
rect 9310 8694 9338 8722
rect 9702 8721 9730 8722
rect 9702 8695 9703 8721
rect 9703 8695 9729 8721
rect 9729 8695 9730 8721
rect 9702 8694 9730 8695
rect 10318 8721 10346 8722
rect 10318 8695 10319 8721
rect 10319 8695 10345 8721
rect 10345 8695 10346 8721
rect 10318 8694 10346 8695
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10150 8638 10178 8666
rect 10022 8610 10050 8611
rect 9142 8078 9170 8106
rect 10374 8022 10402 8050
rect 8806 7769 8834 7770
rect 8806 7743 8807 7769
rect 8807 7743 8833 7769
rect 8833 7743 8834 7769
rect 8806 7742 8834 7743
rect 8078 7686 8106 7714
rect 7854 7601 7882 7602
rect 7854 7575 7855 7601
rect 7855 7575 7881 7601
rect 7881 7575 7882 7601
rect 7854 7574 7882 7575
rect 6678 7126 6706 7154
rect 7518 7153 7546 7154
rect 7518 7127 7519 7153
rect 7519 7127 7545 7153
rect 7545 7127 7546 7153
rect 7518 7126 7546 7127
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 10262 7686 10290 7714
rect 8470 7126 8498 7154
rect 8414 6958 8442 6986
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9478 7630 9506 7658
rect 9758 7657 9786 7658
rect 9758 7631 9759 7657
rect 9759 7631 9785 7657
rect 9785 7631 9786 7657
rect 9758 7630 9786 7631
rect 10094 7630 10122 7658
rect 9030 7070 9058 7098
rect 8862 6958 8890 6986
rect 9422 7126 9450 7154
rect 9198 6958 9226 6986
rect 9366 7070 9394 7098
rect 10094 7153 10122 7154
rect 10094 7127 10095 7153
rect 10095 7127 10121 7153
rect 10121 7127 10122 7153
rect 10094 7126 10122 7127
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 10262 7265 10290 7266
rect 10262 7239 10263 7265
rect 10263 7239 10289 7265
rect 10289 7239 10290 7265
rect 10262 7238 10290 7239
rect 10654 8638 10682 8666
rect 10710 8526 10738 8554
rect 10710 7686 10738 7714
rect 10934 8497 10962 8498
rect 10934 8471 10935 8497
rect 10935 8471 10961 8497
rect 10961 8471 10962 8497
rect 10934 8470 10962 8471
rect 11102 9142 11130 9170
rect 11214 9534 11242 9562
rect 10822 8049 10850 8050
rect 10822 8023 10823 8049
rect 10823 8023 10849 8049
rect 10849 8023 10850 8049
rect 10822 8022 10850 8023
rect 11718 11073 11746 11074
rect 11718 11047 11719 11073
rect 11719 11047 11745 11073
rect 11745 11047 11746 11073
rect 11718 11046 11746 11047
rect 11718 10793 11746 10794
rect 11718 10767 11719 10793
rect 11719 10767 11745 10793
rect 11745 10767 11746 10793
rect 11718 10766 11746 10767
rect 11662 9702 11690 9730
rect 11606 9422 11634 9450
rect 11382 9254 11410 9282
rect 12838 11913 12866 11914
rect 12838 11887 12839 11913
rect 12839 11887 12865 11913
rect 12865 11887 12866 11913
rect 12838 11886 12866 11887
rect 18830 13145 18858 13146
rect 18830 13119 18831 13145
rect 18831 13119 18857 13145
rect 18857 13119 18858 13145
rect 18830 13118 18858 13119
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 20006 12782 20034 12810
rect 13342 12614 13370 12642
rect 13174 11830 13202 11858
rect 13286 11913 13314 11914
rect 13286 11887 13287 11913
rect 13287 11887 13313 11913
rect 13313 11887 13314 11913
rect 13286 11886 13314 11887
rect 13006 11774 13034 11802
rect 14182 12334 14210 12362
rect 13734 12054 13762 12082
rect 13734 11969 13762 11970
rect 13734 11943 13735 11969
rect 13735 11943 13761 11969
rect 13761 11943 13762 11969
rect 13734 11942 13762 11943
rect 13398 11830 13426 11858
rect 13006 11185 13034 11186
rect 13006 11159 13007 11185
rect 13007 11159 13033 11185
rect 13033 11159 13034 11185
rect 13006 11158 13034 11159
rect 11830 9702 11858 9730
rect 11718 8806 11746 8834
rect 11774 8638 11802 8666
rect 11438 8470 11466 8498
rect 11326 8049 11354 8050
rect 11326 8023 11327 8049
rect 11327 8023 11353 8049
rect 11353 8023 11354 8049
rect 11326 8022 11354 8023
rect 12614 10766 12642 10794
rect 11942 9758 11970 9786
rect 12390 9758 12418 9786
rect 12166 9617 12194 9618
rect 12166 9591 12167 9617
rect 12167 9591 12193 9617
rect 12193 9591 12194 9617
rect 12166 9590 12194 9591
rect 12334 9729 12362 9730
rect 12334 9703 12335 9729
rect 12335 9703 12361 9729
rect 12361 9703 12362 9729
rect 12334 9702 12362 9703
rect 12166 8638 12194 8666
rect 12446 9673 12474 9674
rect 12446 9647 12447 9673
rect 12447 9647 12473 9673
rect 12473 9647 12474 9673
rect 12446 9646 12474 9647
rect 12726 10793 12754 10794
rect 12726 10767 12727 10793
rect 12727 10767 12753 10793
rect 12753 10767 12754 10793
rect 12726 10766 12754 10767
rect 12670 9758 12698 9786
rect 13062 11073 13090 11074
rect 13062 11047 13063 11073
rect 13063 11047 13089 11073
rect 13089 11047 13090 11073
rect 13062 11046 13090 11047
rect 13230 11046 13258 11074
rect 12950 10793 12978 10794
rect 12950 10767 12951 10793
rect 12951 10767 12977 10793
rect 12977 10767 12978 10793
rect 12950 10766 12978 10767
rect 13006 10681 13034 10682
rect 13006 10655 13007 10681
rect 13007 10655 13033 10681
rect 13033 10655 13034 10681
rect 13006 10654 13034 10655
rect 13734 10766 13762 10794
rect 13622 10737 13650 10738
rect 13622 10711 13623 10737
rect 13623 10711 13649 10737
rect 13649 10711 13650 10737
rect 13622 10710 13650 10711
rect 13454 10345 13482 10346
rect 13454 10319 13455 10345
rect 13455 10319 13481 10345
rect 13481 10319 13482 10345
rect 13454 10318 13482 10319
rect 13118 9982 13146 10010
rect 12838 9870 12866 9898
rect 12726 9702 12754 9730
rect 12446 8078 12474 8106
rect 11214 7601 11242 7602
rect 11214 7575 11215 7601
rect 11215 7575 11241 7601
rect 11241 7575 11242 7601
rect 11214 7574 11242 7575
rect 11494 7630 11522 7658
rect 11886 7574 11914 7602
rect 10934 7265 10962 7266
rect 10934 7239 10935 7265
rect 10935 7239 10961 7265
rect 10961 7239 10962 7265
rect 10934 7238 10962 7239
rect 10878 7153 10906 7154
rect 10878 7127 10879 7153
rect 10879 7127 10905 7153
rect 10905 7127 10906 7153
rect 10878 7126 10906 7127
rect 11158 7153 11186 7154
rect 11158 7127 11159 7153
rect 11159 7127 11185 7153
rect 11185 7127 11186 7153
rect 11158 7126 11186 7127
rect 10206 6958 10234 6986
rect 10766 6958 10794 6986
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 11830 6985 11858 6986
rect 11830 6959 11831 6985
rect 11831 6959 11857 6985
rect 11857 6959 11858 6985
rect 11830 6958 11858 6959
rect 11214 6734 11242 6762
rect 11606 6734 11634 6762
rect 12894 9422 12922 9450
rect 13174 9870 13202 9898
rect 13118 9254 13146 9282
rect 13286 9422 13314 9450
rect 13622 9982 13650 10010
rect 13510 9590 13538 9618
rect 13622 9870 13650 9898
rect 13174 9225 13202 9226
rect 13174 9199 13175 9225
rect 13175 9199 13201 9225
rect 13201 9199 13202 9225
rect 13174 9198 13202 9199
rect 13342 9198 13370 9226
rect 12502 7742 12530 7770
rect 12614 8526 12642 8554
rect 13118 8553 13146 8554
rect 13118 8527 13119 8553
rect 13119 8527 13145 8553
rect 13145 8527 13146 8553
rect 13118 8526 13146 8527
rect 14070 11969 14098 11970
rect 14070 11943 14071 11969
rect 14071 11943 14097 11969
rect 14097 11943 14098 11969
rect 14070 11942 14098 11943
rect 13846 11913 13874 11914
rect 13846 11887 13847 11913
rect 13847 11887 13873 11913
rect 13873 11887 13874 11913
rect 13846 11886 13874 11887
rect 18830 12361 18858 12362
rect 18830 12335 18831 12361
rect 18831 12335 18857 12361
rect 18857 12335 18858 12361
rect 18830 12334 18858 12335
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 20006 12110 20034 12138
rect 14294 11942 14322 11970
rect 18830 11969 18858 11970
rect 18830 11943 18831 11969
rect 18831 11943 18857 11969
rect 18857 11943 18858 11969
rect 18830 11942 18858 11943
rect 20006 11774 20034 11802
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 13846 10766 13874 10794
rect 14686 10766 14714 10794
rect 18830 10793 18858 10794
rect 18830 10767 18831 10793
rect 18831 10767 18857 10793
rect 18857 10767 18858 10793
rect 18830 10766 18858 10767
rect 20118 10766 20146 10794
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 20006 10430 20034 10458
rect 13902 9982 13930 10010
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 14294 9590 14322 9618
rect 18830 9617 18858 9618
rect 18830 9591 18831 9617
rect 18831 9591 18857 9617
rect 18857 9591 18858 9617
rect 18830 9590 18858 9591
rect 20006 9422 20034 9450
rect 13678 9225 13706 9226
rect 13678 9199 13679 9225
rect 13679 9199 13705 9225
rect 13705 9199 13706 9225
rect 13678 9198 13706 9199
rect 14126 9337 14154 9338
rect 14126 9311 14127 9337
rect 14127 9311 14153 9337
rect 14153 9311 14154 9337
rect 14126 9310 14154 9311
rect 14742 9310 14770 9338
rect 14070 9281 14098 9282
rect 14070 9255 14071 9281
rect 14071 9255 14097 9281
rect 14097 9255 14098 9281
rect 14070 9254 14098 9255
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 14742 8806 14770 8834
rect 13678 8497 13706 8498
rect 13678 8471 13679 8497
rect 13679 8471 13705 8497
rect 13705 8471 13706 8497
rect 13678 8470 13706 8471
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 20006 8750 20034 8778
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 12558 7630 12586 7658
rect 13342 7769 13370 7770
rect 13342 7743 13343 7769
rect 13343 7743 13369 7769
rect 13369 7743 13370 7769
rect 13342 7742 13370 7743
rect 13006 7686 13034 7714
rect 12614 7265 12642 7266
rect 12614 7239 12615 7265
rect 12615 7239 12641 7265
rect 12641 7239 12642 7265
rect 12614 7238 12642 7239
rect 12502 7153 12530 7154
rect 12502 7127 12503 7153
rect 12503 7127 12529 7153
rect 12529 7127 12530 7153
rect 12502 7126 12530 7127
rect 12334 6985 12362 6986
rect 12334 6959 12335 6985
rect 12335 6959 12361 6985
rect 12361 6959 12362 6985
rect 12334 6958 12362 6959
rect 13566 7713 13594 7714
rect 13566 7687 13567 7713
rect 13567 7687 13593 7713
rect 13593 7687 13594 7713
rect 13566 7686 13594 7687
rect 13678 7686 13706 7714
rect 13062 7630 13090 7658
rect 13118 7601 13146 7602
rect 13118 7575 13119 7601
rect 13119 7575 13145 7601
rect 13145 7575 13146 7601
rect 13118 7574 13146 7575
rect 13398 7657 13426 7658
rect 13398 7631 13399 7657
rect 13399 7631 13425 7657
rect 13425 7631 13426 7657
rect 13398 7630 13426 7631
rect 13734 7657 13762 7658
rect 13734 7631 13735 7657
rect 13735 7631 13761 7657
rect 13761 7631 13762 7657
rect 13734 7630 13762 7631
rect 14294 7630 14322 7658
rect 14070 7574 14098 7602
rect 13006 7238 13034 7266
rect 12670 6958 12698 6986
rect 13006 7126 13034 7154
rect 18830 7657 18858 7658
rect 18830 7631 18831 7657
rect 18831 7631 18857 7657
rect 18857 7631 18858 7657
rect 18830 7630 18858 7631
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 20006 7406 20034 7434
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 12278 6734 12306 6762
rect 10430 2030 10458 2058
rect 8078 1694 8106 1722
rect 9254 1721 9282 1722
rect 9254 1695 9255 1721
rect 9255 1695 9281 1721
rect 9281 1695 9282 1721
rect 9254 1694 9282 1695
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 11046 2057 11074 2058
rect 11046 2031 11047 2057
rect 11047 2031 11073 2057
rect 11073 2031 11074 2057
rect 11046 2030 11074 2031
rect 11438 1806 11466 1834
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 8409 19110 8414 19138
rect 8442 19110 9030 19138
rect 9058 19110 9063 19138
rect 12105 19110 12110 19138
rect 12138 19110 12782 19138
rect 12810 19110 12815 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 10761 18718 10766 18746
rect 10794 18718 11382 18746
rect 11410 18718 11415 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 7345 13790 7350 13818
rect 7378 13790 7910 13818
rect 7938 13790 7943 13818
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 0 13482 400 13496
rect 0 13454 2086 13482
rect 2114 13454 2119 13482
rect 0 13440 400 13454
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 2137 13230 2142 13258
rect 2170 13230 5782 13258
rect 5810 13230 5815 13258
rect 13057 13174 13062 13202
rect 13090 13174 13454 13202
rect 0 13146 400 13160
rect 13426 13146 13454 13174
rect 0 13118 966 13146
rect 994 13118 999 13146
rect 2137 13118 2142 13146
rect 2170 13118 6062 13146
rect 6090 13118 6095 13146
rect 8409 13118 8414 13146
rect 8442 13118 9366 13146
rect 9394 13118 9399 13146
rect 13426 13118 14014 13146
rect 14042 13118 18830 13146
rect 18858 13118 18863 13146
rect 0 13104 400 13118
rect 7513 13062 7518 13090
rect 7546 13062 8750 13090
rect 8778 13062 9590 13090
rect 9618 13062 10262 13090
rect 10290 13062 10934 13090
rect 10962 13062 11270 13090
rect 11298 13062 11494 13090
rect 11522 13062 12614 13090
rect 12642 13062 12647 13090
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 0 12810 400 12824
rect 20600 12810 21000 12824
rect 0 12782 966 12810
rect 994 12782 999 12810
rect 8129 12782 8134 12810
rect 8162 12782 9142 12810
rect 9170 12782 10654 12810
rect 10682 12782 10687 12810
rect 20001 12782 20006 12810
rect 20034 12782 21000 12810
rect 0 12768 400 12782
rect 20600 12768 21000 12782
rect 7345 12726 7350 12754
rect 7378 12726 7518 12754
rect 7546 12726 8414 12754
rect 8442 12726 8447 12754
rect 5777 12670 5782 12698
rect 5810 12670 7294 12698
rect 7322 12670 7327 12698
rect 7793 12670 7798 12698
rect 7826 12670 8190 12698
rect 8218 12670 9646 12698
rect 9674 12670 9679 12698
rect 10705 12670 10710 12698
rect 10738 12670 11046 12698
rect 11074 12670 11079 12698
rect 6057 12614 6062 12642
rect 6090 12614 7574 12642
rect 7602 12614 7607 12642
rect 9193 12614 9198 12642
rect 9226 12614 9758 12642
rect 9786 12614 9791 12642
rect 12665 12614 12670 12642
rect 12698 12614 13342 12642
rect 13370 12614 13375 12642
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 7849 12334 7854 12362
rect 7882 12334 10150 12362
rect 10178 12334 10183 12362
rect 14177 12334 14182 12362
rect 14210 12334 18830 12362
rect 18858 12334 18863 12362
rect 7121 12278 7126 12306
rect 7154 12278 7910 12306
rect 7938 12278 7943 12306
rect 10369 12278 10374 12306
rect 10402 12278 11102 12306
rect 11130 12278 12978 12306
rect 12950 12250 12978 12278
rect 12945 12222 12950 12250
rect 12978 12222 12983 12250
rect 12721 12166 12726 12194
rect 12754 12166 13062 12194
rect 13090 12166 13095 12194
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 20600 12138 21000 12152
rect 20001 12110 20006 12138
rect 20034 12110 21000 12138
rect 20600 12096 21000 12110
rect 8185 12054 8190 12082
rect 8218 12054 11214 12082
rect 11242 12054 13734 12082
rect 13762 12054 13767 12082
rect 10369 11998 10374 12026
rect 10402 11998 10878 12026
rect 10906 11998 10911 12026
rect 9585 11942 9590 11970
rect 9618 11942 11550 11970
rect 11578 11942 11830 11970
rect 11858 11942 11863 11970
rect 13729 11942 13734 11970
rect 13762 11942 14070 11970
rect 14098 11942 14294 11970
rect 14322 11942 18830 11970
rect 18858 11942 18863 11970
rect 8353 11886 8358 11914
rect 8386 11886 9898 11914
rect 9977 11886 9982 11914
rect 10010 11886 10374 11914
rect 10402 11886 10407 11914
rect 11265 11886 11270 11914
rect 11298 11886 12838 11914
rect 12866 11886 13286 11914
rect 13314 11886 13319 11914
rect 13841 11886 13846 11914
rect 13874 11886 13879 11914
rect 9870 11858 9898 11886
rect 9870 11830 10206 11858
rect 10234 11830 10239 11858
rect 10761 11830 10766 11858
rect 10794 11830 11438 11858
rect 11466 11830 13174 11858
rect 13202 11830 13398 11858
rect 13426 11830 13431 11858
rect 13846 11802 13874 11886
rect 20600 11802 21000 11816
rect 9193 11774 9198 11802
rect 9226 11774 9366 11802
rect 9394 11774 9814 11802
rect 9842 11774 9847 11802
rect 13001 11774 13006 11802
rect 13034 11774 13874 11802
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 20600 11760 21000 11774
rect 6785 11662 6790 11690
rect 6818 11662 7630 11690
rect 7658 11662 8330 11690
rect 7177 11550 7182 11578
rect 7210 11550 7742 11578
rect 7770 11550 7775 11578
rect 8302 11522 8330 11662
rect 9081 11606 9086 11634
rect 9114 11606 9422 11634
rect 9450 11606 9455 11634
rect 8297 11494 8302 11522
rect 8330 11494 10094 11522
rect 10122 11494 10127 11522
rect 6673 11438 6678 11466
rect 6706 11438 7126 11466
rect 7154 11438 7159 11466
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 8857 11270 8862 11298
rect 8890 11270 9310 11298
rect 9338 11270 9343 11298
rect 961 11214 966 11242
rect 994 11214 999 11242
rect 7681 11214 7686 11242
rect 7714 11214 8414 11242
rect 8442 11214 8447 11242
rect 8801 11214 8806 11242
rect 8834 11214 8839 11242
rect 0 11130 400 11144
rect 966 11130 994 11214
rect 2137 11158 2142 11186
rect 2170 11158 5614 11186
rect 5642 11158 7574 11186
rect 7602 11158 7607 11186
rect 7686 11130 7714 11214
rect 8806 11186 8834 11214
rect 8633 11158 8638 11186
rect 8666 11158 9114 11186
rect 9417 11158 9422 11186
rect 9450 11158 9702 11186
rect 9730 11158 9735 11186
rect 9809 11158 9814 11186
rect 9842 11158 9982 11186
rect 10010 11158 11662 11186
rect 11690 11158 13006 11186
rect 13034 11158 13039 11186
rect 9086 11130 9114 11158
rect 0 11102 994 11130
rect 7345 11102 7350 11130
rect 7378 11102 7714 11130
rect 8185 11102 8190 11130
rect 8218 11102 8806 11130
rect 8834 11102 8839 11130
rect 9081 11102 9086 11130
rect 9114 11102 9926 11130
rect 9954 11102 10430 11130
rect 10458 11102 10463 11130
rect 0 11088 400 11102
rect 7737 11046 7742 11074
rect 7770 11046 8022 11074
rect 8050 11046 8055 11074
rect 8451 11046 8470 11074
rect 8498 11046 8503 11074
rect 10593 11046 10598 11074
rect 10626 11046 11046 11074
rect 11074 11046 11550 11074
rect 11578 11046 11583 11074
rect 11713 11046 11718 11074
rect 11746 11046 13062 11074
rect 13090 11046 13230 11074
rect 13258 11046 13263 11074
rect 10649 10990 10654 11018
rect 10682 10990 10878 11018
rect 10906 10990 10911 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 7737 10934 7742 10962
rect 7770 10934 8022 10962
rect 8050 10934 8694 10962
rect 8722 10934 8727 10962
rect 10145 10934 10150 10962
rect 10178 10934 10262 10962
rect 10290 10934 10822 10962
rect 10850 10934 11214 10962
rect 11242 10934 11247 10962
rect 7121 10878 7126 10906
rect 7154 10878 8078 10906
rect 8106 10878 8111 10906
rect 9921 10878 9926 10906
rect 9954 10878 10374 10906
rect 10402 10878 10878 10906
rect 10906 10878 10911 10906
rect 7065 10822 7070 10850
rect 7098 10822 7518 10850
rect 7546 10822 7910 10850
rect 7938 10822 8750 10850
rect 8778 10822 8783 10850
rect 10145 10822 10150 10850
rect 10178 10822 10822 10850
rect 10850 10822 11158 10850
rect 11186 10822 11191 10850
rect 20600 10794 21000 10808
rect 2137 10766 2142 10794
rect 2170 10766 4998 10794
rect 5026 10766 5031 10794
rect 9865 10766 9870 10794
rect 9898 10766 10206 10794
rect 10234 10766 10542 10794
rect 10570 10766 10575 10794
rect 11713 10766 11718 10794
rect 11746 10766 12614 10794
rect 12642 10766 12726 10794
rect 12754 10766 12759 10794
rect 12945 10766 12950 10794
rect 12978 10766 13734 10794
rect 13762 10766 13767 10794
rect 13841 10766 13846 10794
rect 13874 10766 14686 10794
rect 14714 10766 18830 10794
rect 18858 10766 18863 10794
rect 20113 10766 20118 10794
rect 20146 10766 21000 10794
rect 20600 10752 21000 10766
rect 6057 10710 6062 10738
rect 6090 10710 7294 10738
rect 7322 10710 7327 10738
rect 7401 10710 7406 10738
rect 7434 10710 7854 10738
rect 7882 10710 7887 10738
rect 9585 10710 9590 10738
rect 9618 10710 10598 10738
rect 10626 10710 10631 10738
rect 13426 10710 13622 10738
rect 13650 10710 13655 10738
rect 13426 10682 13454 10710
rect 13001 10654 13006 10682
rect 13034 10654 13454 10682
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 2081 10486 2086 10514
rect 2114 10486 9702 10514
rect 9730 10486 10934 10514
rect 10962 10486 10967 10514
rect 0 10458 400 10472
rect 20600 10458 21000 10472
rect 0 10430 966 10458
rect 994 10430 999 10458
rect 4993 10430 4998 10458
rect 5026 10430 6958 10458
rect 6986 10430 6991 10458
rect 7961 10430 7966 10458
rect 7994 10430 9870 10458
rect 9898 10430 9903 10458
rect 20001 10430 20006 10458
rect 20034 10430 21000 10458
rect 0 10416 400 10430
rect 20600 10416 21000 10430
rect 6449 10374 6454 10402
rect 6482 10374 6790 10402
rect 6818 10374 7238 10402
rect 7266 10374 7271 10402
rect 9809 10374 9814 10402
rect 9842 10374 10150 10402
rect 10178 10374 10183 10402
rect 9249 10318 9254 10346
rect 9282 10318 13454 10346
rect 13482 10318 13487 10346
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 8409 10094 8414 10122
rect 8442 10094 8918 10122
rect 8946 10094 8951 10122
rect 7569 10038 7574 10066
rect 7602 10038 8078 10066
rect 8106 10038 8111 10066
rect 8129 9982 8134 10010
rect 8162 9982 8918 10010
rect 8946 9982 8951 10010
rect 10033 9982 10038 10010
rect 10066 9982 10878 10010
rect 10906 9982 10911 10010
rect 13113 9982 13118 10010
rect 13146 9982 13622 10010
rect 13650 9982 13902 10010
rect 13930 9982 13935 10010
rect 7569 9926 7574 9954
rect 7602 9926 7742 9954
rect 7770 9926 7775 9954
rect 7849 9926 7854 9954
rect 7882 9926 9254 9954
rect 9282 9926 9287 9954
rect 9417 9926 9422 9954
rect 9450 9926 10654 9954
rect 10682 9926 10687 9954
rect 9254 9898 9282 9926
rect 9254 9870 10206 9898
rect 10234 9870 10239 9898
rect 10929 9870 10934 9898
rect 10962 9870 12838 9898
rect 12866 9870 13174 9898
rect 13202 9870 13622 9898
rect 13650 9870 13655 9898
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 7686 9758 10766 9786
rect 10794 9758 10799 9786
rect 11937 9758 11942 9786
rect 11970 9758 12390 9786
rect 12418 9758 12670 9786
rect 12698 9758 12703 9786
rect 7686 9674 7714 9758
rect 8969 9702 8974 9730
rect 9002 9702 9814 9730
rect 9842 9702 11662 9730
rect 11690 9702 11830 9730
rect 11858 9702 11863 9730
rect 12329 9702 12334 9730
rect 12362 9702 12726 9730
rect 12754 9702 12759 9730
rect 7233 9646 7238 9674
rect 7266 9646 7686 9674
rect 7714 9646 7719 9674
rect 9305 9646 9310 9674
rect 9338 9646 9926 9674
rect 9954 9646 9959 9674
rect 10089 9646 10094 9674
rect 10122 9646 10430 9674
rect 10458 9646 10463 9674
rect 10705 9646 10710 9674
rect 10738 9646 11102 9674
rect 11130 9646 12446 9674
rect 12474 9646 12479 9674
rect 9641 9590 9646 9618
rect 9674 9590 9982 9618
rect 10010 9590 10015 9618
rect 10313 9590 10318 9618
rect 10346 9590 12166 9618
rect 12194 9590 12199 9618
rect 13505 9590 13510 9618
rect 13538 9590 14294 9618
rect 14322 9590 18830 9618
rect 18858 9590 18863 9618
rect 9361 9534 9366 9562
rect 9394 9534 9702 9562
rect 9730 9534 9735 9562
rect 9814 9534 10878 9562
rect 10906 9534 11214 9562
rect 11242 9534 11247 9562
rect 9366 9506 9394 9534
rect 6673 9478 6678 9506
rect 6706 9478 7294 9506
rect 7322 9478 7327 9506
rect 8409 9478 8414 9506
rect 8442 9478 9394 9506
rect 0 9450 400 9464
rect 9814 9450 9842 9534
rect 10089 9478 10094 9506
rect 10122 9478 10710 9506
rect 10738 9478 10743 9506
rect 20600 9450 21000 9464
rect 0 9422 966 9450
rect 994 9422 999 9450
rect 8073 9422 8078 9450
rect 8106 9422 9842 9450
rect 11601 9422 11606 9450
rect 11634 9422 12894 9450
rect 12922 9422 13286 9450
rect 13314 9422 13319 9450
rect 20001 9422 20006 9450
rect 20034 9422 21000 9450
rect 0 9408 400 9422
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 20600 9408 21000 9422
rect 7625 9366 7630 9394
rect 7658 9366 7910 9394
rect 7938 9366 7943 9394
rect 7569 9310 7574 9338
rect 7602 9310 8918 9338
rect 8946 9310 8951 9338
rect 9137 9310 9142 9338
rect 9170 9310 9646 9338
rect 9674 9310 9679 9338
rect 14121 9310 14126 9338
rect 14154 9310 14742 9338
rect 14770 9310 14775 9338
rect 7681 9254 7686 9282
rect 7714 9254 7719 9282
rect 9305 9254 9310 9282
rect 9338 9254 9343 9282
rect 9753 9254 9758 9282
rect 9786 9254 10318 9282
rect 10346 9254 10351 9282
rect 10481 9254 10486 9282
rect 10514 9254 11382 9282
rect 11410 9254 11415 9282
rect 13113 9254 13118 9282
rect 13146 9254 14070 9282
rect 14098 9254 14103 9282
rect 7686 9170 7714 9254
rect 9310 9226 9338 9254
rect 13342 9226 13370 9254
rect 8409 9198 8414 9226
rect 8442 9198 8862 9226
rect 8890 9198 8895 9226
rect 9025 9198 9030 9226
rect 9058 9198 9338 9226
rect 9478 9198 9702 9226
rect 9730 9198 9735 9226
rect 10425 9198 10430 9226
rect 10458 9198 11046 9226
rect 11074 9198 13174 9226
rect 13202 9198 13207 9226
rect 13337 9198 13342 9226
rect 13370 9198 13375 9226
rect 13659 9198 13678 9226
rect 13706 9198 13711 9226
rect 9478 9170 9506 9198
rect 2137 9142 2142 9170
rect 2170 9142 5614 9170
rect 5642 9142 5647 9170
rect 7233 9142 7238 9170
rect 7266 9142 8050 9170
rect 8241 9142 8246 9170
rect 8274 9142 9254 9170
rect 9282 9142 9506 9170
rect 9585 9142 9590 9170
rect 9618 9142 11102 9170
rect 11130 9142 11135 9170
rect 8022 9114 8050 9142
rect 8017 9086 8022 9114
rect 8050 9086 9534 9114
rect 9562 9086 10038 9114
rect 10066 9086 10071 9114
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 7961 8974 7966 9002
rect 7994 8974 10038 9002
rect 10066 8974 10071 9002
rect 7065 8862 7070 8890
rect 7098 8862 7350 8890
rect 7378 8862 7383 8890
rect 7793 8862 7798 8890
rect 7826 8862 8246 8890
rect 8274 8862 8279 8890
rect 8857 8806 8862 8834
rect 8890 8806 9366 8834
rect 9394 8806 9399 8834
rect 10257 8806 10262 8834
rect 10290 8806 11718 8834
rect 11746 8806 11751 8834
rect 14737 8806 14742 8834
rect 14770 8806 18830 8834
rect 18858 8806 18863 8834
rect 20600 8778 21000 8792
rect 5609 8750 5614 8778
rect 5642 8750 7182 8778
rect 7210 8750 7215 8778
rect 7737 8750 7742 8778
rect 7770 8750 8246 8778
rect 8274 8750 8470 8778
rect 8498 8750 8503 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 20600 8736 21000 8750
rect 9305 8694 9310 8722
rect 9338 8694 9702 8722
rect 9730 8694 10318 8722
rect 10346 8694 10351 8722
rect 10145 8638 10150 8666
rect 10178 8638 10654 8666
rect 10682 8638 11774 8666
rect 11802 8638 12166 8666
rect 12194 8638 12199 8666
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 7233 8526 7238 8554
rect 7266 8526 10710 8554
rect 10738 8526 10743 8554
rect 12609 8526 12614 8554
rect 12642 8526 13118 8554
rect 13146 8526 13151 8554
rect 7546 8470 7630 8498
rect 7658 8470 7663 8498
rect 10929 8470 10934 8498
rect 10962 8470 11438 8498
rect 11466 8470 11471 8498
rect 13659 8470 13678 8498
rect 13706 8470 13711 8498
rect 7546 8442 7574 8470
rect 2137 8414 2142 8442
rect 2170 8414 5950 8442
rect 5978 8414 7574 8442
rect 7121 8358 7126 8386
rect 7154 8358 7574 8386
rect 7602 8358 7607 8386
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 0 8106 400 8120
rect 0 8078 966 8106
rect 994 8078 999 8106
rect 8017 8078 8022 8106
rect 8050 8078 9142 8106
rect 9170 8078 12446 8106
rect 12474 8078 12479 8106
rect 0 8064 400 8078
rect 10369 8022 10374 8050
rect 10402 8022 10822 8050
rect 10850 8022 11326 8050
rect 11354 8022 11359 8050
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 8465 7742 8470 7770
rect 8498 7742 8806 7770
rect 8834 7742 8839 7770
rect 12497 7742 12502 7770
rect 12530 7742 13342 7770
rect 13370 7742 13375 7770
rect 7625 7686 7630 7714
rect 7658 7686 8078 7714
rect 8106 7686 8111 7714
rect 10257 7686 10262 7714
rect 10290 7686 10710 7714
rect 10738 7686 10743 7714
rect 13001 7686 13006 7714
rect 13034 7686 13566 7714
rect 13594 7686 13599 7714
rect 13673 7686 13678 7714
rect 13706 7686 14322 7714
rect 14294 7658 14322 7686
rect 9473 7630 9478 7658
rect 9506 7630 9758 7658
rect 9786 7630 10094 7658
rect 10122 7630 10127 7658
rect 11489 7630 11494 7658
rect 11522 7630 11527 7658
rect 12553 7630 12558 7658
rect 12586 7630 13062 7658
rect 13090 7630 13095 7658
rect 13393 7630 13398 7658
rect 13426 7630 13734 7658
rect 13762 7630 13767 7658
rect 14289 7630 14294 7658
rect 14322 7630 18830 7658
rect 18858 7630 18863 7658
rect 11494 7602 11522 7630
rect 7457 7574 7462 7602
rect 7490 7574 7854 7602
rect 7882 7574 7887 7602
rect 11209 7574 11214 7602
rect 11242 7574 11886 7602
rect 11914 7574 11919 7602
rect 13113 7574 13118 7602
rect 13146 7574 14070 7602
rect 14098 7574 14103 7602
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 20600 7434 21000 7448
rect 20001 7406 20006 7434
rect 20034 7406 21000 7434
rect 20600 7392 21000 7406
rect 10257 7238 10262 7266
rect 10290 7238 10934 7266
rect 10962 7238 12614 7266
rect 12642 7238 13006 7266
rect 13034 7238 13039 7266
rect 6673 7126 6678 7154
rect 6706 7126 7518 7154
rect 7546 7126 8470 7154
rect 8498 7126 8503 7154
rect 9417 7126 9422 7154
rect 9450 7126 10094 7154
rect 10122 7126 10127 7154
rect 10873 7126 10878 7154
rect 10906 7126 11158 7154
rect 11186 7126 11191 7154
rect 12497 7126 12502 7154
rect 12530 7126 13006 7154
rect 13034 7126 13039 7154
rect 9025 7070 9030 7098
rect 9058 7070 9366 7098
rect 9394 7070 9399 7098
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 8409 6958 8414 6986
rect 8442 6958 8862 6986
rect 8890 6958 9198 6986
rect 9226 6958 9231 6986
rect 10201 6958 10206 6986
rect 10234 6958 10766 6986
rect 10794 6958 11830 6986
rect 11858 6958 12334 6986
rect 12362 6958 12670 6986
rect 12698 6958 12703 6986
rect 11209 6734 11214 6762
rect 11242 6734 11606 6762
rect 11634 6734 12278 6762
rect 12306 6734 12311 6762
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 10425 2030 10430 2058
rect 10458 2030 11046 2058
rect 11074 2030 11079 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 11433 1806 11438 1834
rect 11466 1806 12782 1834
rect 12810 1806 12815 1834
rect 8073 1694 8078 1722
rect 8106 1694 9254 1722
rect 9282 1694 9287 1722
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 8470 11046 8498 11074
rect 10878 10990 10906 11018
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 10878 9534 10906 9562
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 13678 9198 13706 9226
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 8470 8750 8498 8778
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 13678 8470 13706 8498
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 8470 7742 8498 7770
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 8470 11074 8498 11079
rect 8470 8778 8498 11046
rect 8470 7770 8498 8750
rect 8470 7737 8498 7742
rect 9904 10990 10064 11746
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 10878 11018 10906 11023
rect 10878 9562 10906 10990
rect 10878 9529 10906 9534
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 13678 9226 13706 9231
rect 13678 8498 13706 9198
rect 13678 8465 13706 8470
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9856 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8176 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8680 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9128 0 1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_
timestamp 1698175906
transform -1 0 10472 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_
timestamp 1698175906
transform 1 0 11144 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1698175906
transform -1 0 10808 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10136 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _112_
timestamp 1698175906
transform -1 0 11368 0 1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8176 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform -1 0 9576 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7448 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8064 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _118_
timestamp 1698175906
transform -1 0 7448 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _119_
timestamp 1698175906
transform 1 0 9072 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8736 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _121_
timestamp 1698175906
transform -1 0 10192 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8736 0 -1 11760
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _123_
timestamp 1698175906
transform -1 0 7168 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8568 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform -1 0 8232 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _126_
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _127_
timestamp 1698175906
transform -1 0 10024 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698175906
transform -1 0 8512 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _129_
timestamp 1698175906
transform -1 0 10472 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _130_
timestamp 1698175906
transform -1 0 9464 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _131_
timestamp 1698175906
transform 1 0 8288 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _132_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7504 0 -1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _133_
timestamp 1698175906
transform -1 0 7616 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _134_
timestamp 1698175906
transform -1 0 7392 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _135_
timestamp 1698175906
transform 1 0 11088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _136_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11984 0 1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _137_
timestamp 1698175906
transform -1 0 12264 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _138_
timestamp 1698175906
transform -1 0 9184 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _139_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8568 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _140_
timestamp 1698175906
transform -1 0 9968 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _141_
timestamp 1698175906
transform -1 0 9296 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _142_
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _143_
timestamp 1698175906
transform -1 0 8960 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _144_
timestamp 1698175906
transform -1 0 8232 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _145_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9968 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _146_
timestamp 1698175906
transform 1 0 13384 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _147_
timestamp 1698175906
transform -1 0 13384 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_
timestamp 1698175906
transform 1 0 13496 0 -1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _149_
timestamp 1698175906
transform -1 0 13496 0 -1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _150_
timestamp 1698175906
transform -1 0 9968 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _151_
timestamp 1698175906
transform -1 0 11144 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _152_
timestamp 1698175906
transform 1 0 8008 0 -1 13328
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _153_
timestamp 1698175906
transform -1 0 8064 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _154_
timestamp 1698175906
transform -1 0 10360 0 1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _155_
timestamp 1698175906
transform -1 0 9520 0 -1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _156_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11760 0 1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _157_
timestamp 1698175906
transform 1 0 11480 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _158_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _159_
timestamp 1698175906
transform 1 0 13104 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _160_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9128 0 -1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _161_
timestamp 1698175906
transform 1 0 9912 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _162_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13552 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _163_
timestamp 1698175906
transform 1 0 14000 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _164_
timestamp 1698175906
transform 1 0 13552 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _165_
timestamp 1698175906
transform 1 0 11144 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _166_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _167_
timestamp 1698175906
transform -1 0 14000 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _168_
timestamp 1698175906
transform 1 0 9520 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _169_
timestamp 1698175906
transform 1 0 12936 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _170_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13160 0 -1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _171_
timestamp 1698175906
transform -1 0 11312 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _172_
timestamp 1698175906
transform 1 0 9296 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _173_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10920 0 -1 9408
box -43 -43 1107 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _174_
timestamp 1698175906
transform 1 0 9968 0 1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _175_
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _176_
timestamp 1698175906
transform -1 0 7840 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform -1 0 8176 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _178_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7896 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _179_
timestamp 1698175906
transform 1 0 7056 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _180_
timestamp 1698175906
transform 1 0 6888 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _181_
timestamp 1698175906
transform -1 0 8344 0 -1 10192
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _182_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7784 0 -1 10976
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _183_
timestamp 1698175906
transform 1 0 9016 0 -1 13328
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _184_
timestamp 1698175906
transform -1 0 9408 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _185_
timestamp 1698175906
transform 1 0 10136 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _186_
timestamp 1698175906
transform -1 0 9744 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _187_
timestamp 1698175906
transform -1 0 12040 0 -1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _188_
timestamp 1698175906
transform 1 0 11088 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _189_
timestamp 1698175906
transform 1 0 8848 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _190_
timestamp 1698175906
transform -1 0 7728 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _191_
timestamp 1698175906
transform 1 0 7784 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _192_
timestamp 1698175906
transform 1 0 9576 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _193_
timestamp 1698175906
transform -1 0 11704 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _194_
timestamp 1698175906
transform -1 0 10864 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _195_
timestamp 1698175906
transform 1 0 9912 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _196_
timestamp 1698175906
transform -1 0 7336 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _197_
timestamp 1698175906
transform 1 0 7056 0 1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _198_
timestamp 1698175906
transform -1 0 13216 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _199_
timestamp 1698175906
transform 1 0 11704 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _200_
timestamp 1698175906
transform 1 0 12656 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _201_
timestamp 1698175906
transform -1 0 12936 0 1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _202_
timestamp 1698175906
transform 1 0 12544 0 1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _203_
timestamp 1698175906
transform 1 0 13496 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _204_
timestamp 1698175906
transform 1 0 13048 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _205_
timestamp 1698175906
transform -1 0 13216 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _206_
timestamp 1698175906
transform -1 0 12600 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _207_
timestamp 1698175906
transform 1 0 12264 0 1 7056
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7616 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform -1 0 7336 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform -1 0 7168 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 10808 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform -1 0 12656 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform -1 0 9352 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 12768 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 6888 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 8792 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 12768 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 13216 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 9688 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 13160 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 10080 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform -1 0 7504 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform -1 0 6552 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 8512 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 10864 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform -1 0 8232 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 9520 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform -1 0 7168 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 12488 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 12768 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _236_
timestamp 1698175906
transform -1 0 11144 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _237_
timestamp 1698175906
transform 1 0 13944 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__117__A2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8176 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__164__A1
timestamp 1698175906
transform -1 0 13552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__A2
timestamp 1698175906
transform -1 0 8008 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__A2
timestamp 1698175906
transform 1 0 10864 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__B1
timestamp 1698175906
transform 1 0 7672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__A2
timestamp 1698175906
transform 1 0 13328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__A2
timestamp 1698175906
transform 1 0 13384 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 7616 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 7448 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 7224 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 10024 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 10920 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 9464 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 8288 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 8736 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform -1 0 10808 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 13104 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 11424 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 11816 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 7616 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 6776 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 10248 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 11256 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 8344 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 11480 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 7448 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 12320 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 9912 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 12432 0 -1 8624
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform -1 0 12264 0 -1 11760
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_104 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_112 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6944 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_114 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7056 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_119 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7336 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_135
timestamp 1698175906
transform 1 0 8232 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_164 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9856 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_168
timestamp 1698175906
transform 1 0 10080 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_245
timestamp 1698175906
transform 1 0 14392 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_261
timestamp 1698175906
transform 1 0 15288 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_269
timestamp 1698175906
transform 1 0 15736 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_271
timestamp 1698175906
transform 1 0 15848 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_174
timestamp 1698175906
transform 1 0 10416 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_201
timestamp 1698175906
transform 1 0 11928 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_220
timestamp 1698175906
transform 1 0 12992 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_222
timestamp 1698175906
transform 1 0 13104 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_249
timestamp 1698175906
transform 1 0 14616 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_265
timestamp 1698175906
transform 1 0 15512 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_273
timestamp 1698175906
transform 1 0 15960 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_277
timestamp 1698175906
transform 1 0 16184 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698175906
transform 1 0 16296 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_139
timestamp 1698175906
transform 1 0 8456 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_143
timestamp 1698175906
transform 1 0 8680 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 10416 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_181
timestamp 1698175906
transform 1 0 10808 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_104
timestamp 1698175906
transform 1 0 6496 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_135
timestamp 1698175906
transform 1 0 8232 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698175906
transform 1 0 8456 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_150
timestamp 1698175906
transform 1 0 9072 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_152
timestamp 1698175906
transform 1 0 9184 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_158
timestamp 1698175906
transform 1 0 9520 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_166
timestamp 1698175906
transform 1 0 9968 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_197
timestamp 1698175906
transform 1 0 11704 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_201
timestamp 1698175906
transform 1 0 11928 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_205
timestamp 1698175906
transform 1 0 12152 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_207
timestamp 1698175906
transform 1 0 12264 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_241
timestamp 1698175906
transform 1 0 14168 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_273
timestamp 1698175906
transform 1 0 15960 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_277
timestamp 1698175906
transform 1 0 16184 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698175906
transform 1 0 16296 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_115
timestamp 1698175906
transform 1 0 7112 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_119
timestamp 1698175906
transform 1 0 7336 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_155
timestamp 1698175906
transform 1 0 9352 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_159
timestamp 1698175906
transform 1 0 9576 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_167
timestamp 1698175906
transform 1 0 10024 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698175906
transform 1 0 10360 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_190
timestamp 1698175906
transform 1 0 11312 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_206
timestamp 1698175906
transform 1 0 12208 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_88
timestamp 1698175906
transform 1 0 5600 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_92
timestamp 1698175906
transform 1 0 5824 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_122
timestamp 1698175906
transform 1 0 7504 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_126
timestamp 1698175906
transform 1 0 7728 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_133
timestamp 1698175906
transform 1 0 8120 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698175906
transform 1 0 8344 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698175906
transform 1 0 8456 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_150
timestamp 1698175906
transform 1 0 9072 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_158
timestamp 1698175906
transform 1 0 9520 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_160
timestamp 1698175906
transform 1 0 9632 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_190
timestamp 1698175906
transform 1 0 11312 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_194
timestamp 1698175906
transform 1 0 11536 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_216
timestamp 1698175906
transform 1 0 12768 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_234
timestamp 1698175906
transform 1 0 13776 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_266
timestamp 1698175906
transform 1 0 15568 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_274
timestamp 1698175906
transform 1 0 16016 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698175906
transform 1 0 16240 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_314
timestamp 1698175906
transform 1 0 18256 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_322
timestamp 1698175906
transform 1 0 18704 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_139
timestamp 1698175906
transform 1 0 8456 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_147
timestamp 1698175906
transform 1 0 8904 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_154
timestamp 1698175906
transform 1 0 9296 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_170
timestamp 1698175906
transform 1 0 10192 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 10416 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_195
timestamp 1698175906
transform 1 0 11592 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_203
timestamp 1698175906
transform 1 0 12040 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_213
timestamp 1698175906
transform 1 0 12600 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_227
timestamp 1698175906
transform 1 0 13384 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 14280 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 2240 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 4032 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 4480 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_104
timestamp 1698175906
transform 1 0 6496 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_112
timestamp 1698175906
transform 1 0 6944 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_128
timestamp 1698175906
transform 1 0 7840 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698175906
transform 1 0 8288 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_158
timestamp 1698175906
transform 1 0 9520 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_220
timestamp 1698175906
transform 1 0 12992 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_253
timestamp 1698175906
transform 1 0 14840 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_269
timestamp 1698175906
transform 1 0 15736 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698175906
transform 1 0 16184 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 16296 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 20048 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 20160 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_111
timestamp 1698175906
transform 1 0 6888 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_113
timestamp 1698175906
transform 1 0 7000 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_119
timestamp 1698175906
transform 1 0 7336 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_123
timestamp 1698175906
transform 1 0 7560 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_127
timestamp 1698175906
transform 1 0 7784 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_131
timestamp 1698175906
transform 1 0 8008 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_133
timestamp 1698175906
transform 1 0 8120 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_140
timestamp 1698175906
transform 1 0 8512 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_144
timestamp 1698175906
transform 1 0 8736 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_177
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_181
timestamp 1698175906
transform 1 0 10808 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_214
timestamp 1698175906
transform 1 0 12656 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_222
timestamp 1698175906
transform 1 0 13104 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_226
timestamp 1698175906
transform 1 0 13328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_230
timestamp 1698175906
transform 1 0 13552 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_238
timestamp 1698175906
transform 1 0 14000 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_242
timestamp 1698175906
transform 1 0 14224 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 14336 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_80
timestamp 1698175906
transform 1 0 5152 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_84
timestamp 1698175906
transform 1 0 5376 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_86
timestamp 1698175906
transform 1 0 5488 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_116
timestamp 1698175906
transform 1 0 7168 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_118
timestamp 1698175906
transform 1 0 7280 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_183
timestamp 1698175906
transform 1 0 10920 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_191
timestamp 1698175906
transform 1 0 11368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_195
timestamp 1698175906
transform 1 0 11592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_202
timestamp 1698175906
transform 1 0 11984 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698175906
transform 1 0 12264 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 12376 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_216
timestamp 1698175906
transform 1 0 12768 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_220
timestamp 1698175906
transform 1 0 12992 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_243
timestamp 1698175906
transform 1 0 14280 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_275
timestamp 1698175906
transform 1 0 16072 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 16296 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 20048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 20160 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698175906
transform 1 0 2240 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698175906
transform 1 0 2464 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_111
timestamp 1698175906
transform 1 0 6888 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_113
timestamp 1698175906
transform 1 0 7000 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_123
timestamp 1698175906
transform 1 0 7560 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_127
timestamp 1698175906
transform 1 0 7784 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_164
timestamp 1698175906
transform 1 0 9856 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698175906
transform 1 0 10360 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_185
timestamp 1698175906
transform 1 0 11032 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_190
timestamp 1698175906
transform 1 0 11312 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_198
timestamp 1698175906
transform 1 0 11760 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_215
timestamp 1698175906
transform 1 0 12712 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_104
timestamp 1698175906
transform 1 0 6496 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_120
timestamp 1698175906
transform 1 0 7392 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_137
timestamp 1698175906
transform 1 0 8344 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 8456 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_158
timestamp 1698175906
transform 1 0 9520 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_162
timestamp 1698175906
transform 1 0 9744 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_165
timestamp 1698175906
transform 1 0 9912 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_230
timestamp 1698175906
transform 1 0 13552 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_262
timestamp 1698175906
transform 1 0 15344 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 16240 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 20048 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 20160 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 4536 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 4760 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 4872 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_115
timestamp 1698175906
transform 1 0 7112 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_124
timestamp 1698175906
transform 1 0 7616 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_132
timestamp 1698175906
transform 1 0 8064 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_140
timestamp 1698175906
transform 1 0 8512 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_156
timestamp 1698175906
transform 1 0 9408 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_160
timestamp 1698175906
transform 1 0 9632 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_238
timestamp 1698175906
transform 1 0 14000 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1698175906
transform 1 0 14224 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 14336 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 2240 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 4032 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 4480 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_80
timestamp 1698175906
transform 1 0 5152 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_84
timestamp 1698175906
transform 1 0 5376 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_86
timestamp 1698175906
transform 1 0 5488 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_135
timestamp 1698175906
transform 1 0 8232 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698175906
transform 1 0 8456 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_142
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_152
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_156
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_198
timestamp 1698175906
transform 1 0 11760 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698175906
transform 1 0 12208 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_252
timestamp 1698175906
transform 1 0 14784 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_268
timestamp 1698175906
transform 1 0 15680 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698175906
transform 1 0 16128 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 2240 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 2464 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_148
timestamp 1698175906
transform 1 0 8960 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_157
timestamp 1698175906
transform 1 0 9464 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_168
timestamp 1698175906
transform 1 0 10080 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_199
timestamp 1698175906
transform 1 0 11816 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_207
timestamp 1698175906
transform 1 0 12264 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_211
timestamp 1698175906
transform 1 0 12488 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_224
timestamp 1698175906
transform 1 0 13216 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_228
timestamp 1698175906
transform 1 0 13440 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 14336 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_333
timestamp 1698175906
transform 1 0 19320 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_341
timestamp 1698175906
transform 1 0 19768 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_104
timestamp 1698175906
transform 1 0 6496 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_112
timestamp 1698175906
transform 1 0 6944 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_120
timestamp 1698175906
transform 1 0 7392 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_131
timestamp 1698175906
transform 1 0 8008 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_135
timestamp 1698175906
transform 1 0 8232 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698175906
transform 1 0 8400 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698175906
transform 1 0 12264 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_220
timestamp 1698175906
transform 1 0 12992 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_224
timestamp 1698175906
transform 1 0 13216 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_226
timestamp 1698175906
transform 1 0 13328 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_229
timestamp 1698175906
transform 1 0 13496 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_261
timestamp 1698175906
transform 1 0 15288 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 16184 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 16296 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 20048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 20160 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_123
timestamp 1698175906
transform 1 0 7560 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_126
timestamp 1698175906
transform 1 0 7728 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_148
timestamp 1698175906
transform 1 0 8960 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_181
timestamp 1698175906
transform 1 0 10808 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_197
timestamp 1698175906
transform 1 0 11704 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_205
timestamp 1698175906
transform 1 0 12152 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_209
timestamp 1698175906
transform 1 0 12376 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_211
timestamp 1698175906
transform 1 0 12488 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 14280 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_88
timestamp 1698175906
transform 1 0 5600 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_92
timestamp 1698175906
transform 1 0 5824 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_94
timestamp 1698175906
transform 1 0 5936 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_132
timestamp 1698175906
transform 1 0 8064 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698175906
transform 1 0 8288 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_150
timestamp 1698175906
transform 1 0 9072 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_152
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_159
timestamp 1698175906
transform 1 0 9576 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_167
timestamp 1698175906
transform 1 0 10024 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_175
timestamp 1698175906
transform 1 0 10472 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_179
timestamp 1698175906
transform 1 0 10696 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_181
timestamp 1698175906
transform 1 0 10808 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_184
timestamp 1698175906
transform 1 0 10976 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_203
timestamp 1698175906
transform 1 0 12040 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_207
timestamp 1698175906
transform 1 0 12264 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698175906
transform 1 0 12376 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_245
timestamp 1698175906
transform 1 0 14392 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698175906
transform 1 0 16184 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 16296 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 18256 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 18704 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_126
timestamp 1698175906
transform 1 0 7728 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_158
timestamp 1698175906
transform 1 0 9520 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_173
timestamp 1698175906
transform 1 0 10360 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_240
timestamp 1698175906
transform 1 0 14112 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 14336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 2240 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 4032 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 4480 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_88
timestamp 1698175906
transform 1 0 5600 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_119
timestamp 1698175906
transform 1 0 7336 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_123
timestamp 1698175906
transform 1 0 7560 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_146
timestamp 1698175906
transform 1 0 8848 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_148
timestamp 1698175906
transform 1 0 8960 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_187
timestamp 1698175906
transform 1 0 11144 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_191
timestamp 1698175906
transform 1 0 11368 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_195
timestamp 1698175906
transform 1 0 11592 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_203
timestamp 1698175906
transform 1 0 12040 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698175906
transform 1 0 12264 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 12376 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_216
timestamp 1698175906
transform 1 0 12768 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_218
timestamp 1698175906
transform 1 0 12880 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_224
timestamp 1698175906
transform 1 0 13216 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_228
timestamp 1698175906
transform 1 0 13440 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_260
timestamp 1698175906
transform 1 0 15232 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 16128 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 2240 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 2464 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_169
timestamp 1698175906
transform 1 0 10136 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698175906
transform 1 0 10360 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_187
timestamp 1698175906
transform 1 0 11144 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_219
timestamp 1698175906
transform 1 0 12936 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_235
timestamp 1698175906
transform 1 0 13832 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698175906
transform 1 0 14280 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_104
timestamp 1698175906
transform 1 0 6496 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_120
timestamp 1698175906
transform 1 0 7392 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_132
timestamp 1698175906
transform 1 0 8064 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_150
timestamp 1698175906
transform 1 0 9072 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_156
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_188
timestamp 1698175906
transform 1 0 11200 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_204
timestamp 1698175906
transform 1 0 12096 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698175906
transform 1 0 12320 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_150
timestamp 1698175906
transform 1 0 9072 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_154
timestamp 1698175906
transform 1 0 9296 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 16128 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_165
timestamp 1698175906
transform 1 0 9912 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_169
timestamp 1698175906
transform 1 0 10136 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita62_24 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14392 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita62_25
timestamp 1698175906
transform 1 0 19992 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita62_26
timestamp 1698175906
transform -1 0 7336 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14616 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform -1 0 2240 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 10640 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 2240 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 10808 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 2240 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 18760 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 12096 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 10472 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 8456 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 18760 0 -1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform -1 0 2240 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 2240 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 9352 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 2240 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13440 400 13496 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 14112 0 14168 400 0 FreeSans 224 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 13104 0 13160 400 0 FreeSans 224 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 20600 10416 21000 10472 0 FreeSans 224 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 11424 0 11480 400 0 FreeSans 224 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 0 8064 400 8120 0 FreeSans 224 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 0 10416 400 10472 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 20600 10752 21000 10808 0 FreeSans 224 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 10752 20600 10808 21000 0 FreeSans 224 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 7056 0 7112 400 0 FreeSans 224 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 0 9408 400 9464 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 20600 12096 21000 12152 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 10752 0 10808 400 0 FreeSans 224 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 12096 20600 12152 21000 0 FreeSans 224 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 8064 0 8120 400 0 FreeSans 224 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 20600 9408 21000 9464 0 FreeSans 224 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 10416 0 10472 400 0 FreeSans 224 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 8400 20600 8456 21000 0 FreeSans 224 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 20600 7392 21000 7448 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 0 11088 400 11144 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 13104 400 13160 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 9744 20600 9800 21000 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 0 12768 400 12824 0 FreeSans 224 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 7140 11004 7140 11004 0 _000_
rlabel metal2 13244 7476 13244 7476 0 _001_
rlabel metal2 7364 13692 7364 13692 0 _002_
rlabel metal2 9268 6692 9268 6692 0 _003_
rlabel metal2 13356 9436 13356 9436 0 _004_
rlabel metal4 13692 8848 13692 8848 0 _005_
rlabel metal2 10220 7700 10220 7700 0 _006_
rlabel metal3 13230 10668 13230 10668 0 _007_
rlabel metal2 10556 7000 10556 7000 0 _008_
rlabel metal2 7112 7700 7112 7700 0 _009_
rlabel metal2 6076 10584 6076 10584 0 _010_
rlabel metal2 8988 13692 8988 13692 0 _011_
rlabel metal2 11284 12572 11284 12572 0 _012_
rlabel metal2 7756 7028 7756 7028 0 _013_
rlabel metal2 10052 12936 10052 12936 0 _014_
rlabel metal2 6692 9352 6692 9352 0 _015_
rlabel metal2 12908 12348 12908 12348 0 _016_
rlabel metal2 13244 12068 13244 12068 0 _017_
rlabel metal2 13020 7028 13020 7028 0 _018_
rlabel metal3 7532 12292 7532 12292 0 _019_
rlabel metal2 6916 12908 6916 12908 0 _020_
rlabel metal2 6692 11144 6692 11144 0 _021_
rlabel metal2 11256 9716 11256 9716 0 _022_
rlabel metal2 10164 8680 10164 8680 0 _023_
rlabel metal2 8876 7336 8876 7336 0 _024_
rlabel metal2 9436 7028 9436 7028 0 _025_
rlabel metal2 12824 10780 12824 10780 0 _026_
rlabel metal2 11704 11060 11704 11060 0 _027_
rlabel metal2 12852 9940 12852 9940 0 _028_
rlabel metal2 13412 9604 13412 9604 0 _029_
rlabel metal3 9828 9604 9828 9604 0 _030_
rlabel metal2 10976 8148 10976 8148 0 _031_
rlabel metal2 13972 9156 13972 9156 0 _032_
rlabel metal2 11060 7952 11060 7952 0 _033_
rlabel metal2 13748 10584 13748 10584 0 _034_
rlabel metal2 11676 11760 11676 11760 0 _035_
rlabel metal2 13104 10836 13104 10836 0 _036_
rlabel metal3 11032 7140 11032 7140 0 _037_
rlabel metal2 7252 8988 7252 8988 0 _038_
rlabel metal2 10808 7252 10808 7252 0 _039_
rlabel metal2 10640 7252 10640 7252 0 _040_
rlabel metal2 7140 8400 7140 8400 0 _041_
rlabel metal2 7924 9352 7924 9352 0 _042_
rlabel metal2 7504 8428 7504 8428 0 _043_
rlabel metal2 7028 10528 7028 10528 0 _044_
rlabel metal2 7476 9842 7476 9842 0 _045_
rlabel metal2 9324 13650 9324 13650 0 _046_
rlabel metal2 11116 12320 11116 12320 0 _047_
rlabel metal3 10584 11956 10584 11956 0 _048_
rlabel metal2 11452 12432 11452 12432 0 _049_
rlabel metal2 9184 8708 9184 8708 0 _050_
rlabel metal2 7476 7476 7476 7476 0 _051_
rlabel metal2 9996 12768 9996 12768 0 _052_
rlabel metal2 7252 9632 7252 9632 0 _053_
rlabel metal2 10472 12740 10472 12740 0 _054_
rlabel metal2 7196 9268 7196 9268 0 _055_
rlabel metal2 12740 12068 12740 12068 0 _056_
rlabel metal2 11956 9492 11956 9492 0 _057_
rlabel metal2 12936 11172 12936 11172 0 _058_
rlabel metal2 12628 11564 12628 11564 0 _059_
rlabel metal2 13468 11984 13468 11984 0 _060_
rlabel metal3 12824 7644 12824 7644 0 _061_
rlabel metal2 12348 7406 12348 7406 0 _062_
rlabel metal3 9548 9548 9548 9548 0 _063_
rlabel metal2 8484 9996 8484 9996 0 _064_
rlabel metal2 9324 9436 9324 9436 0 _065_
rlabel metal2 7448 10332 7448 10332 0 _066_
rlabel metal2 10836 11060 10836 11060 0 _067_
rlabel metal3 13076 11900 13076 11900 0 _068_
rlabel via2 10220 10780 10220 10780 0 _069_
rlabel metal2 10332 11060 10332 11060 0 _070_
rlabel metal2 8204 12180 8204 12180 0 _071_
rlabel via2 8876 9212 8876 9212 0 _072_
rlabel metal2 8988 10066 8988 10066 0 _073_
rlabel metal3 7448 12740 7448 12740 0 _074_
rlabel metal2 7700 12488 7700 12488 0 _075_
rlabel metal2 7028 12740 7028 12740 0 _076_
rlabel metal2 10668 10220 10668 10220 0 _077_
rlabel metal2 9324 11788 9324 11788 0 _078_
rlabel metal2 9380 11676 9380 11676 0 _079_
rlabel metal2 7084 11760 7084 11760 0 _080_
rlabel metal2 8064 9604 8064 9604 0 _081_
rlabel metal2 7980 9240 7980 9240 0 _082_
rlabel metal2 10164 10640 10164 10640 0 _083_
rlabel metal2 7980 10808 7980 10808 0 _084_
rlabel metal3 8372 8764 8372 8764 0 _085_
rlabel metal3 10052 11844 10052 11844 0 _086_
rlabel metal2 9940 11144 9940 11144 0 _087_
rlabel metal2 7364 10948 7364 10948 0 _088_
rlabel metal2 7196 11592 7196 11592 0 _089_
rlabel metal2 7476 11116 7476 11116 0 _090_
rlabel metal2 12348 9492 12348 9492 0 _091_
rlabel metal2 8708 7896 8708 7896 0 _092_
rlabel metal2 8960 9716 8960 9716 0 _093_
rlabel metal3 11088 8036 11088 8036 0 _094_
rlabel metal3 9212 7084 9212 7084 0 _095_
rlabel metal2 7588 9296 7588 9296 0 _096_
rlabel metal3 12236 10780 12236 10780 0 _097_
rlabel metal3 13356 9240 13356 9240 0 _098_
rlabel metal3 10612 7252 10612 7252 0 _099_
rlabel metal3 13580 7644 13580 7644 0 _100_
rlabel metal2 11564 9380 11564 9380 0 _101_
rlabel metal2 10668 11060 10668 11060 0 _102_
rlabel metal2 8120 13860 8120 13860 0 _103_
rlabel metal3 1239 13468 1239 13468 0 clk
rlabel metal2 11900 9380 11900 9380 0 clknet_0_clk
rlabel metal3 12516 6972 12516 6972 0 clknet_1_0__leaf_clk
rlabel metal2 7476 13104 7476 13104 0 clknet_1_1__leaf_clk
rlabel metal2 10332 9632 10332 9632 0 dut62.count\[0\]
rlabel metal2 11116 9268 11116 9268 0 dut62.count\[1\]
rlabel metal2 8260 9044 8260 9044 0 dut62.count\[2\]
rlabel metal2 8204 10808 8204 10808 0 dut62.count\[3\]
rlabel metal2 14084 6776 14084 6776 0 net1
rlabel metal2 14196 12124 14196 12124 0 net10
rlabel metal3 16464 11956 16464 11956 0 net11
rlabel metal2 11788 2982 11788 2982 0 net12
rlabel metal2 12404 12600 12404 12600 0 net13
rlabel metal3 8008 7140 8008 7140 0 net14
rlabel metal2 14756 8596 14756 8596 0 net15
rlabel metal2 14308 9632 14308 9632 0 net16
rlabel metal2 10556 3178 10556 3178 0 net17
rlabel metal2 8428 14770 8428 14770 0 net18
rlabel metal3 16576 7644 16576 7644 0 net19
rlabel metal2 14700 10752 14700 10752 0 net2
rlabel metal2 5628 10948 5628 10948 0 net20
rlabel metal2 2156 13384 2156 13384 0 net21
rlabel metal2 9744 13580 9744 13580 0 net22
rlabel metal2 6076 12712 6076 12712 0 net23
rlabel metal2 14140 1015 14140 1015 0 net24
rlabel metal2 20132 10920 20132 10920 0 net25
rlabel metal2 7084 1015 7084 1015 0 net26
rlabel metal2 11620 6776 11620 6776 0 net3
rlabel metal2 5964 8008 5964 8008 0 net4
rlabel metal2 10892 16240 10892 16240 0 net5
rlabel metal3 5992 10444 5992 10444 0 net6
rlabel metal2 11032 13524 11032 13524 0 net7
rlabel metal2 2156 9380 2156 9380 0 net8
rlabel metal3 13258 13188 13258 13188 0 net9
rlabel metal2 13132 1211 13132 1211 0 segm[10]
rlabel metal2 20020 10556 20020 10556 0 segm[11]
rlabel metal2 11452 1099 11452 1099 0 segm[12]
rlabel metal3 679 8092 679 8092 0 segm[13]
rlabel metal2 11116 19873 11116 19873 0 segm[1]
rlabel metal3 679 10444 679 10444 0 segm[2]
rlabel metal2 10780 19677 10780 19677 0 segm[4]
rlabel metal3 679 9436 679 9436 0 segm[6]
rlabel metal2 20020 12908 20020 12908 0 segm[7]
rlabel metal2 20020 12180 20020 12180 0 segm[8]
rlabel metal2 20020 11900 20020 11900 0 segm[9]
rlabel metal2 10780 1099 10780 1099 0 sel[0]
rlabel metal2 12124 19873 12124 19873 0 sel[10]
rlabel metal2 8092 1043 8092 1043 0 sel[11]
rlabel metal2 20020 8820 20020 8820 0 sel[1]
rlabel metal2 20020 9548 20020 9548 0 sel[2]
rlabel metal2 10444 1211 10444 1211 0 sel[3]
rlabel metal2 8428 19873 8428 19873 0 sel[4]
rlabel metal2 20020 7504 20020 7504 0 sel[5]
rlabel metal3 679 11116 679 11116 0 sel[6]
rlabel metal3 679 13132 679 13132 0 sel[7]
rlabel metal2 9884 18732 9884 18732 0 sel[8]
rlabel metal3 679 12796 679 12796 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
