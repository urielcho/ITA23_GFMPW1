magic
tech gf180mcuD
magscale 1 5
timestamp 1699642253
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9031 19137 9057 19143
rect 9031 19105 9057 19111
rect 11047 19137 11073 19143
rect 11047 19105 11073 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 8521 18999 8527 19025
rect 8553 18999 8559 19025
rect 10537 18999 10543 19025
rect 10569 18999 10575 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 3151 18969 3177 18975
rect 3151 18937 3177 18943
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 9199 18745 9225 18751
rect 9199 18713 9225 18719
rect 10711 18745 10737 18751
rect 10711 18713 10737 18719
rect 13119 18745 13145 18751
rect 13119 18713 13145 18719
rect 8857 18607 8863 18633
rect 8889 18607 8895 18633
rect 10201 18607 10207 18633
rect 10233 18607 10239 18633
rect 12609 18607 12615 18633
rect 12641 18607 12647 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 20119 18185 20145 18191
rect 20119 18153 20145 18159
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 8303 14041 8329 14047
rect 8303 14009 8329 14015
rect 8023 13985 8049 13991
rect 8023 13953 8049 13959
rect 8079 13929 8105 13935
rect 8079 13897 8105 13903
rect 8191 13929 8217 13935
rect 8191 13897 8217 13903
rect 8359 13929 8385 13935
rect 9081 13903 9087 13929
rect 9113 13903 9119 13929
rect 8359 13897 8385 13903
rect 8807 13873 8833 13879
rect 10711 13873 10737 13879
rect 9417 13847 9423 13873
rect 9449 13847 9455 13873
rect 10481 13847 10487 13873
rect 10513 13847 10519 13873
rect 8807 13841 8833 13847
rect 10711 13841 10737 13847
rect 8023 13817 8049 13823
rect 8023 13785 8049 13791
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 10319 13649 10345 13655
rect 10319 13617 10345 13623
rect 10711 13593 10737 13599
rect 20007 13593 20033 13599
rect 7401 13567 7407 13593
rect 7433 13567 7439 13593
rect 8465 13567 8471 13593
rect 8497 13567 8503 13593
rect 10089 13567 10095 13593
rect 10121 13567 10127 13593
rect 12497 13567 12503 13593
rect 12529 13567 12535 13593
rect 10711 13561 10737 13567
rect 20007 13561 20033 13567
rect 13903 13537 13929 13543
rect 7065 13511 7071 13537
rect 7097 13511 7103 13537
rect 8689 13511 8695 13537
rect 8721 13511 8727 13537
rect 11041 13511 11047 13537
rect 11073 13511 11079 13537
rect 18825 13511 18831 13537
rect 18857 13511 18863 13537
rect 13903 13505 13929 13511
rect 10263 13481 10289 13487
rect 13847 13481 13873 13487
rect 9025 13455 9031 13481
rect 9057 13455 9063 13481
rect 11433 13455 11439 13481
rect 11465 13455 11471 13481
rect 10263 13449 10289 13455
rect 13847 13449 13873 13455
rect 10319 13425 10345 13431
rect 10319 13393 10345 13399
rect 12727 13425 12753 13431
rect 12727 13393 12753 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 9535 13257 9561 13263
rect 9535 13225 9561 13231
rect 9927 13257 9953 13263
rect 9927 13225 9953 13231
rect 10039 13257 10065 13263
rect 10039 13225 10065 13231
rect 10207 13257 10233 13263
rect 10207 13225 10233 13231
rect 11887 13257 11913 13263
rect 11887 13225 11913 13231
rect 12167 13257 12193 13263
rect 12167 13225 12193 13231
rect 8751 13201 8777 13207
rect 8751 13169 8777 13175
rect 8807 13201 8833 13207
rect 8807 13169 8833 13175
rect 9647 13201 9673 13207
rect 9647 13169 9673 13175
rect 9871 13201 9897 13207
rect 9871 13169 9897 13175
rect 10151 13201 10177 13207
rect 10151 13169 10177 13175
rect 9703 13145 9729 13151
rect 6953 13119 6959 13145
rect 6985 13119 6991 13145
rect 9703 13113 9729 13119
rect 10319 13145 10345 13151
rect 14575 13145 14601 13151
rect 12273 13119 12279 13145
rect 12305 13119 12311 13145
rect 12889 13119 12895 13145
rect 12921 13119 12927 13145
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 10319 13113 10345 13119
rect 14575 13113 14601 13119
rect 7289 13063 7295 13089
rect 7321 13063 7327 13089
rect 8353 13063 8359 13089
rect 8385 13063 8391 13089
rect 13281 13063 13287 13089
rect 13313 13063 13319 13089
rect 14345 13063 14351 13089
rect 14377 13063 14383 13089
rect 8751 13033 8777 13039
rect 8751 13001 8777 13007
rect 11775 13033 11801 13039
rect 11775 13001 11801 13007
rect 11943 13033 11969 13039
rect 11943 13001 11969 13007
rect 12111 13033 12137 13039
rect 12111 13001 12137 13007
rect 20007 13033 20033 13039
rect 20007 13001 20033 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 14631 12809 14657 12815
rect 12609 12783 12615 12809
rect 12641 12783 12647 12809
rect 14289 12783 14295 12809
rect 14321 12783 14327 12809
rect 14631 12777 14657 12783
rect 7911 12753 7937 12759
rect 7911 12721 7937 12727
rect 8079 12753 8105 12759
rect 12447 12753 12473 12759
rect 10761 12727 10767 12753
rect 10793 12727 10799 12753
rect 8079 12721 8105 12727
rect 12447 12721 12473 12727
rect 12559 12753 12585 12759
rect 12665 12727 12671 12753
rect 12697 12727 12703 12753
rect 12833 12727 12839 12753
rect 12865 12727 12871 12753
rect 12559 12721 12585 12727
rect 10879 12697 10905 12703
rect 9249 12671 9255 12697
rect 9281 12671 9287 12697
rect 10879 12665 10905 12671
rect 10935 12697 10961 12703
rect 12335 12697 12361 12703
rect 11153 12671 11159 12697
rect 11185 12671 11191 12697
rect 13225 12671 13231 12697
rect 13257 12671 13263 12697
rect 10935 12665 10961 12671
rect 12335 12665 12361 12671
rect 8023 12641 8049 12647
rect 8023 12609 8049 12615
rect 8471 12641 8497 12647
rect 8471 12609 8497 12615
rect 9423 12641 9449 12647
rect 9423 12609 9449 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 12223 12473 12249 12479
rect 12223 12441 12249 12447
rect 13175 12473 13201 12479
rect 13175 12441 13201 12447
rect 13231 12473 13257 12479
rect 13231 12441 13257 12447
rect 14071 12417 14097 12423
rect 12833 12391 12839 12417
rect 12865 12391 12871 12417
rect 14071 12385 14097 12391
rect 12671 12361 12697 12367
rect 13287 12361 13313 12367
rect 14015 12361 14041 12367
rect 2137 12335 2143 12361
rect 2169 12335 2175 12361
rect 10593 12335 10599 12361
rect 10625 12335 10631 12361
rect 13057 12335 13063 12361
rect 13089 12335 13095 12361
rect 13393 12335 13399 12361
rect 13425 12335 13431 12361
rect 12671 12329 12697 12335
rect 13287 12329 13313 12335
rect 14015 12329 14041 12335
rect 10929 12279 10935 12305
rect 10961 12279 10967 12305
rect 11993 12279 11999 12305
rect 12025 12279 12031 12305
rect 967 12249 993 12255
rect 967 12217 993 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 9815 12081 9841 12087
rect 9815 12049 9841 12055
rect 10431 12081 10457 12087
rect 10431 12049 10457 12055
rect 10767 12081 10793 12087
rect 12497 12055 12503 12081
rect 12529 12055 12535 12081
rect 10767 12049 10793 12055
rect 6729 11999 6735 12025
rect 6761 11999 6767 12025
rect 10711 11969 10737 11975
rect 8129 11943 8135 11969
rect 8161 11943 8167 11969
rect 10711 11937 10737 11943
rect 10935 11969 10961 11975
rect 10935 11937 10961 11943
rect 11495 11969 11521 11975
rect 11495 11937 11521 11943
rect 11831 11969 11857 11975
rect 11831 11937 11857 11943
rect 12223 11969 12249 11975
rect 12223 11937 12249 11943
rect 12335 11969 12361 11975
rect 12335 11937 12361 11943
rect 8471 11913 8497 11919
rect 7793 11887 7799 11913
rect 7825 11887 7831 11913
rect 8471 11881 8497 11887
rect 9759 11913 9785 11919
rect 9759 11881 9785 11887
rect 10151 11913 10177 11919
rect 10151 11881 10177 11887
rect 11047 11913 11073 11919
rect 11047 11881 11073 11887
rect 11551 11913 11577 11919
rect 11551 11881 11577 11887
rect 8303 11857 8329 11863
rect 8303 11825 8329 11831
rect 8415 11857 8441 11863
rect 8415 11825 8441 11831
rect 8695 11857 8721 11863
rect 8695 11825 8721 11831
rect 9815 11857 9841 11863
rect 9815 11825 9841 11831
rect 10263 11857 10289 11863
rect 10263 11825 10289 11831
rect 10375 11857 10401 11863
rect 10375 11825 10401 11831
rect 10823 11857 10849 11863
rect 10823 11825 10849 11831
rect 11663 11857 11689 11863
rect 11663 11825 11689 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 7407 11689 7433 11695
rect 7407 11657 7433 11663
rect 7631 11689 7657 11695
rect 7631 11657 7657 11663
rect 7967 11689 7993 11695
rect 7967 11657 7993 11663
rect 9087 11689 9113 11695
rect 9087 11657 9113 11663
rect 9703 11689 9729 11695
rect 13231 11689 13257 11695
rect 12049 11663 12055 11689
rect 12081 11663 12087 11689
rect 9703 11657 9729 11663
rect 13231 11657 13257 11663
rect 6959 11633 6985 11639
rect 6959 11601 6985 11607
rect 7911 11633 7937 11639
rect 9591 11633 9617 11639
rect 11159 11633 11185 11639
rect 8913 11607 8919 11633
rect 8945 11607 8951 11633
rect 9977 11607 9983 11633
rect 10009 11607 10015 11633
rect 10313 11607 10319 11633
rect 10345 11607 10351 11633
rect 10873 11607 10879 11633
rect 10905 11607 10911 11633
rect 7911 11601 7937 11607
rect 9591 11601 9617 11607
rect 11159 11601 11185 11607
rect 7015 11577 7041 11583
rect 2137 11551 2143 11577
rect 2169 11551 2175 11577
rect 6729 11551 6735 11577
rect 6761 11551 6767 11577
rect 7015 11545 7041 11551
rect 8079 11577 8105 11583
rect 9535 11577 9561 11583
rect 8185 11551 8191 11577
rect 8217 11551 8223 11577
rect 8079 11545 8105 11551
rect 9535 11545 9561 11551
rect 9815 11577 9841 11583
rect 9815 11545 9841 11551
rect 10151 11577 10177 11583
rect 11887 11577 11913 11583
rect 10761 11551 10767 11577
rect 10793 11551 10799 11577
rect 11321 11551 11327 11577
rect 11353 11551 11359 11577
rect 13393 11551 13399 11577
rect 13425 11551 13431 11577
rect 10151 11545 10177 11551
rect 11887 11545 11913 11551
rect 7351 11521 7377 11527
rect 5273 11495 5279 11521
rect 5305 11495 5311 11521
rect 6337 11495 6343 11521
rect 6369 11495 6375 11521
rect 7351 11489 7377 11495
rect 8023 11521 8049 11527
rect 8023 11489 8049 11495
rect 9367 11521 9393 11527
rect 13785 11495 13791 11521
rect 13817 11495 13823 11521
rect 14849 11495 14855 11521
rect 14881 11495 14887 11521
rect 9367 11489 9393 11495
rect 967 11465 993 11471
rect 967 11433 993 11439
rect 6959 11465 6985 11471
rect 6959 11433 6985 11439
rect 11327 11465 11353 11471
rect 11327 11433 11353 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 967 11241 993 11247
rect 6791 11241 6817 11247
rect 4993 11215 4999 11241
rect 5025 11215 5031 11241
rect 967 11209 993 11215
rect 6791 11209 6817 11215
rect 7519 11241 7545 11247
rect 20007 11241 20033 11247
rect 7849 11215 7855 11241
rect 7881 11215 7887 11241
rect 8465 11215 8471 11241
rect 8497 11215 8503 11241
rect 9529 11215 9535 11241
rect 9561 11215 9567 11241
rect 13561 11215 13567 11241
rect 13593 11215 13599 11241
rect 7519 11209 7545 11215
rect 20007 11209 20033 11215
rect 7295 11185 7321 11191
rect 10095 11185 10121 11191
rect 2137 11159 2143 11185
rect 2169 11159 2175 11185
rect 6449 11159 6455 11185
rect 6481 11159 6487 11185
rect 7681 11159 7687 11185
rect 7713 11159 7719 11185
rect 8129 11159 8135 11185
rect 8161 11159 8167 11185
rect 7295 11153 7321 11159
rect 10095 11153 10121 11159
rect 10655 11185 10681 11191
rect 11831 11185 11857 11191
rect 10985 11159 10991 11185
rect 11017 11159 11023 11185
rect 11377 11159 11383 11185
rect 11409 11159 11415 11185
rect 11657 11159 11663 11185
rect 11689 11159 11695 11185
rect 13617 11159 13623 11185
rect 13649 11159 13655 11185
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 10655 11153 10681 11159
rect 11831 11153 11857 11159
rect 6959 11129 6985 11135
rect 6057 11103 6063 11129
rect 6089 11103 6095 11129
rect 6959 11097 6985 11103
rect 7239 11129 7265 11135
rect 7239 11097 7265 11103
rect 9927 11129 9953 11135
rect 9927 11097 9953 11103
rect 10263 11129 10289 11135
rect 10263 11097 10289 11103
rect 10375 11129 10401 11135
rect 13287 11129 13313 11135
rect 10929 11103 10935 11129
rect 10961 11103 10967 11129
rect 11265 11103 11271 11129
rect 11297 11103 11303 11129
rect 10375 11097 10401 11103
rect 13287 11097 13313 11103
rect 14631 11129 14657 11135
rect 14631 11097 14657 11103
rect 6735 11073 6761 11079
rect 6735 11041 6761 11047
rect 6847 11073 6873 11079
rect 6847 11041 6873 11047
rect 7127 11073 7153 11079
rect 7127 11041 7153 11047
rect 7799 11073 7825 11079
rect 7799 11041 7825 11047
rect 7911 11073 7937 11079
rect 7911 11041 7937 11047
rect 9815 11073 9841 11079
rect 9815 11041 9841 11047
rect 9871 11073 9897 11079
rect 9871 11041 9897 11047
rect 10207 11073 10233 11079
rect 10207 11041 10233 11047
rect 10711 11073 10737 11079
rect 13399 11073 13425 11079
rect 11993 11047 11999 11073
rect 12025 11047 12031 11073
rect 10711 11041 10737 11047
rect 13399 11041 13425 11047
rect 13511 11073 13537 11079
rect 13511 11041 13537 11047
rect 14575 11073 14601 11079
rect 14575 11041 14601 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 6399 10905 6425 10911
rect 6399 10873 6425 10879
rect 7687 10905 7713 10911
rect 7687 10873 7713 10879
rect 7855 10905 7881 10911
rect 7855 10873 7881 10879
rect 11551 10905 11577 10911
rect 11551 10873 11577 10879
rect 12727 10905 12753 10911
rect 12727 10873 12753 10879
rect 13119 10905 13145 10911
rect 13119 10873 13145 10879
rect 6847 10849 6873 10855
rect 6847 10817 6873 10823
rect 7183 10849 7209 10855
rect 7183 10817 7209 10823
rect 7239 10849 7265 10855
rect 7239 10817 7265 10823
rect 7743 10849 7769 10855
rect 11831 10849 11857 10855
rect 9361 10823 9367 10849
rect 9393 10823 9399 10849
rect 7743 10817 7769 10823
rect 11831 10817 11857 10823
rect 11943 10849 11969 10855
rect 11943 10817 11969 10823
rect 6567 10793 6593 10799
rect 6567 10761 6593 10767
rect 6735 10793 6761 10799
rect 6735 10761 6761 10767
rect 7071 10793 7097 10799
rect 7071 10761 7097 10767
rect 8023 10793 8049 10799
rect 11999 10793 12025 10799
rect 11153 10767 11159 10793
rect 11185 10767 11191 10793
rect 11657 10767 11663 10793
rect 11689 10767 11695 10793
rect 8023 10761 8049 10767
rect 11999 10761 12025 10767
rect 12055 10793 12081 10799
rect 12055 10761 12081 10767
rect 12111 10793 12137 10799
rect 13007 10793 13033 10799
rect 12889 10767 12895 10793
rect 12921 10767 12927 10793
rect 13225 10767 13231 10793
rect 13257 10767 13263 10793
rect 13449 10767 13455 10793
rect 13481 10767 13487 10793
rect 18825 10767 18831 10793
rect 18857 10767 18863 10793
rect 12111 10761 12137 10767
rect 13007 10761 13033 10767
rect 13063 10737 13089 10743
rect 20007 10737 20033 10743
rect 13785 10711 13791 10737
rect 13817 10711 13823 10737
rect 14849 10711 14855 10737
rect 14881 10711 14887 10737
rect 13063 10705 13089 10711
rect 20007 10705 20033 10711
rect 6455 10681 6481 10687
rect 6455 10649 6481 10655
rect 11495 10681 11521 10687
rect 11495 10649 11521 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 7799 10513 7825 10519
rect 7799 10481 7825 10487
rect 10655 10513 10681 10519
rect 10655 10481 10681 10487
rect 14575 10513 14601 10519
rect 14575 10481 14601 10487
rect 14015 10457 14041 10463
rect 8185 10431 8191 10457
rect 8217 10431 8223 10457
rect 13449 10431 13455 10457
rect 13481 10431 13487 10457
rect 14015 10425 14041 10431
rect 8303 10401 8329 10407
rect 7513 10375 7519 10401
rect 7545 10375 7551 10401
rect 8303 10369 8329 10375
rect 8471 10401 8497 10407
rect 8471 10369 8497 10375
rect 8639 10401 8665 10407
rect 8639 10369 8665 10375
rect 8695 10401 8721 10407
rect 8695 10369 8721 10375
rect 8863 10401 8889 10407
rect 8863 10369 8889 10375
rect 10207 10401 10233 10407
rect 10207 10369 10233 10375
rect 10823 10401 10849 10407
rect 11153 10375 11159 10401
rect 11185 10375 11191 10401
rect 10823 10369 10849 10375
rect 7407 10345 7433 10351
rect 7407 10313 7433 10319
rect 7855 10345 7881 10351
rect 7855 10313 7881 10319
rect 8191 10345 8217 10351
rect 8191 10313 8217 10319
rect 8527 10345 8553 10351
rect 8527 10313 8553 10319
rect 8807 10345 8833 10351
rect 9423 10345 9449 10351
rect 9025 10319 9031 10345
rect 9057 10319 9063 10345
rect 8807 10313 8833 10319
rect 9423 10313 9449 10319
rect 9535 10345 9561 10351
rect 10935 10345 10961 10351
rect 9865 10319 9871 10345
rect 9897 10319 9903 10345
rect 9977 10319 9983 10345
rect 10009 10319 10015 10345
rect 9535 10313 9561 10319
rect 10935 10313 10961 10319
rect 14631 10345 14657 10351
rect 14631 10313 14657 10319
rect 9199 10289 9225 10295
rect 9199 10257 9225 10263
rect 9479 10289 9505 10295
rect 10201 10263 10207 10289
rect 10233 10263 10239 10289
rect 9479 10257 9505 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 9255 10121 9281 10127
rect 13393 10095 13399 10121
rect 13425 10095 13431 10121
rect 9255 10089 9281 10095
rect 8023 10065 8049 10071
rect 7289 10039 7295 10065
rect 7321 10039 7327 10065
rect 8023 10033 8049 10039
rect 8135 10065 8161 10071
rect 12615 10065 12641 10071
rect 11153 10039 11159 10065
rect 11185 10039 11191 10065
rect 8135 10033 8161 10039
rect 12615 10033 12641 10039
rect 12839 10065 12865 10071
rect 12839 10033 12865 10039
rect 7127 10009 7153 10015
rect 7127 9977 7153 9983
rect 7463 10009 7489 10015
rect 7463 9977 7489 9983
rect 7743 10009 7769 10015
rect 7743 9977 7769 9983
rect 8807 10009 8833 10015
rect 12727 10009 12753 10015
rect 9417 9983 9423 10009
rect 9449 9983 9455 10009
rect 8807 9977 8833 9983
rect 12727 9977 12753 9983
rect 12895 10009 12921 10015
rect 12895 9977 12921 9983
rect 13231 10009 13257 10015
rect 13561 9983 13567 10009
rect 13593 9983 13599 10009
rect 18825 9983 18831 10009
rect 18857 9983 18863 10009
rect 13231 9977 13257 9983
rect 6567 9953 6593 9959
rect 6567 9921 6593 9927
rect 8079 9953 8105 9959
rect 13119 9953 13145 9959
rect 9025 9927 9031 9953
rect 9057 9927 9063 9953
rect 13953 9927 13959 9953
rect 13985 9927 13991 9953
rect 15017 9927 15023 9953
rect 15049 9927 15055 9953
rect 8079 9921 8105 9927
rect 13119 9921 13145 9927
rect 12895 9897 12921 9903
rect 12895 9865 12921 9871
rect 20007 9897 20033 9903
rect 20007 9865 20033 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 12105 9703 12111 9729
rect 12137 9703 12143 9729
rect 20007 9673 20033 9679
rect 5385 9647 5391 9673
rect 5417 9647 5423 9673
rect 6449 9647 6455 9673
rect 6481 9647 6487 9673
rect 13785 9647 13791 9673
rect 13817 9647 13823 9673
rect 20007 9641 20033 9647
rect 7519 9617 7545 9623
rect 5049 9591 5055 9617
rect 5081 9591 5087 9617
rect 7401 9591 7407 9617
rect 7433 9591 7439 9617
rect 7519 9585 7545 9591
rect 9143 9617 9169 9623
rect 9143 9585 9169 9591
rect 9759 9617 9785 9623
rect 9759 9585 9785 9591
rect 10039 9617 10065 9623
rect 10039 9585 10065 9591
rect 10095 9617 10121 9623
rect 11495 9617 11521 9623
rect 13175 9617 13201 9623
rect 14183 9617 14209 9623
rect 10985 9591 10991 9617
rect 11017 9591 11023 9617
rect 11713 9591 11719 9617
rect 11745 9591 11751 9617
rect 13505 9591 13511 9617
rect 13537 9591 13543 9617
rect 10095 9585 10121 9591
rect 11495 9585 11521 9591
rect 13175 9585 13201 9591
rect 14183 9585 14209 9591
rect 14239 9617 14265 9623
rect 18937 9591 18943 9617
rect 18969 9591 18975 9617
rect 14239 9585 14265 9591
rect 6735 9561 6761 9567
rect 6735 9529 6761 9535
rect 6903 9561 6929 9567
rect 6903 9529 6929 9535
rect 7071 9561 7097 9567
rect 7071 9529 7097 9535
rect 7911 9561 7937 9567
rect 7911 9529 7937 9535
rect 8079 9561 8105 9567
rect 8079 9529 8105 9535
rect 8303 9561 8329 9567
rect 8303 9529 8329 9535
rect 9255 9561 9281 9567
rect 9255 9529 9281 9535
rect 9311 9561 9337 9567
rect 9311 9529 9337 9535
rect 9983 9561 10009 9567
rect 13735 9561 13761 9567
rect 10929 9535 10935 9561
rect 10961 9535 10967 9561
rect 12665 9535 12671 9561
rect 12697 9535 12703 9561
rect 12833 9535 12839 9561
rect 12865 9535 12871 9561
rect 9983 9529 10009 9535
rect 13735 9529 13761 9535
rect 14015 9561 14041 9567
rect 14015 9529 14041 9535
rect 8359 9505 8385 9511
rect 8359 9473 8385 9479
rect 9479 9505 9505 9511
rect 12503 9505 12529 9511
rect 10313 9479 10319 9505
rect 10345 9479 10351 9505
rect 9479 9473 9505 9479
rect 12503 9473 12529 9479
rect 13007 9505 13033 9511
rect 13007 9473 13033 9479
rect 13343 9505 13369 9511
rect 13343 9473 13369 9479
rect 13623 9505 13649 9511
rect 13623 9473 13649 9479
rect 13791 9505 13817 9511
rect 13791 9473 13817 9479
rect 14071 9505 14097 9511
rect 14071 9473 14097 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 9647 9337 9673 9343
rect 7233 9311 7239 9337
rect 7265 9311 7271 9337
rect 7569 9311 7575 9337
rect 7601 9311 7607 9337
rect 9647 9305 9673 9311
rect 9983 9337 10009 9343
rect 9983 9305 10009 9311
rect 10095 9337 10121 9343
rect 12839 9337 12865 9343
rect 11937 9311 11943 9337
rect 11969 9311 11975 9337
rect 10095 9305 10121 9311
rect 12839 9305 12865 9311
rect 13455 9337 13481 9343
rect 13455 9305 13481 9311
rect 11327 9281 11353 9287
rect 7905 9255 7911 9281
rect 7937 9255 7943 9281
rect 11327 9249 11353 9255
rect 12783 9281 12809 9287
rect 12783 9249 12809 9255
rect 13287 9281 13313 9287
rect 13287 9249 13313 9255
rect 13343 9281 13369 9287
rect 13953 9255 13959 9281
rect 13985 9255 13991 9281
rect 15353 9255 15359 9281
rect 15385 9255 15391 9281
rect 13343 9249 13369 9255
rect 7407 9225 7433 9231
rect 9591 9225 9617 9231
rect 11159 9225 11185 9231
rect 5273 9199 5279 9225
rect 5305 9199 5311 9225
rect 7121 9199 7127 9225
rect 7153 9199 7159 9225
rect 8129 9199 8135 9225
rect 8161 9199 8167 9225
rect 8353 9199 8359 9225
rect 8385 9199 8391 9225
rect 9865 9199 9871 9225
rect 9897 9199 9903 9225
rect 10201 9199 10207 9225
rect 10233 9199 10239 9225
rect 10929 9199 10935 9225
rect 10961 9199 10967 9225
rect 13561 9199 13567 9225
rect 13593 9199 13599 9225
rect 15241 9199 15247 9225
rect 15273 9199 15279 9225
rect 18825 9199 18831 9225
rect 18857 9199 18863 9225
rect 7407 9193 7433 9199
rect 9591 9193 9617 9199
rect 11159 9193 11185 9199
rect 6903 9169 6929 9175
rect 10039 9169 10065 9175
rect 11663 9169 11689 9175
rect 5609 9143 5615 9169
rect 5641 9143 5647 9169
rect 6673 9143 6679 9169
rect 6705 9143 6711 9169
rect 8185 9143 8191 9169
rect 8217 9143 8223 9169
rect 11041 9143 11047 9169
rect 11073 9143 11079 9169
rect 6903 9137 6929 9143
rect 10039 9137 10065 9143
rect 11663 9137 11689 9143
rect 13119 9169 13145 9175
rect 15017 9143 15023 9169
rect 15049 9143 15055 9169
rect 13119 9137 13145 9143
rect 11775 9113 11801 9119
rect 11775 9081 11801 9087
rect 12839 9113 12865 9119
rect 12839 9081 12865 9087
rect 20007 9113 20033 9119
rect 20007 9081 20033 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 7911 8945 7937 8951
rect 7911 8913 7937 8919
rect 9647 8945 9673 8951
rect 9647 8913 9673 8919
rect 10655 8945 10681 8951
rect 10655 8913 10681 8919
rect 10711 8945 10737 8951
rect 10711 8913 10737 8919
rect 10823 8945 10849 8951
rect 10823 8913 10849 8919
rect 10879 8945 10905 8951
rect 10879 8913 10905 8919
rect 11607 8945 11633 8951
rect 11607 8913 11633 8919
rect 9535 8889 9561 8895
rect 13847 8889 13873 8895
rect 11489 8863 11495 8889
rect 11521 8863 11527 8889
rect 9535 8857 9561 8863
rect 13847 8857 13873 8863
rect 20007 8889 20033 8895
rect 20007 8857 20033 8863
rect 9927 8833 9953 8839
rect 12615 8833 12641 8839
rect 10145 8807 10151 8833
rect 10177 8807 10183 8833
rect 11433 8807 11439 8833
rect 11465 8807 11471 8833
rect 9927 8801 9953 8807
rect 12615 8801 12641 8807
rect 12839 8833 12865 8839
rect 12839 8801 12865 8807
rect 12951 8833 12977 8839
rect 12951 8801 12977 8807
rect 13735 8833 13761 8839
rect 13735 8801 13761 8807
rect 13903 8833 13929 8839
rect 13903 8801 13929 8807
rect 14071 8833 14097 8839
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 14071 8801 14097 8807
rect 9255 8777 9281 8783
rect 9255 8745 9281 8751
rect 9367 8777 9393 8783
rect 9367 8745 9393 8751
rect 9423 8777 9449 8783
rect 9423 8745 9449 8751
rect 9871 8777 9897 8783
rect 9871 8745 9897 8751
rect 7799 8721 7825 8727
rect 7799 8689 7825 8695
rect 7855 8721 7881 8727
rect 7855 8689 7881 8695
rect 8415 8721 8441 8727
rect 8415 8689 8441 8695
rect 12783 8721 12809 8727
rect 12783 8689 12809 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 9031 8553 9057 8559
rect 9031 8521 9057 8527
rect 10319 8553 10345 8559
rect 10319 8521 10345 8527
rect 12223 8553 12249 8559
rect 12223 8521 12249 8527
rect 12335 8553 12361 8559
rect 12335 8521 12361 8527
rect 8863 8497 8889 8503
rect 7233 8471 7239 8497
rect 7265 8471 7271 8497
rect 8863 8465 8889 8471
rect 8919 8497 8945 8503
rect 8919 8465 8945 8471
rect 11383 8497 11409 8503
rect 11383 8465 11409 8471
rect 11495 8497 11521 8503
rect 11495 8465 11521 8471
rect 12111 8497 12137 8503
rect 13001 8471 13007 8497
rect 13033 8471 13039 8497
rect 12111 8465 12137 8471
rect 9759 8441 9785 8447
rect 14295 8441 14321 8447
rect 6897 8415 6903 8441
rect 6929 8415 6935 8441
rect 9529 8415 9535 8441
rect 9561 8415 9567 8441
rect 12665 8415 12671 8441
rect 12697 8415 12703 8441
rect 9759 8409 9785 8415
rect 14295 8409 14321 8415
rect 10207 8385 10233 8391
rect 8297 8359 8303 8385
rect 8329 8359 8335 8385
rect 10207 8353 10233 8359
rect 12391 8385 12417 8391
rect 14065 8359 14071 8385
rect 14097 8359 14103 8385
rect 12391 8353 12417 8359
rect 10375 8329 10401 8335
rect 10375 8297 10401 8303
rect 11551 8329 11577 8335
rect 11551 8297 11577 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 12167 8105 12193 8111
rect 7681 8079 7687 8105
rect 7713 8079 7719 8105
rect 8745 8079 8751 8105
rect 8777 8079 8783 8105
rect 12167 8073 12193 8079
rect 11551 8049 11577 8055
rect 11943 8049 11969 8055
rect 7345 8023 7351 8049
rect 7377 8023 7383 8049
rect 9865 8023 9871 8049
rect 9897 8023 9903 8049
rect 11769 8023 11775 8049
rect 11801 8023 11807 8049
rect 12105 8023 12111 8049
rect 12137 8023 12143 8049
rect 11551 8017 11577 8023
rect 11943 8017 11969 8023
rect 11383 7993 11409 7999
rect 9977 7967 9983 7993
rect 10009 7967 10015 7993
rect 11383 7961 11409 7967
rect 11439 7993 11465 7999
rect 11439 7961 11465 7967
rect 11663 7993 11689 7999
rect 11663 7961 11689 7967
rect 8975 7937 9001 7943
rect 8975 7905 9001 7911
rect 11607 7937 11633 7943
rect 11607 7905 11633 7911
rect 12223 7937 12249 7943
rect 12223 7905 12249 7911
rect 12335 7937 12361 7943
rect 12335 7905 12361 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 9535 7713 9561 7719
rect 9535 7681 9561 7687
rect 9703 7657 9729 7663
rect 10767 7657 10793 7663
rect 9809 7631 9815 7657
rect 9841 7631 9847 7657
rect 9703 7625 9729 7631
rect 10767 7625 10793 7631
rect 9591 7601 9617 7607
rect 9591 7569 9617 7575
rect 10655 7601 10681 7607
rect 10655 7569 10681 7575
rect 10599 7545 10625 7551
rect 9809 7519 9815 7545
rect 9841 7519 9847 7545
rect 10599 7513 10625 7519
rect 10823 7545 10849 7551
rect 10823 7513 10849 7519
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 9759 7377 9785 7383
rect 9759 7345 9785 7351
rect 10207 7377 10233 7383
rect 10207 7345 10233 7351
rect 10711 7321 10737 7327
rect 8521 7295 8527 7321
rect 8553 7295 8559 7321
rect 9585 7295 9591 7321
rect 9617 7295 9623 7321
rect 11881 7295 11887 7321
rect 11913 7295 11919 7321
rect 12945 7295 12951 7321
rect 12977 7295 12983 7321
rect 10711 7289 10737 7295
rect 10767 7265 10793 7271
rect 8185 7239 8191 7265
rect 8217 7239 8223 7265
rect 10369 7239 10375 7265
rect 10401 7239 10407 7265
rect 10767 7233 10793 7239
rect 10935 7265 10961 7271
rect 11489 7239 11495 7265
rect 11521 7239 11527 7265
rect 10935 7233 10961 7239
rect 9815 7209 9841 7215
rect 9815 7177 9841 7183
rect 10655 7209 10681 7215
rect 10655 7177 10681 7183
rect 10039 7153 10065 7159
rect 10039 7121 10065 7127
rect 10263 7153 10289 7159
rect 10263 7121 10289 7127
rect 13175 7153 13201 7159
rect 13175 7121 13201 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 9983 6985 10009 6991
rect 9983 6953 10009 6959
rect 9703 6929 9729 6935
rect 9703 6897 9729 6903
rect 10039 6929 10065 6935
rect 10817 6903 10823 6929
rect 10849 6903 10855 6929
rect 12329 6903 12335 6929
rect 12361 6903 12367 6929
rect 10039 6897 10065 6903
rect 9871 6873 9897 6879
rect 12167 6873 12193 6879
rect 10257 6847 10263 6873
rect 10289 6847 10295 6873
rect 10481 6847 10487 6873
rect 10513 6847 10519 6873
rect 9871 6841 9897 6847
rect 12167 6841 12193 6847
rect 9647 6817 9673 6823
rect 9647 6785 9673 6791
rect 9927 6817 9953 6823
rect 11937 6791 11943 6817
rect 11969 6791 11975 6817
rect 9927 6785 9953 6791
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 10711 6537 10737 6543
rect 9305 6511 9311 6537
rect 9337 6511 9343 6537
rect 10369 6511 10375 6537
rect 10401 6511 10407 6537
rect 10711 6505 10737 6511
rect 12167 6537 12193 6543
rect 12167 6505 12193 6511
rect 8969 6455 8975 6481
rect 9001 6455 9007 6481
rect 11601 6455 11607 6481
rect 11633 6455 11639 6481
rect 11713 6343 11719 6369
rect 11745 6343 11751 6369
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 12391 2617 12417 2623
rect 12391 2585 12417 2591
rect 11881 2535 11887 2561
rect 11913 2535 11919 2561
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 8857 2143 8863 2169
rect 8889 2143 8895 2169
rect 10537 2143 10543 2169
rect 10569 2143 10575 2169
rect 12665 2143 12671 2169
rect 12697 2143 12703 2169
rect 9367 2057 9393 2063
rect 9367 2025 9393 2031
rect 11047 2057 11073 2063
rect 11047 2025 11073 2031
rect 13119 2057 13145 2063
rect 13119 2025 13145 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 9865 1751 9871 1777
rect 9897 1751 9903 1777
rect 11769 1751 11775 1777
rect 11801 1751 11807 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 11097 1695 11103 1721
rect 11129 1695 11135 1721
rect 9591 1665 9617 1671
rect 9591 1633 9617 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9031 19111 9057 19137
rect 11047 19111 11073 19137
rect 12783 19111 12809 19137
rect 8527 18999 8553 19025
rect 10543 18999 10569 19025
rect 12279 18999 12305 19025
rect 3151 18943 3177 18969
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 9199 18719 9225 18745
rect 10711 18719 10737 18745
rect 13119 18719 13145 18745
rect 8863 18607 8889 18633
rect 10207 18607 10233 18633
rect 12615 18607 12641 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 20119 18159 20145 18185
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 8303 14015 8329 14041
rect 8023 13959 8049 13985
rect 8079 13903 8105 13929
rect 8191 13903 8217 13929
rect 8359 13903 8385 13929
rect 9087 13903 9113 13929
rect 8807 13847 8833 13873
rect 9423 13847 9449 13873
rect 10487 13847 10513 13873
rect 10711 13847 10737 13873
rect 8023 13791 8049 13817
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 10319 13623 10345 13649
rect 7407 13567 7433 13593
rect 8471 13567 8497 13593
rect 10095 13567 10121 13593
rect 10711 13567 10737 13593
rect 12503 13567 12529 13593
rect 20007 13567 20033 13593
rect 7071 13511 7097 13537
rect 8695 13511 8721 13537
rect 11047 13511 11073 13537
rect 13903 13511 13929 13537
rect 18831 13511 18857 13537
rect 9031 13455 9057 13481
rect 10263 13455 10289 13481
rect 11439 13455 11465 13481
rect 13847 13455 13873 13481
rect 10319 13399 10345 13425
rect 12727 13399 12753 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 9535 13231 9561 13257
rect 9927 13231 9953 13257
rect 10039 13231 10065 13257
rect 10207 13231 10233 13257
rect 11887 13231 11913 13257
rect 12167 13231 12193 13257
rect 8751 13175 8777 13201
rect 8807 13175 8833 13201
rect 9647 13175 9673 13201
rect 9871 13175 9897 13201
rect 10151 13175 10177 13201
rect 6959 13119 6985 13145
rect 9703 13119 9729 13145
rect 10319 13119 10345 13145
rect 12279 13119 12305 13145
rect 12895 13119 12921 13145
rect 14575 13119 14601 13145
rect 18831 13119 18857 13145
rect 7295 13063 7321 13089
rect 8359 13063 8385 13089
rect 13287 13063 13313 13089
rect 14351 13063 14377 13089
rect 8751 13007 8777 13033
rect 11775 13007 11801 13033
rect 11943 13007 11969 13033
rect 12111 13007 12137 13033
rect 20007 13007 20033 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 12615 12783 12641 12809
rect 14295 12783 14321 12809
rect 14631 12783 14657 12809
rect 7911 12727 7937 12753
rect 8079 12727 8105 12753
rect 10767 12727 10793 12753
rect 12447 12727 12473 12753
rect 12559 12727 12585 12753
rect 12671 12727 12697 12753
rect 12839 12727 12865 12753
rect 9255 12671 9281 12697
rect 10879 12671 10905 12697
rect 10935 12671 10961 12697
rect 11159 12671 11185 12697
rect 12335 12671 12361 12697
rect 13231 12671 13257 12697
rect 8023 12615 8049 12641
rect 8471 12615 8497 12641
rect 9423 12615 9449 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 12223 12447 12249 12473
rect 13175 12447 13201 12473
rect 13231 12447 13257 12473
rect 12839 12391 12865 12417
rect 14071 12391 14097 12417
rect 2143 12335 2169 12361
rect 10599 12335 10625 12361
rect 12671 12335 12697 12361
rect 13063 12335 13089 12361
rect 13287 12335 13313 12361
rect 13399 12335 13425 12361
rect 14015 12335 14041 12361
rect 10935 12279 10961 12305
rect 11999 12279 12025 12305
rect 967 12223 993 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 9815 12055 9841 12081
rect 10431 12055 10457 12081
rect 10767 12055 10793 12081
rect 12503 12055 12529 12081
rect 6735 11999 6761 12025
rect 8135 11943 8161 11969
rect 10711 11943 10737 11969
rect 10935 11943 10961 11969
rect 11495 11943 11521 11969
rect 11831 11943 11857 11969
rect 12223 11943 12249 11969
rect 12335 11943 12361 11969
rect 7799 11887 7825 11913
rect 8471 11887 8497 11913
rect 9759 11887 9785 11913
rect 10151 11887 10177 11913
rect 11047 11887 11073 11913
rect 11551 11887 11577 11913
rect 8303 11831 8329 11857
rect 8415 11831 8441 11857
rect 8695 11831 8721 11857
rect 9815 11831 9841 11857
rect 10263 11831 10289 11857
rect 10375 11831 10401 11857
rect 10823 11831 10849 11857
rect 11663 11831 11689 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 7407 11663 7433 11689
rect 7631 11663 7657 11689
rect 7967 11663 7993 11689
rect 9087 11663 9113 11689
rect 9703 11663 9729 11689
rect 12055 11663 12081 11689
rect 13231 11663 13257 11689
rect 6959 11607 6985 11633
rect 7911 11607 7937 11633
rect 8919 11607 8945 11633
rect 9591 11607 9617 11633
rect 9983 11607 10009 11633
rect 10319 11607 10345 11633
rect 10879 11607 10905 11633
rect 11159 11607 11185 11633
rect 2143 11551 2169 11577
rect 6735 11551 6761 11577
rect 7015 11551 7041 11577
rect 8079 11551 8105 11577
rect 8191 11551 8217 11577
rect 9535 11551 9561 11577
rect 9815 11551 9841 11577
rect 10151 11551 10177 11577
rect 10767 11551 10793 11577
rect 11327 11551 11353 11577
rect 11887 11551 11913 11577
rect 13399 11551 13425 11577
rect 5279 11495 5305 11521
rect 6343 11495 6369 11521
rect 7351 11495 7377 11521
rect 8023 11495 8049 11521
rect 9367 11495 9393 11521
rect 13791 11495 13817 11521
rect 14855 11495 14881 11521
rect 967 11439 993 11465
rect 6959 11439 6985 11465
rect 11327 11439 11353 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 967 11215 993 11241
rect 4999 11215 5025 11241
rect 6791 11215 6817 11241
rect 7519 11215 7545 11241
rect 7855 11215 7881 11241
rect 8471 11215 8497 11241
rect 9535 11215 9561 11241
rect 13567 11215 13593 11241
rect 20007 11215 20033 11241
rect 2143 11159 2169 11185
rect 6455 11159 6481 11185
rect 7295 11159 7321 11185
rect 7687 11159 7713 11185
rect 8135 11159 8161 11185
rect 10095 11159 10121 11185
rect 10655 11159 10681 11185
rect 10991 11159 11017 11185
rect 11383 11159 11409 11185
rect 11663 11159 11689 11185
rect 11831 11159 11857 11185
rect 13623 11159 13649 11185
rect 18831 11159 18857 11185
rect 6063 11103 6089 11129
rect 6959 11103 6985 11129
rect 7239 11103 7265 11129
rect 9927 11103 9953 11129
rect 10263 11103 10289 11129
rect 10375 11103 10401 11129
rect 10935 11103 10961 11129
rect 11271 11103 11297 11129
rect 13287 11103 13313 11129
rect 14631 11103 14657 11129
rect 6735 11047 6761 11073
rect 6847 11047 6873 11073
rect 7127 11047 7153 11073
rect 7799 11047 7825 11073
rect 7911 11047 7937 11073
rect 9815 11047 9841 11073
rect 9871 11047 9897 11073
rect 10207 11047 10233 11073
rect 10711 11047 10737 11073
rect 11999 11047 12025 11073
rect 13399 11047 13425 11073
rect 13511 11047 13537 11073
rect 14575 11047 14601 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 6399 10879 6425 10905
rect 7687 10879 7713 10905
rect 7855 10879 7881 10905
rect 11551 10879 11577 10905
rect 12727 10879 12753 10905
rect 13119 10879 13145 10905
rect 6847 10823 6873 10849
rect 7183 10823 7209 10849
rect 7239 10823 7265 10849
rect 7743 10823 7769 10849
rect 9367 10823 9393 10849
rect 11831 10823 11857 10849
rect 11943 10823 11969 10849
rect 6567 10767 6593 10793
rect 6735 10767 6761 10793
rect 7071 10767 7097 10793
rect 8023 10767 8049 10793
rect 11159 10767 11185 10793
rect 11663 10767 11689 10793
rect 11999 10767 12025 10793
rect 12055 10767 12081 10793
rect 12111 10767 12137 10793
rect 12895 10767 12921 10793
rect 13007 10767 13033 10793
rect 13231 10767 13257 10793
rect 13455 10767 13481 10793
rect 18831 10767 18857 10793
rect 13063 10711 13089 10737
rect 13791 10711 13817 10737
rect 14855 10711 14881 10737
rect 20007 10711 20033 10737
rect 6455 10655 6481 10681
rect 11495 10655 11521 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 7799 10487 7825 10513
rect 10655 10487 10681 10513
rect 14575 10487 14601 10513
rect 8191 10431 8217 10457
rect 13455 10431 13481 10457
rect 14015 10431 14041 10457
rect 7519 10375 7545 10401
rect 8303 10375 8329 10401
rect 8471 10375 8497 10401
rect 8639 10375 8665 10401
rect 8695 10375 8721 10401
rect 8863 10375 8889 10401
rect 10207 10375 10233 10401
rect 10823 10375 10849 10401
rect 11159 10375 11185 10401
rect 7407 10319 7433 10345
rect 7855 10319 7881 10345
rect 8191 10319 8217 10345
rect 8527 10319 8553 10345
rect 8807 10319 8833 10345
rect 9031 10319 9057 10345
rect 9423 10319 9449 10345
rect 9535 10319 9561 10345
rect 9871 10319 9897 10345
rect 9983 10319 10009 10345
rect 10935 10319 10961 10345
rect 14631 10319 14657 10345
rect 9199 10263 9225 10289
rect 9479 10263 9505 10289
rect 10207 10263 10233 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 9255 10095 9281 10121
rect 13399 10095 13425 10121
rect 7295 10039 7321 10065
rect 8023 10039 8049 10065
rect 8135 10039 8161 10065
rect 11159 10039 11185 10065
rect 12615 10039 12641 10065
rect 12839 10039 12865 10065
rect 7127 9983 7153 10009
rect 7463 9983 7489 10009
rect 7743 9983 7769 10009
rect 8807 9983 8833 10009
rect 9423 9983 9449 10009
rect 12727 9983 12753 10009
rect 12895 9983 12921 10009
rect 13231 9983 13257 10009
rect 13567 9983 13593 10009
rect 18831 9983 18857 10009
rect 6567 9927 6593 9953
rect 8079 9927 8105 9953
rect 9031 9927 9057 9953
rect 13119 9927 13145 9953
rect 13959 9927 13985 9953
rect 15023 9927 15049 9953
rect 12895 9871 12921 9897
rect 20007 9871 20033 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 12111 9703 12137 9729
rect 5391 9647 5417 9673
rect 6455 9647 6481 9673
rect 13791 9647 13817 9673
rect 20007 9647 20033 9673
rect 5055 9591 5081 9617
rect 7407 9591 7433 9617
rect 7519 9591 7545 9617
rect 9143 9591 9169 9617
rect 9759 9591 9785 9617
rect 10039 9591 10065 9617
rect 10095 9591 10121 9617
rect 10991 9591 11017 9617
rect 11495 9591 11521 9617
rect 11719 9591 11745 9617
rect 13175 9591 13201 9617
rect 13511 9591 13537 9617
rect 14183 9591 14209 9617
rect 14239 9591 14265 9617
rect 18943 9591 18969 9617
rect 6735 9535 6761 9561
rect 6903 9535 6929 9561
rect 7071 9535 7097 9561
rect 7911 9535 7937 9561
rect 8079 9535 8105 9561
rect 8303 9535 8329 9561
rect 9255 9535 9281 9561
rect 9311 9535 9337 9561
rect 9983 9535 10009 9561
rect 10935 9535 10961 9561
rect 12671 9535 12697 9561
rect 12839 9535 12865 9561
rect 13735 9535 13761 9561
rect 14015 9535 14041 9561
rect 8359 9479 8385 9505
rect 9479 9479 9505 9505
rect 10319 9479 10345 9505
rect 12503 9479 12529 9505
rect 13007 9479 13033 9505
rect 13343 9479 13369 9505
rect 13623 9479 13649 9505
rect 13791 9479 13817 9505
rect 14071 9479 14097 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 7239 9311 7265 9337
rect 7575 9311 7601 9337
rect 9647 9311 9673 9337
rect 9983 9311 10009 9337
rect 10095 9311 10121 9337
rect 11943 9311 11969 9337
rect 12839 9311 12865 9337
rect 13455 9311 13481 9337
rect 7911 9255 7937 9281
rect 11327 9255 11353 9281
rect 12783 9255 12809 9281
rect 13287 9255 13313 9281
rect 13343 9255 13369 9281
rect 13959 9255 13985 9281
rect 15359 9255 15385 9281
rect 5279 9199 5305 9225
rect 7127 9199 7153 9225
rect 7407 9199 7433 9225
rect 8135 9199 8161 9225
rect 8359 9199 8385 9225
rect 9591 9199 9617 9225
rect 9871 9199 9897 9225
rect 10207 9199 10233 9225
rect 10935 9199 10961 9225
rect 11159 9199 11185 9225
rect 13567 9199 13593 9225
rect 15247 9199 15273 9225
rect 18831 9199 18857 9225
rect 5615 9143 5641 9169
rect 6679 9143 6705 9169
rect 6903 9143 6929 9169
rect 8191 9143 8217 9169
rect 10039 9143 10065 9169
rect 11047 9143 11073 9169
rect 11663 9143 11689 9169
rect 13119 9143 13145 9169
rect 15023 9143 15049 9169
rect 11775 9087 11801 9113
rect 12839 9087 12865 9113
rect 20007 9087 20033 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 7911 8919 7937 8945
rect 9647 8919 9673 8945
rect 10655 8919 10681 8945
rect 10711 8919 10737 8945
rect 10823 8919 10849 8945
rect 10879 8919 10905 8945
rect 11607 8919 11633 8945
rect 9535 8863 9561 8889
rect 11495 8863 11521 8889
rect 13847 8863 13873 8889
rect 20007 8863 20033 8889
rect 9927 8807 9953 8833
rect 10151 8807 10177 8833
rect 11439 8807 11465 8833
rect 12615 8807 12641 8833
rect 12839 8807 12865 8833
rect 12951 8807 12977 8833
rect 13735 8807 13761 8833
rect 13903 8807 13929 8833
rect 14071 8807 14097 8833
rect 18831 8807 18857 8833
rect 9255 8751 9281 8777
rect 9367 8751 9393 8777
rect 9423 8751 9449 8777
rect 9871 8751 9897 8777
rect 7799 8695 7825 8721
rect 7855 8695 7881 8721
rect 8415 8695 8441 8721
rect 12783 8695 12809 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 9031 8527 9057 8553
rect 10319 8527 10345 8553
rect 12223 8527 12249 8553
rect 12335 8527 12361 8553
rect 7239 8471 7265 8497
rect 8863 8471 8889 8497
rect 8919 8471 8945 8497
rect 11383 8471 11409 8497
rect 11495 8471 11521 8497
rect 12111 8471 12137 8497
rect 13007 8471 13033 8497
rect 6903 8415 6929 8441
rect 9535 8415 9561 8441
rect 9759 8415 9785 8441
rect 12671 8415 12697 8441
rect 14295 8415 14321 8441
rect 8303 8359 8329 8385
rect 10207 8359 10233 8385
rect 12391 8359 12417 8385
rect 14071 8359 14097 8385
rect 10375 8303 10401 8329
rect 11551 8303 11577 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 7687 8079 7713 8105
rect 8751 8079 8777 8105
rect 12167 8079 12193 8105
rect 7351 8023 7377 8049
rect 9871 8023 9897 8049
rect 11551 8023 11577 8049
rect 11775 8023 11801 8049
rect 11943 8023 11969 8049
rect 12111 8023 12137 8049
rect 9983 7967 10009 7993
rect 11383 7967 11409 7993
rect 11439 7967 11465 7993
rect 11663 7967 11689 7993
rect 8975 7911 9001 7937
rect 11607 7911 11633 7937
rect 12223 7911 12249 7937
rect 12335 7911 12361 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 9535 7687 9561 7713
rect 9703 7631 9729 7657
rect 9815 7631 9841 7657
rect 10767 7631 10793 7657
rect 9591 7575 9617 7601
rect 10655 7575 10681 7601
rect 9815 7519 9841 7545
rect 10599 7519 10625 7545
rect 10823 7519 10849 7545
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 9759 7351 9785 7377
rect 10207 7351 10233 7377
rect 8527 7295 8553 7321
rect 9591 7295 9617 7321
rect 10711 7295 10737 7321
rect 11887 7295 11913 7321
rect 12951 7295 12977 7321
rect 8191 7239 8217 7265
rect 10375 7239 10401 7265
rect 10767 7239 10793 7265
rect 10935 7239 10961 7265
rect 11495 7239 11521 7265
rect 9815 7183 9841 7209
rect 10655 7183 10681 7209
rect 10039 7127 10065 7153
rect 10263 7127 10289 7153
rect 13175 7127 13201 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 9983 6959 10009 6985
rect 9703 6903 9729 6929
rect 10039 6903 10065 6929
rect 10823 6903 10849 6929
rect 12335 6903 12361 6929
rect 9871 6847 9897 6873
rect 10263 6847 10289 6873
rect 10487 6847 10513 6873
rect 12167 6847 12193 6873
rect 9647 6791 9673 6817
rect 9927 6791 9953 6817
rect 11943 6791 11969 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9311 6511 9337 6537
rect 10375 6511 10401 6537
rect 10711 6511 10737 6537
rect 12167 6511 12193 6537
rect 8975 6455 9001 6481
rect 11607 6455 11633 6481
rect 11719 6343 11745 6369
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 12391 2591 12417 2617
rect 11887 2535 11913 2561
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 8863 2143 8889 2169
rect 10543 2143 10569 2169
rect 12671 2143 12697 2169
rect 9367 2031 9393 2057
rect 11047 2031 11073 2057
rect 13119 2031 13145 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 12783 1807 12809 1833
rect 9871 1751 9897 1777
rect 11775 1751 11801 1777
rect 12279 1751 12305 1777
rect 11103 1695 11129 1721
rect 9591 1639 9617 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 3024 20600 3080 21000
rect 8064 20600 8120 21000
rect 8400 20600 8456 21000
rect 10080 20600 10136 21000
rect 10416 20600 10472 21000
rect 11760 20600 11816 21000
rect 12432 20600 12488 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 3038 18970 3066 20600
rect 3150 18970 3178 18975
rect 3038 18969 3178 18970
rect 3038 18943 3151 18969
rect 3177 18943 3178 18969
rect 3038 18942 3178 18943
rect 3150 18937 3178 18942
rect 8078 18746 8106 20600
rect 8414 19138 8442 20600
rect 8414 19105 8442 19110
rect 9030 19138 9058 19143
rect 9030 19091 9058 19110
rect 8078 18713 8106 18718
rect 8526 19025 8554 19031
rect 8526 18999 8527 19025
rect 8553 18999 8554 19025
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 8526 15974 8554 18999
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 9198 18746 9226 18751
rect 9198 18699 9226 18718
rect 10094 18746 10122 20600
rect 10430 19138 10458 20600
rect 10430 19105 10458 19110
rect 11046 19138 11074 19143
rect 11046 19091 11074 19110
rect 11774 19138 11802 20600
rect 11774 19105 11802 19110
rect 10094 18713 10122 18718
rect 10542 19025 10570 19031
rect 10542 18999 10543 19025
rect 10569 18999 10570 19025
rect 8414 15946 8554 15974
rect 8862 18633 8890 18639
rect 8862 18607 8863 18633
rect 8889 18607 8890 18633
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 8414 14266 8442 15946
rect 8302 14238 8498 14266
rect 8302 14041 8330 14238
rect 8302 14015 8303 14041
rect 8329 14015 8330 14041
rect 8302 14009 8330 14015
rect 8022 13985 8050 13991
rect 8022 13959 8023 13985
rect 8049 13959 8050 13985
rect 8022 13930 8050 13959
rect 7742 13902 8050 13930
rect 8078 13930 8106 13935
rect 8190 13930 8218 13935
rect 8078 13929 8218 13930
rect 8078 13903 8079 13929
rect 8105 13903 8191 13929
rect 8217 13903 8218 13929
rect 8078 13902 8218 13903
rect 7406 13818 7434 13823
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 7406 13593 7434 13790
rect 7406 13567 7407 13593
rect 7433 13567 7434 13593
rect 7406 13561 7434 13567
rect 7070 13537 7098 13543
rect 7070 13511 7071 13537
rect 7097 13511 7098 13537
rect 2086 13482 2114 13487
rect 966 12250 994 12255
rect 966 12203 994 12222
rect 966 11466 994 11471
rect 966 11419 994 11438
rect 966 11242 994 11247
rect 966 11195 994 11214
rect 2086 9954 2114 13454
rect 6958 13146 6986 13151
rect 7070 13146 7098 13511
rect 6958 13145 7098 13146
rect 6958 13119 6959 13145
rect 6985 13119 7098 13145
rect 6958 13118 7098 13119
rect 6958 13113 6986 13118
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 2142 12362 2170 12367
rect 2142 12315 2170 12334
rect 6734 12362 6762 12367
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 6734 12026 6762 12334
rect 6734 11979 6762 11998
rect 6454 11690 6482 11695
rect 5278 11634 5306 11639
rect 2142 11578 2170 11583
rect 2142 11531 2170 11550
rect 5278 11521 5306 11606
rect 5278 11495 5279 11521
rect 5305 11495 5306 11521
rect 5278 11489 5306 11495
rect 6342 11522 6370 11527
rect 6342 11475 6370 11494
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 4998 11241 5026 11247
rect 4998 11215 4999 11241
rect 5025 11215 5026 11241
rect 2142 11186 2170 11191
rect 2142 11139 2170 11158
rect 4998 11130 5026 11215
rect 6454 11186 6482 11662
rect 6734 11690 6762 11695
rect 6734 11577 6762 11662
rect 7070 11690 7098 13118
rect 7294 13090 7322 13095
rect 7294 13043 7322 13062
rect 7742 12698 7770 13902
rect 8078 13897 8106 13902
rect 8190 13897 8218 13902
rect 8358 13929 8386 13935
rect 8358 13903 8359 13929
rect 8385 13903 8386 13929
rect 8022 13818 8050 13823
rect 8022 13771 8050 13790
rect 8358 13314 8386 13903
rect 8470 13593 8498 14238
rect 8806 13874 8834 13879
rect 8470 13567 8471 13593
rect 8497 13567 8498 13593
rect 8470 13561 8498 13567
rect 8694 13846 8806 13874
rect 8694 13538 8722 13846
rect 8806 13827 8834 13846
rect 8862 13762 8890 18607
rect 10206 18633 10234 18639
rect 10206 18607 10207 18633
rect 10233 18607 10234 18633
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 10206 15974 10234 18607
rect 10542 15974 10570 18999
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 10710 18746 10738 18751
rect 10710 18699 10738 18718
rect 12278 15974 12306 18999
rect 12446 18746 12474 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 12446 18713 12474 18718
rect 13118 18746 13146 18751
rect 13118 18699 13146 18718
rect 10094 15946 10234 15974
rect 10486 15946 10570 15974
rect 11886 15946 12306 15974
rect 12614 18633 12642 18639
rect 12614 18607 12615 18633
rect 12641 18607 12642 18633
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9086 13929 9114 13935
rect 9086 13903 9087 13929
rect 9113 13903 9114 13929
rect 9086 13874 9114 13903
rect 9086 13841 9114 13846
rect 9422 13873 9450 13879
rect 9422 13847 9423 13873
rect 9449 13847 9450 13873
rect 8358 13281 8386 13286
rect 8526 13537 8722 13538
rect 8526 13511 8695 13537
rect 8721 13511 8722 13537
rect 8526 13510 8722 13511
rect 8358 13202 8386 13207
rect 7910 13090 7938 13095
rect 7910 12753 7938 13062
rect 8358 13089 8386 13174
rect 8358 13063 8359 13089
rect 8385 13063 8386 13089
rect 8358 13057 8386 13063
rect 7910 12727 7911 12753
rect 7937 12727 7938 12753
rect 7910 12721 7938 12727
rect 8078 13034 8106 13039
rect 8078 12753 8106 13006
rect 8078 12727 8079 12753
rect 8105 12727 8106 12753
rect 8078 12721 8106 12727
rect 7070 11657 7098 11662
rect 7406 11914 7434 11919
rect 7406 11689 7434 11886
rect 7574 11690 7602 11695
rect 7630 11690 7658 11695
rect 7406 11663 7407 11689
rect 7433 11663 7434 11689
rect 7406 11657 7434 11663
rect 7518 11662 7574 11690
rect 7602 11689 7658 11690
rect 7602 11663 7631 11689
rect 7657 11663 7658 11689
rect 7602 11662 7658 11663
rect 6958 11634 6986 11639
rect 6958 11587 6986 11606
rect 6734 11551 6735 11577
rect 6761 11551 6762 11577
rect 6734 11545 6762 11551
rect 7014 11578 7042 11583
rect 7014 11531 7042 11550
rect 7294 11578 7322 11583
rect 6790 11522 6818 11527
rect 6790 11241 6818 11494
rect 6790 11215 6791 11241
rect 6817 11215 6818 11241
rect 6790 11209 6818 11215
rect 6958 11465 6986 11471
rect 6958 11439 6959 11465
rect 6985 11439 6986 11465
rect 6454 11185 6538 11186
rect 6454 11159 6455 11185
rect 6481 11159 6538 11185
rect 6454 11158 6538 11159
rect 6454 11153 6482 11158
rect 4998 11097 5026 11102
rect 6062 11130 6090 11135
rect 6062 11129 6426 11130
rect 6062 11103 6063 11129
rect 6089 11103 6426 11129
rect 6062 11102 6426 11103
rect 6062 11097 6090 11102
rect 6398 10905 6426 11102
rect 6398 10879 6399 10905
rect 6425 10879 6426 10905
rect 6398 10873 6426 10879
rect 5390 10794 5418 10799
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 2086 9921 2114 9926
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 5390 9673 5418 10766
rect 6454 10682 6482 10687
rect 6454 10635 6482 10654
rect 6510 10094 6538 11158
rect 6958 11129 6986 11439
rect 7294 11185 7322 11550
rect 7350 11522 7378 11527
rect 7350 11475 7378 11494
rect 7518 11241 7546 11662
rect 7574 11657 7602 11662
rect 7630 11657 7658 11662
rect 7518 11215 7519 11241
rect 7545 11215 7546 11241
rect 7518 11209 7546 11215
rect 7686 11466 7714 11471
rect 7294 11159 7295 11185
rect 7321 11159 7322 11185
rect 7294 11153 7322 11159
rect 7686 11185 7714 11438
rect 7686 11159 7687 11185
rect 7713 11159 7714 11185
rect 7686 11153 7714 11159
rect 6958 11103 6959 11129
rect 6985 11103 6986 11129
rect 6958 11097 6986 11103
rect 7238 11130 7266 11135
rect 7238 11083 7266 11102
rect 6734 11073 6762 11079
rect 6846 11074 6874 11079
rect 7126 11074 7154 11079
rect 7742 11074 7770 12670
rect 8022 12641 8050 12647
rect 8022 12615 8023 12641
rect 8049 12615 8050 12641
rect 7966 12026 7994 12031
rect 7798 11914 7826 11919
rect 7798 11867 7826 11886
rect 7854 11802 7882 11807
rect 7854 11241 7882 11774
rect 7966 11689 7994 11998
rect 8022 11802 8050 12615
rect 8470 12642 8498 12647
rect 8526 12642 8554 13510
rect 8694 13505 8722 13510
rect 8750 13734 8890 13762
rect 8750 13202 8778 13734
rect 9422 13650 9450 13847
rect 9422 13617 9450 13622
rect 10094 13594 10122 15946
rect 10486 13873 10514 15946
rect 10486 13847 10487 13873
rect 10513 13847 10514 13873
rect 10318 13650 10346 13655
rect 10318 13603 10346 13622
rect 10094 13593 10234 13594
rect 10094 13567 10095 13593
rect 10121 13567 10234 13593
rect 10094 13566 10234 13567
rect 10094 13561 10122 13566
rect 9030 13481 9058 13487
rect 9030 13455 9031 13481
rect 9057 13455 9058 13481
rect 8750 13155 8778 13174
rect 8806 13314 8834 13319
rect 8806 13201 8834 13286
rect 9030 13258 9058 13455
rect 10094 13482 10122 13487
rect 9918 13342 10050 13347
rect 9030 13225 9058 13230
rect 9254 13314 9282 13319
rect 8806 13175 8807 13201
rect 8833 13175 8834 13201
rect 8806 13169 8834 13175
rect 8750 13034 8778 13039
rect 8750 12987 8778 13006
rect 9254 12697 9282 13286
rect 9814 13314 9842 13319
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9534 13258 9562 13263
rect 9534 13211 9562 13230
rect 9254 12671 9255 12697
rect 9281 12671 9282 12697
rect 9254 12665 9282 12671
rect 9646 13201 9674 13207
rect 9646 13175 9647 13201
rect 9673 13175 9674 13201
rect 8470 12641 8554 12642
rect 8470 12615 8471 12641
rect 8497 12615 8554 12641
rect 8470 12614 8554 12615
rect 8470 12609 8498 12614
rect 8022 11769 8050 11774
rect 8134 11969 8162 11975
rect 8134 11943 8135 11969
rect 8161 11943 8162 11969
rect 8134 11858 8162 11943
rect 8470 11913 8498 11919
rect 8470 11887 8471 11913
rect 8497 11887 8498 11913
rect 7966 11663 7967 11689
rect 7993 11663 7994 11689
rect 7966 11657 7994 11663
rect 8134 11690 8162 11830
rect 8302 11858 8330 11863
rect 8302 11857 8386 11858
rect 8302 11831 8303 11857
rect 8329 11831 8386 11857
rect 8302 11830 8386 11831
rect 8302 11825 8330 11830
rect 7910 11634 7938 11639
rect 7910 11587 7938 11606
rect 8078 11577 8106 11583
rect 8078 11551 8079 11577
rect 8105 11551 8106 11577
rect 8022 11522 8050 11527
rect 8022 11475 8050 11494
rect 8078 11466 8106 11551
rect 8078 11433 8106 11438
rect 7854 11215 7855 11241
rect 7881 11215 7882 11241
rect 7854 11209 7882 11215
rect 8134 11185 8162 11662
rect 8134 11159 8135 11185
rect 8161 11159 8162 11185
rect 8134 11153 8162 11159
rect 8190 11578 8218 11583
rect 6734 11047 6735 11073
rect 6761 11047 6762 11073
rect 6566 10906 6594 10911
rect 6734 10906 6762 11047
rect 6566 10793 6594 10878
rect 6566 10767 6567 10793
rect 6593 10767 6594 10793
rect 6566 10761 6594 10767
rect 6678 10878 6762 10906
rect 6790 11073 6874 11074
rect 6790 11047 6847 11073
rect 6873 11047 6874 11073
rect 6790 11046 6874 11047
rect 6678 10682 6706 10878
rect 6790 10850 6818 11046
rect 6846 11041 6874 11046
rect 7014 11073 7154 11074
rect 7014 11047 7127 11073
rect 7153 11047 7154 11073
rect 7014 11046 7154 11047
rect 7014 10906 7042 11046
rect 7126 11041 7154 11046
rect 7686 11046 7770 11074
rect 7798 11073 7826 11079
rect 7798 11047 7799 11073
rect 7825 11047 7826 11073
rect 6790 10817 6818 10822
rect 6846 10878 7042 10906
rect 7238 10906 7266 10911
rect 6846 10849 6874 10878
rect 6846 10823 6847 10849
rect 6873 10823 6874 10849
rect 6846 10817 6874 10823
rect 7126 10850 7154 10855
rect 6734 10794 6762 10799
rect 6734 10747 6762 10766
rect 7070 10794 7098 10799
rect 7126 10794 7154 10822
rect 7070 10793 7154 10794
rect 7070 10767 7071 10793
rect 7097 10767 7154 10793
rect 7070 10766 7154 10767
rect 7182 10849 7210 10855
rect 7182 10823 7183 10849
rect 7209 10823 7210 10849
rect 7182 10794 7210 10823
rect 7238 10849 7266 10878
rect 7238 10823 7239 10849
rect 7265 10823 7266 10849
rect 7238 10817 7266 10823
rect 7406 10906 7434 10911
rect 7070 10761 7098 10766
rect 7182 10761 7210 10766
rect 6734 10682 6762 10687
rect 6678 10654 6734 10682
rect 6734 10649 6762 10654
rect 7406 10345 7434 10878
rect 7686 10905 7714 11046
rect 7686 10879 7687 10905
rect 7713 10879 7714 10905
rect 7686 10873 7714 10879
rect 7798 10906 7826 11047
rect 7910 11073 7938 11079
rect 7910 11047 7911 11073
rect 7937 11047 7938 11073
rect 7854 10906 7882 10911
rect 7798 10878 7854 10906
rect 7854 10859 7882 10878
rect 7742 10850 7770 10855
rect 7742 10849 7826 10850
rect 7742 10823 7743 10849
rect 7769 10823 7826 10849
rect 7742 10822 7826 10823
rect 7742 10817 7770 10822
rect 7798 10794 7826 10822
rect 7798 10513 7826 10766
rect 7798 10487 7799 10513
rect 7825 10487 7826 10513
rect 7798 10481 7826 10487
rect 7574 10458 7602 10463
rect 7406 10319 7407 10345
rect 7433 10319 7434 10345
rect 7406 10313 7434 10319
rect 7518 10401 7546 10407
rect 7518 10375 7519 10401
rect 7545 10375 7546 10401
rect 6510 10066 6594 10094
rect 5390 9647 5391 9673
rect 5417 9647 5418 9673
rect 5390 9641 5418 9647
rect 6454 10010 6482 10015
rect 6454 9673 6482 9982
rect 6454 9647 6455 9673
rect 6481 9647 6482 9673
rect 6454 9641 6482 9647
rect 6566 9953 6594 10066
rect 7294 10065 7322 10071
rect 7294 10039 7295 10065
rect 7321 10039 7322 10065
rect 7126 10010 7154 10015
rect 7126 9963 7154 9982
rect 6566 9927 6567 9953
rect 6593 9927 6594 9953
rect 5054 9617 5082 9623
rect 5054 9591 5055 9617
rect 5081 9591 5082 9617
rect 5054 9282 5082 9591
rect 5054 9249 5082 9254
rect 5278 9282 5306 9287
rect 5278 9225 5306 9254
rect 6566 9282 6594 9927
rect 6566 9249 6594 9254
rect 6734 9730 6762 9735
rect 6734 9561 6762 9702
rect 7294 9618 7322 10039
rect 7462 10010 7490 10015
rect 7462 9963 7490 9982
rect 7406 9618 7434 9623
rect 7294 9590 7406 9618
rect 7406 9571 7434 9590
rect 7518 9617 7546 10375
rect 7518 9591 7519 9617
rect 7545 9591 7546 9617
rect 6734 9535 6735 9561
rect 6761 9535 6762 9561
rect 5278 9199 5279 9225
rect 5305 9199 5306 9225
rect 5278 9193 5306 9199
rect 6678 9226 6706 9231
rect 5614 9170 5642 9175
rect 5614 9123 5642 9142
rect 6678 9169 6706 9198
rect 6678 9143 6679 9169
rect 6705 9143 6706 9169
rect 6678 9137 6706 9143
rect 6734 9170 6762 9535
rect 6902 9562 6930 9567
rect 7070 9562 7098 9567
rect 6902 9561 7098 9562
rect 6902 9535 6903 9561
rect 6929 9535 7071 9561
rect 7097 9535 7098 9561
rect 6902 9534 7098 9535
rect 6902 9529 6930 9534
rect 7070 9529 7098 9534
rect 7238 9562 7266 9567
rect 7238 9337 7266 9534
rect 7518 9562 7546 9591
rect 7518 9529 7546 9534
rect 7238 9311 7239 9337
rect 7265 9311 7266 9337
rect 7238 9305 7266 9311
rect 7574 9337 7602 10430
rect 7742 10346 7770 10351
rect 7742 10009 7770 10318
rect 7742 9983 7743 10009
rect 7769 9983 7770 10009
rect 7742 9977 7770 9983
rect 7854 10345 7882 10351
rect 7854 10319 7855 10345
rect 7881 10319 7882 10345
rect 7854 9618 7882 10319
rect 7910 9786 7938 11047
rect 8022 10794 8050 10799
rect 8022 10065 8050 10766
rect 8190 10457 8218 11550
rect 8358 11242 8386 11830
rect 8414 11857 8442 11863
rect 8414 11831 8415 11857
rect 8441 11831 8442 11857
rect 8414 11802 8442 11831
rect 8414 11769 8442 11774
rect 8470 11354 8498 11887
rect 8526 11858 8554 12614
rect 9422 12641 9450 12647
rect 9422 12615 9423 12641
rect 9449 12615 9450 12641
rect 9422 12306 9450 12615
rect 9366 12082 9394 12087
rect 9310 12054 9366 12082
rect 8526 11825 8554 11830
rect 8694 11858 8722 11863
rect 8694 11811 8722 11830
rect 9086 11690 9114 11695
rect 9086 11643 9114 11662
rect 8918 11634 8946 11639
rect 8470 11326 8722 11354
rect 8470 11242 8498 11247
rect 8358 11241 8498 11242
rect 8358 11215 8471 11241
rect 8497 11215 8498 11241
rect 8358 11214 8498 11215
rect 8470 11209 8498 11214
rect 8190 10431 8191 10457
rect 8217 10431 8218 10457
rect 8190 10425 8218 10431
rect 8470 10458 8498 10463
rect 8022 10039 8023 10065
rect 8049 10039 8050 10065
rect 8022 10033 8050 10039
rect 8134 10402 8162 10407
rect 8134 10065 8162 10374
rect 8302 10402 8330 10407
rect 8470 10402 8498 10430
rect 8302 10401 8498 10402
rect 8302 10375 8303 10401
rect 8329 10375 8471 10401
rect 8497 10375 8498 10401
rect 8302 10374 8498 10375
rect 8302 10369 8330 10374
rect 8470 10369 8498 10374
rect 8638 10402 8666 10407
rect 8638 10355 8666 10374
rect 8694 10401 8722 11326
rect 8694 10375 8695 10401
rect 8721 10375 8722 10401
rect 8694 10369 8722 10375
rect 8806 10906 8834 10911
rect 8190 10346 8218 10351
rect 8190 10299 8218 10318
rect 8526 10346 8554 10351
rect 8526 10299 8554 10318
rect 8806 10345 8834 10878
rect 8862 10402 8890 10407
rect 8862 10355 8890 10374
rect 8806 10319 8807 10345
rect 8833 10319 8834 10345
rect 8806 10313 8834 10319
rect 8918 10290 8946 11606
rect 9142 11074 9170 11079
rect 9030 10794 9058 10799
rect 8134 10039 8135 10065
rect 8161 10039 8162 10065
rect 8134 10033 8162 10039
rect 8862 10262 8946 10290
rect 8974 10682 9002 10687
rect 8806 10010 8834 10015
rect 8806 9963 8834 9982
rect 8078 9954 8106 9959
rect 7910 9753 7938 9758
rect 8022 9953 8106 9954
rect 8022 9927 8079 9953
rect 8105 9927 8106 9953
rect 8022 9926 8106 9927
rect 8022 9730 8050 9926
rect 8078 9921 8106 9926
rect 7966 9702 8050 9730
rect 8078 9786 8106 9791
rect 7910 9618 7938 9623
rect 7854 9590 7910 9618
rect 7574 9311 7575 9337
rect 7601 9311 7602 9337
rect 7574 9305 7602 9311
rect 7910 9561 7938 9590
rect 7910 9535 7911 9561
rect 7937 9535 7938 9561
rect 6734 9137 6762 9142
rect 6902 9282 6930 9287
rect 6902 9169 6930 9254
rect 7910 9281 7938 9535
rect 7910 9255 7911 9281
rect 7937 9255 7938 9281
rect 7910 9249 7938 9255
rect 7126 9226 7154 9231
rect 7126 9179 7154 9198
rect 7406 9226 7434 9231
rect 7406 9179 7434 9198
rect 6902 9143 6903 9169
rect 6929 9143 6930 9169
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 6902 8442 6930 9143
rect 7910 8946 7938 8951
rect 7966 8946 7994 9702
rect 8078 9561 8106 9758
rect 8190 9562 8218 9567
rect 8302 9562 8330 9567
rect 8078 9535 8079 9561
rect 8105 9535 8106 9561
rect 8078 9529 8106 9535
rect 8134 9534 8190 9562
rect 8218 9561 8330 9562
rect 8218 9535 8303 9561
rect 8329 9535 8330 9561
rect 8218 9534 8330 9535
rect 8134 9225 8162 9534
rect 8190 9515 8218 9534
rect 8302 9529 8330 9534
rect 8358 9506 8386 9511
rect 8358 9459 8386 9478
rect 8134 9199 8135 9225
rect 8161 9199 8162 9225
rect 8134 9193 8162 9199
rect 8358 9225 8386 9231
rect 8358 9199 8359 9225
rect 8385 9199 8386 9225
rect 7910 8945 7994 8946
rect 7910 8919 7911 8945
rect 7937 8919 7994 8945
rect 7910 8918 7994 8919
rect 8190 9169 8218 9175
rect 8190 9143 8191 9169
rect 8217 9143 8218 9169
rect 7910 8913 7938 8918
rect 7238 8722 7266 8727
rect 7238 8497 7266 8694
rect 7798 8721 7826 8727
rect 7798 8695 7799 8721
rect 7825 8695 7826 8721
rect 7798 8554 7826 8695
rect 7854 8722 7882 8727
rect 7854 8675 7882 8694
rect 7798 8521 7826 8526
rect 8190 8554 8218 9143
rect 8190 8521 8218 8526
rect 7238 8471 7239 8497
rect 7265 8471 7266 8497
rect 7238 8465 7266 8471
rect 7686 8498 7714 8503
rect 6902 8395 6930 8414
rect 7350 8442 7378 8447
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 7350 8049 7378 8414
rect 7686 8105 7714 8470
rect 8302 8386 8330 8391
rect 8358 8386 8386 9199
rect 8302 8385 8358 8386
rect 8302 8359 8303 8385
rect 8329 8359 8358 8385
rect 8302 8358 8358 8359
rect 8302 8353 8330 8358
rect 8358 8353 8386 8358
rect 8414 8721 8442 8727
rect 8414 8695 8415 8721
rect 8441 8695 8442 8721
rect 8414 8442 8442 8695
rect 8862 8497 8890 10262
rect 8974 9842 9002 10654
rect 9030 10345 9058 10766
rect 9030 10319 9031 10345
rect 9057 10319 9058 10345
rect 9030 10313 9058 10319
rect 9142 10122 9170 11046
rect 9198 10290 9226 10295
rect 9198 10243 9226 10262
rect 9254 10122 9282 10127
rect 9142 10121 9282 10122
rect 9142 10095 9255 10121
rect 9281 10095 9282 10121
rect 9142 10094 9282 10095
rect 9254 10089 9282 10094
rect 9310 10066 9338 12054
rect 9366 12049 9394 12054
rect 9366 11858 9394 11863
rect 9366 11521 9394 11830
rect 9366 11495 9367 11521
rect 9393 11495 9394 11521
rect 9366 10849 9394 11495
rect 9422 11690 9450 12278
rect 9646 11690 9674 13175
rect 9814 13202 9842 13286
rect 9926 13258 9954 13263
rect 9926 13211 9954 13230
rect 10038 13258 10066 13263
rect 10094 13258 10122 13454
rect 10038 13257 10122 13258
rect 10038 13231 10039 13257
rect 10065 13231 10122 13257
rect 10038 13230 10122 13231
rect 10206 13257 10234 13566
rect 10262 13482 10290 13487
rect 10262 13435 10290 13454
rect 10318 13426 10346 13431
rect 10318 13425 10458 13426
rect 10318 13399 10319 13425
rect 10345 13399 10458 13425
rect 10318 13398 10458 13399
rect 10318 13393 10346 13398
rect 10206 13231 10207 13257
rect 10233 13231 10234 13257
rect 10038 13225 10066 13230
rect 10206 13225 10234 13231
rect 9870 13202 9898 13207
rect 9814 13174 9870 13202
rect 9870 13155 9898 13174
rect 10150 13202 10178 13207
rect 10150 13155 10178 13174
rect 9702 13146 9730 13151
rect 9702 13099 9730 13118
rect 10318 13146 10346 13151
rect 10318 13099 10346 13118
rect 10430 12810 10458 13398
rect 10486 13258 10514 13847
rect 10710 13874 10738 13879
rect 10710 13593 10738 13846
rect 10710 13567 10711 13593
rect 10737 13567 10738 13593
rect 10710 13561 10738 13567
rect 10486 13225 10514 13230
rect 11046 13537 11074 13543
rect 11046 13511 11047 13537
rect 11073 13511 11074 13537
rect 10430 12782 10794 12810
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9814 12082 9842 12087
rect 9814 12035 9842 12054
rect 10430 12081 10458 12782
rect 10766 12753 10794 12782
rect 10766 12727 10767 12753
rect 10793 12727 10794 12753
rect 10766 12721 10794 12727
rect 10878 12698 10906 12703
rect 10878 12651 10906 12670
rect 10934 12698 10962 12703
rect 10934 12697 11018 12698
rect 10934 12671 10935 12697
rect 10961 12671 11018 12697
rect 10934 12670 11018 12671
rect 10934 12665 10962 12670
rect 10598 12586 10626 12591
rect 10598 12361 10626 12558
rect 10598 12335 10599 12361
rect 10625 12335 10626 12361
rect 10598 12329 10626 12335
rect 10934 12305 10962 12311
rect 10934 12279 10935 12305
rect 10961 12279 10962 12305
rect 10430 12055 10431 12081
rect 10457 12055 10458 12081
rect 9758 11913 9786 11919
rect 9758 11887 9759 11913
rect 9785 11887 9786 11913
rect 9702 11690 9730 11695
rect 9646 11662 9702 11690
rect 9422 11522 9450 11662
rect 9702 11643 9730 11662
rect 9590 11633 9618 11639
rect 9590 11607 9591 11633
rect 9617 11607 9618 11633
rect 9422 11489 9450 11494
rect 9534 11577 9562 11583
rect 9534 11551 9535 11577
rect 9561 11551 9562 11577
rect 9534 11410 9562 11551
rect 9590 11578 9618 11607
rect 9590 11545 9618 11550
rect 9758 11410 9786 11887
rect 10150 11914 10178 11919
rect 10430 11914 10458 12055
rect 10766 12082 10794 12087
rect 10934 12082 10962 12279
rect 10766 12081 10962 12082
rect 10766 12055 10767 12081
rect 10793 12055 10962 12081
rect 10766 12054 10962 12055
rect 10766 12049 10794 12054
rect 10710 11970 10738 11975
rect 10150 11913 10234 11914
rect 10150 11887 10151 11913
rect 10177 11887 10234 11913
rect 10150 11886 10234 11887
rect 10150 11881 10178 11886
rect 9814 11857 9842 11863
rect 9814 11831 9815 11857
rect 9841 11831 9842 11857
rect 9814 11690 9842 11831
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9814 11657 9842 11662
rect 9982 11633 10010 11639
rect 9982 11607 9983 11633
rect 10009 11607 10010 11633
rect 9534 11382 9618 11410
rect 9534 11298 9562 11303
rect 9534 11242 9562 11270
rect 9366 10823 9367 10849
rect 9393 10823 9394 10849
rect 9366 10817 9394 10823
rect 9422 11241 9562 11242
rect 9422 11215 9535 11241
rect 9561 11215 9562 11241
rect 9422 11214 9562 11215
rect 9422 10345 9450 11214
rect 9534 11209 9562 11214
rect 9590 10458 9618 11382
rect 9758 11377 9786 11382
rect 9814 11577 9842 11583
rect 9814 11551 9815 11577
rect 9841 11551 9842 11577
rect 9814 11298 9842 11551
rect 9982 11578 10010 11607
rect 10206 11634 10234 11886
rect 10430 11881 10458 11886
rect 10486 11969 10738 11970
rect 10486 11943 10711 11969
rect 10737 11943 10738 11969
rect 10486 11942 10738 11943
rect 10262 11857 10290 11863
rect 10262 11831 10263 11857
rect 10289 11831 10290 11857
rect 10262 11634 10290 11831
rect 10374 11857 10402 11863
rect 10374 11831 10375 11857
rect 10401 11831 10402 11857
rect 10318 11634 10346 11639
rect 10262 11606 10318 11634
rect 10206 11601 10234 11606
rect 10318 11587 10346 11606
rect 10150 11578 10178 11583
rect 9814 11265 9842 11270
rect 9870 11522 9898 11527
rect 9422 10319 9423 10345
rect 9449 10319 9450 10345
rect 9422 10313 9450 10319
rect 9478 10430 9618 10458
rect 9646 11130 9674 11135
rect 9646 10514 9674 11102
rect 9814 11074 9842 11079
rect 9814 11027 9842 11046
rect 9870 11073 9898 11494
rect 9982 11242 10010 11550
rect 9982 11209 10010 11214
rect 10038 11577 10178 11578
rect 10038 11551 10151 11577
rect 10177 11551 10178 11577
rect 10038 11550 10178 11551
rect 9926 11130 9954 11135
rect 10038 11130 10066 11550
rect 10150 11545 10178 11550
rect 10374 11578 10402 11831
rect 10374 11545 10402 11550
rect 10486 11466 10514 11942
rect 10710 11937 10738 11942
rect 10934 11970 10962 11975
rect 10934 11923 10962 11942
rect 10822 11858 10850 11863
rect 10822 11811 10850 11830
rect 10990 11858 11018 12670
rect 11046 12586 11074 13511
rect 11438 13481 11466 13487
rect 11438 13455 11439 13481
rect 11465 13455 11466 13481
rect 11438 13258 11466 13455
rect 11886 13454 11914 15946
rect 11438 13225 11466 13230
rect 11830 13426 11914 13454
rect 11942 13594 11970 13599
rect 11774 13033 11802 13039
rect 11774 13007 11775 13033
rect 11801 13007 11802 13033
rect 11158 12698 11186 12703
rect 11158 12651 11186 12670
rect 11046 12553 11074 12558
rect 11214 12642 11242 12647
rect 11046 11914 11074 11919
rect 11046 11867 11074 11886
rect 10990 11825 11018 11830
rect 10934 11690 10962 11695
rect 10878 11633 10906 11639
rect 10878 11607 10879 11633
rect 10905 11607 10906 11633
rect 10766 11578 10794 11583
rect 10766 11531 10794 11550
rect 10878 11578 10906 11607
rect 10878 11545 10906 11550
rect 10206 11438 10514 11466
rect 9954 11102 10066 11130
rect 10094 11410 10122 11415
rect 10094 11185 10122 11382
rect 10094 11159 10095 11185
rect 10121 11159 10122 11185
rect 9926 11083 9954 11102
rect 9870 11047 9871 11073
rect 9897 11047 9898 11073
rect 9870 11041 9898 11047
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 10094 10794 10122 11159
rect 10094 10761 10122 10766
rect 10150 11242 10178 11247
rect 10150 10682 10178 11214
rect 10206 11073 10234 11438
rect 10654 11298 10682 11303
rect 10654 11185 10682 11270
rect 10654 11159 10655 11185
rect 10681 11159 10682 11185
rect 10654 11153 10682 11159
rect 10206 11047 10207 11073
rect 10233 11047 10234 11073
rect 10206 11041 10234 11047
rect 10262 11129 10290 11135
rect 10262 11103 10263 11129
rect 10289 11103 10290 11129
rect 9478 10290 9506 10430
rect 9478 10243 9506 10262
rect 9534 10345 9562 10351
rect 9534 10319 9535 10345
rect 9561 10319 9562 10345
rect 9310 10033 9338 10038
rect 9422 10010 9450 10015
rect 9422 9963 9450 9982
rect 9030 9954 9058 9959
rect 9030 9953 9226 9954
rect 9030 9927 9031 9953
rect 9057 9927 9226 9953
rect 9030 9926 9226 9927
rect 9030 9921 9058 9926
rect 8974 9814 9170 9842
rect 9142 9617 9170 9814
rect 9142 9591 9143 9617
rect 9169 9591 9170 9617
rect 9142 9170 9170 9591
rect 9198 9562 9226 9926
rect 9254 9562 9282 9567
rect 9198 9534 9254 9562
rect 9254 9515 9282 9534
rect 9310 9561 9338 9567
rect 9310 9535 9311 9561
rect 9337 9535 9338 9561
rect 9142 9137 9170 9142
rect 9254 8778 9282 8783
rect 9030 8777 9282 8778
rect 9030 8751 9255 8777
rect 9281 8751 9282 8777
rect 9030 8750 9282 8751
rect 9030 8553 9058 8750
rect 9254 8745 9282 8750
rect 9030 8527 9031 8553
rect 9057 8527 9058 8553
rect 9030 8521 9058 8527
rect 8862 8471 8863 8497
rect 8889 8471 8890 8497
rect 8862 8465 8890 8471
rect 8918 8497 8946 8503
rect 8918 8471 8919 8497
rect 8945 8471 8946 8497
rect 7686 8079 7687 8105
rect 7713 8079 7714 8105
rect 7686 8073 7714 8079
rect 7350 8023 7351 8049
rect 7377 8023 7378 8049
rect 7350 8017 7378 8023
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 8190 7266 8218 7271
rect 8190 7219 8218 7238
rect 8414 7266 8442 8414
rect 8750 8106 8778 8111
rect 8918 8106 8946 8471
rect 8750 8105 8946 8106
rect 8750 8079 8751 8105
rect 8777 8079 8946 8105
rect 8750 8078 8946 8079
rect 8526 7602 8554 7607
rect 8526 7321 8554 7574
rect 8526 7295 8527 7321
rect 8553 7295 8554 7321
rect 8526 7289 8554 7295
rect 8414 7233 8442 7238
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 8750 4214 8778 8078
rect 9310 7994 9338 9535
rect 9478 9506 9506 9511
rect 9478 9114 9506 9478
rect 9534 9226 9562 10319
rect 9646 9337 9674 10486
rect 9870 10654 10178 10682
rect 9870 10345 9898 10654
rect 9870 10319 9871 10345
rect 9897 10319 9898 10345
rect 9870 10313 9898 10319
rect 9926 10570 9954 10575
rect 9926 10346 9954 10542
rect 9982 10346 10010 10351
rect 9926 10345 10010 10346
rect 9926 10319 9983 10345
rect 10009 10319 10010 10345
rect 9926 10318 10010 10319
rect 9982 10313 10010 10318
rect 10094 10290 10122 10295
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9814 10122 9842 10127
rect 9758 9618 9786 9623
rect 9758 9571 9786 9590
rect 9646 9311 9647 9337
rect 9673 9311 9674 9337
rect 9646 9305 9674 9311
rect 9814 9338 9842 10094
rect 9870 9786 9898 9791
rect 9870 9562 9898 9758
rect 10038 9618 10066 9623
rect 10038 9571 10066 9590
rect 10094 9617 10122 10262
rect 10094 9591 10095 9617
rect 10121 9591 10122 9617
rect 10094 9585 10122 9591
rect 9982 9562 10010 9567
rect 9870 9561 10010 9562
rect 9870 9535 9983 9561
rect 10009 9535 10010 9561
rect 9870 9534 10010 9535
rect 9982 9506 10010 9534
rect 9982 9478 10122 9506
rect 10094 9450 10122 9478
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9982 9338 10010 9343
rect 9814 9337 10010 9338
rect 9814 9311 9983 9337
rect 10009 9311 10010 9337
rect 9814 9310 10010 9311
rect 9982 9305 10010 9310
rect 10094 9337 10122 9422
rect 10094 9311 10095 9337
rect 10121 9311 10122 9337
rect 10094 9305 10122 9311
rect 9534 9193 9562 9198
rect 9590 9225 9618 9231
rect 9590 9199 9591 9225
rect 9617 9199 9618 9225
rect 9534 9114 9562 9119
rect 9478 9086 9534 9114
rect 9534 9081 9562 9086
rect 9534 8890 9562 8895
rect 9534 8843 9562 8862
rect 9366 8778 9394 8783
rect 9366 8731 9394 8750
rect 9422 8777 9450 8783
rect 9422 8751 9423 8777
rect 9449 8751 9450 8777
rect 9422 8498 9450 8751
rect 9422 8465 9450 8470
rect 9534 8442 9562 8447
rect 9590 8442 9618 9199
rect 9870 9225 9898 9231
rect 9870 9199 9871 9225
rect 9897 9199 9898 9225
rect 9870 9170 9898 9199
rect 9870 9137 9898 9142
rect 9926 9226 9954 9231
rect 9646 8946 9674 8951
rect 9646 8899 9674 8918
rect 9926 8890 9954 9198
rect 10038 9169 10066 9175
rect 10038 9143 10039 9169
rect 10065 9143 10066 9169
rect 10038 8946 10066 9143
rect 10038 8913 10066 8918
rect 9534 8441 9618 8442
rect 9534 8415 9535 8441
rect 9561 8415 9618 8441
rect 9534 8414 9618 8415
rect 9758 8862 9954 8890
rect 9758 8441 9786 8862
rect 9926 8833 9954 8862
rect 9926 8807 9927 8833
rect 9953 8807 9954 8833
rect 9926 8801 9954 8807
rect 10150 8833 10178 10654
rect 10206 10514 10234 10519
rect 10206 10401 10234 10486
rect 10206 10375 10207 10401
rect 10233 10375 10234 10401
rect 10206 10369 10234 10375
rect 10206 10289 10234 10295
rect 10206 10263 10207 10289
rect 10233 10263 10234 10289
rect 10206 10122 10234 10263
rect 10206 10089 10234 10094
rect 10262 9730 10290 11103
rect 10374 11130 10402 11135
rect 10374 11129 10626 11130
rect 10374 11103 10375 11129
rect 10401 11103 10626 11129
rect 10374 11102 10626 11103
rect 10374 11097 10402 11102
rect 10262 9697 10290 9702
rect 10598 9674 10626 11102
rect 10934 11129 10962 11662
rect 11214 11690 11242 12614
rect 11774 12642 11802 13007
rect 11774 12609 11802 12614
rect 11830 12306 11858 13426
rect 11886 13258 11914 13263
rect 11942 13258 11970 13566
rect 12502 13594 12530 13599
rect 12614 13594 12642 18607
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 20118 18186 20146 18191
rect 20118 18139 20146 18158
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 12530 13566 12642 13594
rect 20006 13593 20034 13599
rect 20006 13567 20007 13593
rect 20033 13567 20034 13593
rect 12502 13547 12530 13566
rect 13902 13538 13930 13543
rect 13902 13491 13930 13510
rect 14350 13538 14378 13543
rect 12558 13482 12586 13487
rect 11886 13257 11970 13258
rect 11886 13231 11887 13257
rect 11913 13231 11970 13257
rect 11886 13230 11970 13231
rect 12166 13258 12194 13263
rect 11886 13225 11914 13230
rect 12166 13211 12194 13230
rect 12278 13146 12306 13151
rect 12278 13145 12474 13146
rect 12278 13119 12279 13145
rect 12305 13119 12474 13145
rect 12278 13118 12474 13119
rect 12278 13113 12306 13118
rect 11942 13034 11970 13039
rect 12110 13034 12138 13039
rect 11942 13033 12138 13034
rect 11942 13007 11943 13033
rect 11969 13007 12111 13033
rect 12137 13007 12138 13033
rect 11942 13006 12138 13007
rect 11942 13001 11970 13006
rect 12110 13001 12138 13006
rect 12446 12753 12474 13118
rect 12446 12727 12447 12753
rect 12473 12727 12474 12753
rect 12334 12698 12362 12703
rect 12334 12651 12362 12670
rect 12222 12586 12250 12591
rect 12222 12473 12250 12558
rect 12222 12447 12223 12473
rect 12249 12447 12250 12473
rect 12222 12441 12250 12447
rect 12446 12474 12474 12727
rect 12558 12753 12586 13454
rect 13846 13482 13874 13487
rect 13846 13435 13874 13454
rect 12726 13425 12754 13431
rect 12726 13399 12727 13425
rect 12753 13399 12754 13425
rect 12726 13146 12754 13399
rect 12894 13146 12922 13151
rect 12726 13118 12894 13146
rect 12614 13090 12642 13095
rect 12614 12809 12642 13062
rect 12614 12783 12615 12809
rect 12641 12783 12642 12809
rect 12614 12777 12642 12783
rect 12558 12727 12559 12753
rect 12585 12727 12586 12753
rect 12558 12721 12586 12727
rect 12670 12753 12698 12759
rect 12670 12727 12671 12753
rect 12697 12727 12698 12753
rect 12670 12474 12698 12727
rect 12726 12754 12754 13118
rect 12894 13099 12922 13118
rect 13286 13090 13314 13095
rect 13286 13043 13314 13062
rect 14350 13089 14378 13510
rect 18830 13538 18858 13543
rect 18830 13491 18858 13510
rect 14574 13146 14602 13151
rect 14602 13118 14658 13146
rect 14574 13099 14602 13118
rect 14350 13063 14351 13089
rect 14377 13063 14378 13089
rect 14350 13057 14378 13063
rect 14294 12810 14322 12815
rect 14070 12782 14294 12810
rect 12838 12754 12866 12759
rect 12726 12753 12866 12754
rect 12726 12727 12839 12753
rect 12865 12727 12866 12753
rect 12726 12726 12866 12727
rect 12726 12586 12754 12726
rect 12838 12721 12866 12726
rect 13230 12697 13258 12703
rect 13230 12671 13231 12697
rect 13257 12671 13258 12697
rect 12726 12553 12754 12558
rect 13062 12586 13090 12591
rect 13090 12558 13146 12586
rect 13062 12553 13090 12558
rect 13006 12474 13034 12479
rect 12670 12446 12754 12474
rect 12446 12441 12474 12446
rect 12726 12418 12754 12446
rect 12838 12418 12866 12423
rect 12726 12417 12866 12418
rect 12726 12391 12839 12417
rect 12865 12391 12866 12417
rect 12726 12390 12866 12391
rect 12502 12362 12530 12367
rect 11998 12306 12026 12311
rect 11550 12305 12026 12306
rect 11550 12279 11999 12305
rect 12025 12279 12026 12305
rect 11550 12278 12026 12279
rect 11494 11970 11522 11975
rect 11494 11923 11522 11942
rect 11550 11913 11578 12278
rect 11998 12273 12026 12278
rect 12502 12081 12530 12334
rect 12670 12361 12698 12367
rect 12670 12335 12671 12361
rect 12697 12335 12698 12361
rect 12670 12306 12698 12335
rect 12838 12306 12866 12390
rect 12950 12306 12978 12311
rect 12838 12278 12950 12306
rect 12670 12273 12698 12278
rect 12950 12273 12978 12278
rect 12502 12055 12503 12081
rect 12529 12055 12530 12081
rect 12502 12049 12530 12055
rect 11550 11887 11551 11913
rect 11577 11887 11578 11913
rect 11550 11881 11578 11887
rect 11830 11969 11858 11975
rect 11830 11943 11831 11969
rect 11857 11943 11858 11969
rect 11662 11857 11690 11863
rect 11662 11831 11663 11857
rect 11689 11831 11690 11857
rect 11214 11662 11410 11690
rect 11158 11634 11186 11639
rect 11214 11634 11242 11662
rect 11186 11606 11242 11634
rect 11158 11587 11186 11606
rect 11326 11578 11354 11597
rect 11326 11545 11354 11550
rect 11326 11466 11354 11471
rect 10934 11103 10935 11129
rect 10961 11103 10962 11129
rect 10710 11074 10738 11079
rect 10654 11018 10682 11023
rect 10654 10513 10682 10990
rect 10654 10487 10655 10513
rect 10681 10487 10682 10513
rect 10654 10481 10682 10487
rect 10710 10010 10738 11046
rect 10934 11018 10962 11103
rect 10934 10985 10962 10990
rect 10990 11185 11018 11191
rect 10990 11159 10991 11185
rect 11017 11159 11018 11185
rect 10822 10458 10850 10463
rect 10822 10402 10850 10430
rect 10990 10402 11018 11159
rect 11270 11129 11298 11135
rect 11270 11103 11271 11129
rect 11297 11103 11298 11129
rect 10822 10401 10906 10402
rect 10822 10375 10823 10401
rect 10849 10375 10906 10401
rect 10822 10374 10906 10375
rect 10822 10369 10850 10374
rect 10710 9982 10794 10010
rect 10206 9618 10234 9623
rect 10206 9226 10234 9590
rect 10318 9506 10346 9511
rect 10318 9505 10402 9506
rect 10318 9479 10319 9505
rect 10345 9479 10402 9505
rect 10318 9478 10402 9479
rect 10318 9473 10346 9478
rect 10206 9225 10346 9226
rect 10206 9199 10207 9225
rect 10233 9199 10346 9225
rect 10206 9198 10346 9199
rect 10206 9193 10234 9198
rect 10150 8807 10151 8833
rect 10177 8807 10178 8833
rect 10150 8801 10178 8807
rect 9870 8778 9898 8783
rect 9758 8415 9759 8441
rect 9785 8415 9786 8441
rect 9534 8386 9562 8414
rect 9758 8409 9786 8415
rect 9814 8777 9898 8778
rect 9814 8751 9871 8777
rect 9897 8751 9898 8777
rect 9814 8750 9898 8751
rect 9534 8050 9562 8358
rect 9814 8050 9842 8750
rect 9870 8745 9898 8750
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9926 8554 9954 8559
rect 9534 8017 9562 8022
rect 9758 8022 9842 8050
rect 9870 8050 9898 8055
rect 9310 7961 9338 7966
rect 9590 7994 9618 7999
rect 8974 7937 9002 7943
rect 8974 7911 8975 7937
rect 9001 7911 9002 7937
rect 8974 7266 9002 7911
rect 9534 7714 9562 7719
rect 9590 7714 9618 7966
rect 9534 7713 9618 7714
rect 9534 7687 9535 7713
rect 9561 7687 9618 7713
rect 9534 7686 9618 7687
rect 9534 7681 9562 7686
rect 9702 7657 9730 7663
rect 9702 7631 9703 7657
rect 9729 7631 9730 7657
rect 9590 7602 9618 7621
rect 9590 7569 9618 7574
rect 9702 7378 9730 7631
rect 9758 7658 9786 8022
rect 9870 8003 9898 8022
rect 9926 7938 9954 8526
rect 10318 8553 10346 9198
rect 10318 8527 10319 8553
rect 10345 8527 10346 8553
rect 10318 8521 10346 8527
rect 10374 8778 10402 9478
rect 10598 8946 10626 9646
rect 10766 9170 10794 9982
rect 10878 9450 10906 10374
rect 10990 10369 11018 10374
rect 11158 10793 11186 10799
rect 11158 10767 11159 10793
rect 11185 10767 11186 10793
rect 11158 10401 11186 10767
rect 11270 10682 11298 11103
rect 11326 11074 11354 11438
rect 11382 11185 11410 11662
rect 11382 11159 11383 11185
rect 11409 11159 11410 11185
rect 11382 11153 11410 11159
rect 11662 11578 11690 11831
rect 11830 11774 11858 11943
rect 12222 11969 12250 11975
rect 12222 11943 12223 11969
rect 12249 11943 12250 11969
rect 11830 11746 12082 11774
rect 12054 11690 12082 11746
rect 12054 11643 12082 11662
rect 11662 11186 11690 11550
rect 11886 11578 11914 11583
rect 11830 11186 11858 11191
rect 11662 11185 11858 11186
rect 11662 11159 11663 11185
rect 11689 11159 11831 11185
rect 11857 11159 11858 11185
rect 11662 11158 11858 11159
rect 11662 11153 11690 11158
rect 11830 11153 11858 11158
rect 11326 11041 11354 11046
rect 11550 11130 11578 11135
rect 11550 10905 11578 11102
rect 11550 10879 11551 10905
rect 11577 10879 11578 10905
rect 11550 10873 11578 10879
rect 11830 11074 11858 11079
rect 11830 10849 11858 11046
rect 11830 10823 11831 10849
rect 11857 10823 11858 10849
rect 11830 10817 11858 10823
rect 11662 10793 11690 10799
rect 11662 10767 11663 10793
rect 11689 10767 11690 10793
rect 11662 10738 11690 10767
rect 11494 10682 11522 10687
rect 11270 10681 11522 10682
rect 11270 10655 11495 10681
rect 11521 10655 11522 10681
rect 11270 10654 11522 10655
rect 11158 10375 11159 10401
rect 11185 10375 11186 10401
rect 10934 10346 10962 10351
rect 10934 10299 10962 10318
rect 11158 10065 11186 10375
rect 11158 10039 11159 10065
rect 11185 10039 11186 10065
rect 11158 10033 11186 10039
rect 11494 10010 11522 10654
rect 11382 9982 11522 10010
rect 10990 9617 11018 9623
rect 10990 9591 10991 9617
rect 11017 9591 11018 9617
rect 10934 9562 10962 9567
rect 10934 9515 10962 9534
rect 10878 9422 10962 9450
rect 10934 9225 10962 9422
rect 10934 9199 10935 9225
rect 10961 9199 10962 9225
rect 10934 9193 10962 9199
rect 10990 9226 11018 9591
rect 10822 9170 10850 9175
rect 10766 9142 10822 9170
rect 10710 9114 10738 9119
rect 10654 8946 10682 8951
rect 10598 8945 10682 8946
rect 10598 8919 10655 8945
rect 10681 8919 10682 8945
rect 10598 8918 10682 8919
rect 10654 8913 10682 8918
rect 10710 8945 10738 9086
rect 10710 8919 10711 8945
rect 10737 8919 10738 8945
rect 10710 8913 10738 8919
rect 10822 8945 10850 9142
rect 10990 9114 11018 9198
rect 11158 9562 11186 9567
rect 11158 9338 11186 9534
rect 11158 9225 11186 9310
rect 11326 9282 11354 9287
rect 11326 9235 11354 9254
rect 11158 9199 11159 9225
rect 11185 9199 11186 9225
rect 11158 9193 11186 9199
rect 10822 8919 10823 8945
rect 10849 8919 10850 8945
rect 10822 8913 10850 8919
rect 10878 9086 11018 9114
rect 11046 9169 11074 9175
rect 11046 9143 11047 9169
rect 11073 9143 11074 9169
rect 10878 8945 10906 9086
rect 10878 8919 10879 8945
rect 10905 8919 10906 8945
rect 10878 8913 10906 8919
rect 10374 8442 10402 8750
rect 10430 8442 10458 8447
rect 10374 8414 10430 8442
rect 10430 8409 10458 8414
rect 10934 8442 10962 8447
rect 9982 8386 10010 8391
rect 9982 7994 10010 8358
rect 10206 8386 10234 8391
rect 10206 8339 10234 8358
rect 9982 7947 10010 7966
rect 10374 8329 10402 8335
rect 10374 8303 10375 8329
rect 10401 8303 10402 8329
rect 9814 7910 9954 7938
rect 9814 7770 9842 7910
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9814 7742 9898 7770
rect 9814 7658 9842 7663
rect 9758 7630 9814 7658
rect 9814 7611 9842 7630
rect 9814 7546 9842 7551
rect 9870 7546 9898 7742
rect 9814 7545 9898 7546
rect 9814 7519 9815 7545
rect 9841 7519 9898 7545
rect 9814 7518 9898 7519
rect 10206 7658 10234 7663
rect 9814 7513 9842 7518
rect 9758 7378 9786 7383
rect 9702 7377 9786 7378
rect 9702 7351 9759 7377
rect 9785 7351 9786 7377
rect 9702 7350 9786 7351
rect 9758 7345 9786 7350
rect 10206 7377 10234 7630
rect 10206 7351 10207 7377
rect 10233 7351 10234 7377
rect 10206 7345 10234 7351
rect 10374 7658 10402 8303
rect 8974 6538 9002 7238
rect 9590 7321 9618 7327
rect 9590 7295 9591 7321
rect 9617 7295 9618 7321
rect 9590 7210 9618 7295
rect 10374 7265 10402 7630
rect 10766 7658 10794 7663
rect 10654 7602 10682 7621
rect 10766 7611 10794 7630
rect 10654 7569 10682 7574
rect 10598 7545 10626 7551
rect 10598 7519 10599 7545
rect 10625 7519 10626 7545
rect 10598 7322 10626 7519
rect 10822 7546 10850 7551
rect 10822 7545 10906 7546
rect 10822 7519 10823 7545
rect 10849 7519 10906 7545
rect 10822 7518 10906 7519
rect 10822 7513 10850 7518
rect 10710 7322 10738 7327
rect 10598 7321 10738 7322
rect 10598 7295 10711 7321
rect 10737 7295 10738 7321
rect 10598 7294 10738 7295
rect 10710 7289 10738 7294
rect 10374 7239 10375 7265
rect 10401 7239 10402 7265
rect 10374 7233 10402 7239
rect 10766 7265 10794 7271
rect 10766 7239 10767 7265
rect 10793 7239 10794 7265
rect 9814 7210 9842 7215
rect 9590 7209 9842 7210
rect 9590 7183 9815 7209
rect 9841 7183 9842 7209
rect 9590 7182 9842 7183
rect 9758 6986 9786 6991
rect 9702 6958 9758 6986
rect 9702 6929 9730 6958
rect 9758 6953 9786 6958
rect 9702 6903 9703 6929
rect 9729 6903 9730 6929
rect 9702 6897 9730 6903
rect 9366 6818 9394 6823
rect 8974 6481 9002 6510
rect 9310 6790 9366 6818
rect 9310 6537 9338 6790
rect 9366 6785 9394 6790
rect 9646 6817 9674 6823
rect 9646 6791 9647 6817
rect 9673 6791 9674 6817
rect 9646 6706 9674 6791
rect 9646 6673 9674 6678
rect 9310 6511 9311 6537
rect 9337 6511 9338 6537
rect 9310 6505 9338 6511
rect 8974 6455 8975 6481
rect 9001 6455 9002 6481
rect 8974 6449 9002 6455
rect 8750 4186 8890 4214
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 8862 2169 8890 4186
rect 8862 2143 8863 2169
rect 8889 2143 8890 2169
rect 8862 2137 8890 2143
rect 8750 2058 8778 2063
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8750 400 8778 2030
rect 9366 2058 9394 2063
rect 9366 2011 9394 2030
rect 9814 1778 9842 7182
rect 10654 7209 10682 7215
rect 10654 7183 10655 7209
rect 10681 7183 10682 7209
rect 10038 7154 10066 7159
rect 10038 7153 10122 7154
rect 10038 7127 10039 7153
rect 10065 7127 10122 7153
rect 10038 7126 10122 7127
rect 10038 7121 10066 7126
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9982 6986 10010 6991
rect 9982 6939 10010 6958
rect 10038 6930 10066 6935
rect 10038 6883 10066 6902
rect 9870 6873 9898 6879
rect 9870 6847 9871 6873
rect 9897 6847 9898 6873
rect 9870 6762 9898 6847
rect 9926 6818 9954 6823
rect 9926 6771 9954 6790
rect 9870 6729 9898 6734
rect 10094 6538 10122 7126
rect 10262 7153 10290 7159
rect 10262 7127 10263 7153
rect 10289 7127 10290 7153
rect 10262 6873 10290 7127
rect 10598 6930 10626 6935
rect 10654 6930 10682 7183
rect 10626 6902 10682 6930
rect 10598 6897 10626 6902
rect 10262 6847 10263 6873
rect 10289 6847 10290 6873
rect 10262 6841 10290 6847
rect 10486 6874 10514 6879
rect 10486 6827 10514 6846
rect 10766 6818 10794 7239
rect 10822 6930 10850 6935
rect 10878 6930 10906 7518
rect 10822 6929 10906 6930
rect 10822 6903 10823 6929
rect 10849 6903 10906 6929
rect 10822 6902 10906 6903
rect 10934 7265 10962 8414
rect 11046 8386 11074 9143
rect 11382 8497 11410 9982
rect 11494 9618 11522 9623
rect 11494 9571 11522 9590
rect 11494 9394 11522 9399
rect 11438 9338 11466 9343
rect 11438 8833 11466 9310
rect 11494 8890 11522 9366
rect 11662 9282 11690 10710
rect 11774 10346 11802 10351
rect 11718 9618 11746 9623
rect 11774 9618 11802 10318
rect 11886 10122 11914 11550
rect 12222 11578 12250 11943
rect 12222 11545 12250 11550
rect 12334 11969 12362 11975
rect 12334 11943 12335 11969
rect 12361 11943 12362 11969
rect 12334 11858 12362 11943
rect 11998 11073 12026 11079
rect 11998 11047 11999 11073
rect 12025 11047 12026 11073
rect 11998 10906 12026 11047
rect 11998 10873 12026 10878
rect 12222 10906 12250 10911
rect 11942 10850 11970 10855
rect 11942 10803 11970 10822
rect 11998 10794 12026 10799
rect 11998 10747 12026 10766
rect 12054 10793 12082 10799
rect 12054 10767 12055 10793
rect 12081 10767 12082 10793
rect 11886 10089 11914 10094
rect 11718 9617 11802 9618
rect 11718 9591 11719 9617
rect 11745 9591 11802 9617
rect 11718 9590 11802 9591
rect 11718 9585 11746 9590
rect 12054 9562 12082 10767
rect 12110 10793 12138 10799
rect 12110 10767 12111 10793
rect 12137 10767 12138 10793
rect 12110 10738 12138 10767
rect 12110 10705 12138 10710
rect 12166 10066 12194 10071
rect 12110 9730 12138 9735
rect 12110 9683 12138 9702
rect 12054 9529 12082 9534
rect 11942 9338 11970 9343
rect 11942 9291 11970 9310
rect 11662 9249 11690 9254
rect 11662 9170 11690 9175
rect 11662 9123 11690 9142
rect 11774 9114 11802 9119
rect 11718 9113 11802 9114
rect 11718 9087 11775 9113
rect 11801 9087 11802 9113
rect 11718 9086 11802 9087
rect 11494 8843 11522 8862
rect 11606 8946 11634 8951
rect 11718 8946 11746 9086
rect 11774 9081 11802 9086
rect 11606 8945 11746 8946
rect 11606 8919 11607 8945
rect 11633 8919 11746 8945
rect 11606 8918 11746 8919
rect 11438 8807 11439 8833
rect 11465 8807 11466 8833
rect 11438 8801 11466 8807
rect 11606 8554 11634 8918
rect 11606 8521 11634 8526
rect 11382 8471 11383 8497
rect 11409 8471 11410 8497
rect 11382 8465 11410 8471
rect 11494 8497 11522 8503
rect 11494 8471 11495 8497
rect 11521 8471 11522 8497
rect 11494 8442 11522 8471
rect 11494 8409 11522 8414
rect 12110 8498 12138 8503
rect 12166 8498 12194 10038
rect 12110 8497 12194 8498
rect 12110 8471 12111 8497
rect 12137 8471 12194 8497
rect 12110 8470 12194 8471
rect 12222 8553 12250 10878
rect 12334 9730 12362 11830
rect 12614 11690 12642 11695
rect 12614 10066 12642 11662
rect 13006 11522 13034 12446
rect 13062 12362 13090 12367
rect 13062 12315 13090 12334
rect 13118 12194 13146 12558
rect 13174 12474 13202 12479
rect 13174 12427 13202 12446
rect 13230 12473 13258 12671
rect 13230 12447 13231 12473
rect 13257 12447 13258 12473
rect 13230 12441 13258 12447
rect 14070 12417 14098 12782
rect 14294 12763 14322 12782
rect 14630 12809 14658 13118
rect 18830 13145 18858 13151
rect 18830 13119 18831 13145
rect 18857 13119 18858 13145
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 14630 12783 14631 12809
rect 14657 12783 14658 12809
rect 14630 12777 14658 12783
rect 18830 12810 18858 13119
rect 20006 13146 20034 13567
rect 20006 13113 20034 13118
rect 18830 12777 18858 12782
rect 20006 13033 20034 13039
rect 20006 13007 20007 13033
rect 20033 13007 20034 13033
rect 20006 12810 20034 13007
rect 20006 12777 20034 12782
rect 14070 12391 14071 12417
rect 14097 12391 14098 12417
rect 14070 12385 14098 12391
rect 13286 12362 13314 12367
rect 13286 12315 13314 12334
rect 13398 12361 13426 12367
rect 13398 12335 13399 12361
rect 13425 12335 13426 12361
rect 13398 12306 13426 12335
rect 14014 12362 14042 12367
rect 14014 12315 14042 12334
rect 13118 12166 13258 12194
rect 13230 11690 13258 12166
rect 13398 11746 13426 12278
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 13398 11718 13538 11746
rect 13230 11689 13426 11690
rect 13230 11663 13231 11689
rect 13257 11663 13426 11689
rect 13230 11662 13426 11663
rect 13230 11657 13258 11662
rect 13398 11578 13426 11662
rect 13398 11577 13482 11578
rect 13398 11551 13399 11577
rect 13425 11551 13482 11577
rect 13398 11550 13482 11551
rect 13398 11545 13426 11550
rect 12838 11494 13034 11522
rect 12726 11074 12754 11079
rect 12726 10905 12754 11046
rect 12726 10879 12727 10905
rect 12753 10879 12754 10905
rect 12726 10873 12754 10879
rect 12614 10019 12642 10038
rect 12838 10065 12866 11494
rect 13230 11186 13258 11191
rect 13118 11018 13146 11023
rect 13118 10905 13146 10990
rect 13118 10879 13119 10905
rect 13145 10879 13146 10905
rect 13118 10873 13146 10879
rect 12894 10794 12922 10799
rect 12894 10747 12922 10766
rect 13006 10793 13034 10799
rect 13006 10767 13007 10793
rect 13033 10767 13034 10793
rect 13006 10626 13034 10767
rect 13230 10793 13258 11158
rect 13286 11130 13314 11135
rect 13286 11083 13314 11102
rect 13230 10767 13231 10793
rect 13257 10767 13258 10793
rect 13230 10761 13258 10767
rect 13398 11073 13426 11079
rect 13398 11047 13399 11073
rect 13425 11047 13426 11073
rect 13062 10738 13090 10743
rect 13062 10691 13090 10710
rect 13398 10626 13426 11047
rect 13006 10598 13426 10626
rect 13398 10121 13426 10598
rect 13398 10095 13399 10121
rect 13425 10095 13426 10121
rect 13398 10089 13426 10095
rect 13454 11074 13482 11550
rect 13510 11186 13538 11718
rect 13790 11522 13818 11527
rect 14854 11522 14882 11527
rect 13566 11521 13818 11522
rect 13566 11495 13791 11521
rect 13817 11495 13818 11521
rect 13566 11494 13818 11495
rect 13566 11241 13594 11494
rect 13790 11489 13818 11494
rect 14798 11521 14882 11522
rect 14798 11495 14855 11521
rect 14881 11495 14882 11521
rect 14798 11494 14882 11495
rect 13566 11215 13567 11241
rect 13593 11215 13594 11241
rect 13566 11209 13594 11215
rect 13510 11153 13538 11158
rect 13622 11186 13650 11191
rect 13622 11139 13650 11158
rect 14630 11129 14658 11135
rect 14630 11103 14631 11129
rect 14657 11103 14658 11129
rect 13454 10793 13482 11046
rect 13454 10767 13455 10793
rect 13481 10767 13482 10793
rect 13454 10457 13482 10767
rect 13510 11073 13538 11079
rect 13510 11047 13511 11073
rect 13537 11047 13538 11073
rect 13510 10514 13538 11047
rect 14014 11074 14042 11079
rect 13790 10738 13818 10743
rect 13790 10691 13818 10710
rect 13510 10481 13538 10486
rect 13454 10431 13455 10457
rect 13481 10431 13482 10457
rect 13454 10094 13482 10431
rect 14014 10457 14042 11046
rect 14574 11073 14602 11079
rect 14574 11047 14575 11073
rect 14601 11047 14602 11073
rect 14574 11018 14602 11047
rect 14574 10985 14602 10990
rect 14630 10962 14658 11103
rect 14630 10929 14658 10934
rect 14574 10514 14602 10519
rect 14574 10467 14602 10486
rect 14014 10431 14015 10457
rect 14041 10431 14042 10457
rect 14014 10425 14042 10431
rect 14630 10346 14658 10351
rect 14798 10346 14826 11494
rect 14854 11489 14882 11494
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 18830 11185 18858 11191
rect 18830 11159 18831 11185
rect 18857 11159 18858 11185
rect 14854 10962 14882 10967
rect 14854 10737 14882 10934
rect 18830 10962 18858 11159
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 18830 10929 18858 10934
rect 14854 10711 14855 10737
rect 14881 10711 14882 10737
rect 14854 10705 14882 10711
rect 18830 10793 18858 10799
rect 18830 10767 18831 10793
rect 18857 10767 18858 10793
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 14854 10346 14882 10351
rect 14798 10318 14854 10346
rect 14630 10299 14658 10318
rect 14854 10313 14882 10318
rect 18830 10346 18858 10767
rect 20006 10794 20034 10799
rect 20006 10737 20034 10766
rect 20006 10711 20007 10737
rect 20033 10711 20034 10737
rect 20006 10705 20034 10711
rect 18830 10313 18858 10318
rect 13454 10066 13594 10094
rect 12838 10039 12839 10065
rect 12865 10039 12866 10065
rect 12334 9697 12362 9702
rect 12726 10009 12754 10015
rect 12726 9983 12727 10009
rect 12753 9983 12754 10009
rect 12726 9730 12754 9983
rect 12726 9697 12754 9702
rect 12670 9562 12698 9567
rect 12698 9534 12754 9562
rect 12670 9515 12698 9534
rect 12502 9505 12530 9511
rect 12502 9479 12503 9505
rect 12529 9479 12530 9505
rect 12502 9450 12530 9479
rect 12502 9417 12530 9422
rect 12726 9394 12754 9534
rect 12838 9561 12866 10039
rect 12894 10010 12922 10015
rect 12894 9963 12922 9982
rect 13230 10010 13258 10015
rect 13230 9963 13258 9982
rect 13566 10009 13594 10066
rect 18830 10010 18858 10015
rect 13566 9983 13567 10009
rect 13593 9983 13594 10009
rect 13118 9953 13146 9959
rect 13118 9927 13119 9953
rect 13145 9927 13146 9953
rect 12894 9898 12922 9903
rect 12894 9851 12922 9870
rect 12838 9535 12839 9561
rect 12865 9535 12866 9561
rect 12838 9529 12866 9535
rect 12950 9506 12978 9511
rect 12726 9366 12866 9394
rect 12838 9337 12866 9366
rect 12838 9311 12839 9337
rect 12865 9311 12866 9337
rect 12838 9305 12866 9311
rect 12782 9282 12810 9287
rect 12782 9235 12810 9254
rect 12838 9113 12866 9119
rect 12838 9087 12839 9113
rect 12865 9087 12866 9113
rect 12614 8834 12642 8839
rect 12390 8833 12642 8834
rect 12390 8807 12615 8833
rect 12641 8807 12642 8833
rect 12390 8806 12642 8807
rect 12222 8527 12223 8553
rect 12249 8527 12250 8553
rect 11046 8353 11074 8358
rect 11494 8330 11522 8335
rect 11382 7993 11410 7999
rect 11382 7967 11383 7993
rect 11409 7967 11410 7993
rect 11382 7658 11410 7967
rect 11438 7994 11466 7999
rect 11494 7994 11522 8302
rect 11550 8330 11578 8335
rect 11550 8329 11802 8330
rect 11550 8303 11551 8329
rect 11577 8303 11802 8329
rect 11550 8302 11802 8303
rect 11550 8297 11578 8302
rect 11550 8050 11578 8055
rect 11550 8049 11690 8050
rect 11550 8023 11551 8049
rect 11577 8023 11690 8049
rect 11550 8022 11690 8023
rect 11550 8017 11578 8022
rect 11438 7993 11522 7994
rect 11438 7967 11439 7993
rect 11465 7967 11522 7993
rect 11438 7966 11522 7967
rect 11662 7993 11690 8022
rect 11774 8049 11802 8302
rect 11774 8023 11775 8049
rect 11801 8023 11802 8049
rect 11774 8017 11802 8023
rect 11942 8049 11970 8055
rect 11942 8023 11943 8049
rect 11969 8023 11970 8049
rect 11662 7967 11663 7993
rect 11689 7967 11690 7993
rect 11438 7961 11466 7966
rect 11662 7961 11690 7967
rect 11382 7625 11410 7630
rect 11606 7937 11634 7943
rect 11606 7911 11607 7937
rect 11633 7911 11634 7937
rect 11606 7574 11634 7911
rect 11942 7882 11970 8023
rect 12110 8049 12138 8470
rect 12222 8330 12250 8527
rect 12334 8554 12362 8559
rect 12334 8507 12362 8526
rect 12390 8385 12418 8806
rect 12614 8801 12642 8806
rect 12838 8833 12866 9087
rect 12838 8807 12839 8833
rect 12865 8807 12866 8833
rect 12838 8801 12866 8807
rect 12950 8834 12978 9478
rect 13006 9506 13034 9511
rect 13118 9506 13146 9927
rect 13510 9898 13538 9903
rect 13174 9674 13202 9679
rect 13174 9617 13202 9646
rect 13174 9591 13175 9617
rect 13201 9591 13202 9617
rect 13174 9585 13202 9591
rect 13510 9617 13538 9870
rect 13510 9591 13511 9617
rect 13537 9591 13538 9617
rect 13510 9585 13538 9591
rect 13006 9505 13146 9506
rect 13006 9479 13007 9505
rect 13033 9479 13146 9505
rect 13006 9478 13146 9479
rect 13342 9506 13370 9511
rect 13006 9338 13034 9478
rect 13342 9459 13370 9478
rect 13454 9506 13482 9511
rect 13006 9305 13034 9310
rect 13286 9394 13314 9399
rect 13286 9281 13314 9366
rect 13454 9337 13482 9478
rect 13454 9311 13455 9337
rect 13481 9311 13482 9337
rect 13454 9305 13482 9311
rect 13286 9255 13287 9281
rect 13313 9255 13314 9281
rect 13286 9249 13314 9255
rect 13342 9281 13370 9287
rect 13342 9255 13343 9281
rect 13369 9255 13370 9281
rect 13342 9226 13370 9255
rect 13342 9193 13370 9198
rect 13566 9225 13594 9983
rect 18774 10009 18858 10010
rect 18774 9983 18831 10009
rect 18857 9983 18858 10009
rect 18774 9982 18858 9983
rect 13958 9954 13986 9959
rect 13846 9953 13986 9954
rect 13846 9927 13959 9953
rect 13985 9927 13986 9953
rect 13846 9926 13986 9927
rect 13790 9673 13818 9679
rect 13790 9647 13791 9673
rect 13817 9647 13818 9673
rect 13790 9618 13818 9647
rect 13790 9585 13818 9590
rect 13734 9562 13762 9567
rect 13622 9506 13650 9511
rect 13622 9459 13650 9478
rect 13734 9450 13762 9534
rect 13734 9417 13762 9422
rect 13790 9506 13818 9511
rect 13566 9199 13567 9225
rect 13593 9199 13594 9225
rect 12950 8787 12978 8806
rect 13118 9170 13146 9175
rect 12782 8722 12810 8727
rect 12782 8721 12922 8722
rect 12782 8695 12783 8721
rect 12809 8695 12922 8721
rect 12782 8694 12922 8695
rect 12782 8689 12810 8694
rect 12894 8554 12922 8694
rect 12894 8526 13034 8554
rect 13006 8497 13034 8526
rect 13006 8471 13007 8497
rect 13033 8471 13034 8497
rect 13006 8465 13034 8471
rect 12390 8359 12391 8385
rect 12417 8359 12418 8385
rect 12390 8353 12418 8359
rect 12670 8442 12698 8447
rect 12250 8302 12306 8330
rect 12222 8297 12250 8302
rect 12110 8023 12111 8049
rect 12137 8023 12138 8049
rect 12110 8017 12138 8023
rect 12166 8105 12194 8111
rect 12166 8079 12167 8105
rect 12193 8079 12194 8105
rect 12166 7882 12194 8079
rect 12222 7938 12250 7943
rect 12278 7938 12306 8302
rect 12222 7937 12306 7938
rect 12222 7911 12223 7937
rect 12249 7911 12306 7937
rect 12222 7910 12306 7911
rect 12334 7938 12362 7943
rect 12222 7905 12250 7910
rect 12334 7891 12362 7910
rect 11942 7854 12194 7882
rect 11606 7546 11746 7574
rect 11718 7518 11914 7546
rect 11886 7321 11914 7518
rect 11886 7295 11887 7321
rect 11913 7295 11914 7321
rect 11886 7289 11914 7295
rect 10934 7239 10935 7265
rect 10961 7239 10962 7265
rect 10822 6897 10850 6902
rect 10822 6818 10850 6823
rect 10766 6790 10822 6818
rect 10822 6785 10850 6790
rect 10934 6762 10962 7239
rect 11494 7265 11522 7271
rect 11494 7239 11495 7265
rect 11521 7239 11522 7265
rect 11494 6874 11522 7239
rect 12334 6929 12362 6935
rect 12334 6903 12335 6929
rect 12361 6903 12362 6929
rect 11494 6841 11522 6846
rect 12110 6874 12138 6879
rect 10934 6729 10962 6734
rect 11606 6818 11634 6823
rect 10094 6505 10122 6510
rect 10374 6706 10402 6711
rect 10374 6537 10402 6678
rect 10374 6511 10375 6537
rect 10401 6511 10402 6537
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 10374 4214 10402 6511
rect 10710 6538 10738 6543
rect 10710 6491 10738 6510
rect 11606 6481 11634 6790
rect 11942 6818 11970 6823
rect 11942 6771 11970 6790
rect 12110 6538 12138 6846
rect 12166 6873 12194 6879
rect 12166 6847 12167 6873
rect 12193 6847 12194 6873
rect 12166 6818 12194 6847
rect 12166 6785 12194 6790
rect 12166 6538 12194 6543
rect 12110 6537 12194 6538
rect 12110 6511 12167 6537
rect 12193 6511 12194 6537
rect 12110 6510 12194 6511
rect 12166 6505 12194 6510
rect 11606 6455 11607 6481
rect 11633 6455 11634 6481
rect 11606 5866 11634 6455
rect 11718 6370 11746 6375
rect 11718 6369 11914 6370
rect 11718 6343 11719 6369
rect 11745 6343 11914 6369
rect 11718 6342 11914 6343
rect 11718 6337 11746 6342
rect 11606 5838 11802 5866
rect 10374 4186 10570 4214
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 10542 2169 10570 4186
rect 10542 2143 10543 2169
rect 10569 2143 10570 2169
rect 10542 2137 10570 2143
rect 10430 2058 10458 2063
rect 9870 1778 9898 1783
rect 9814 1777 9898 1778
rect 9814 1751 9871 1777
rect 9897 1751 9898 1777
rect 9814 1750 9898 1751
rect 9870 1745 9898 1750
rect 9590 1666 9618 1671
rect 9590 1665 9786 1666
rect 9590 1639 9591 1665
rect 9617 1639 9786 1665
rect 9590 1638 9786 1639
rect 9590 1633 9618 1638
rect 9758 400 9786 1638
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10430 400 10458 2030
rect 11046 2058 11074 2063
rect 11046 2011 11074 2030
rect 11438 1834 11466 1839
rect 11102 1721 11130 1727
rect 11102 1695 11103 1721
rect 11129 1695 11130 1721
rect 11102 400 11130 1695
rect 11438 400 11466 1806
rect 11774 1777 11802 5838
rect 11774 1751 11775 1777
rect 11801 1751 11802 1777
rect 11774 1745 11802 1751
rect 11830 2618 11858 2623
rect 11830 490 11858 2590
rect 11886 2561 11914 6342
rect 12334 4214 12362 6903
rect 12670 6874 12698 8414
rect 13118 8442 13146 9142
rect 13566 9170 13594 9199
rect 13566 9137 13594 9142
rect 13734 8834 13762 8839
rect 13790 8834 13818 9478
rect 13846 8889 13874 9926
rect 13958 9921 13986 9926
rect 14182 9954 14210 9959
rect 13958 9618 13986 9623
rect 13846 8863 13847 8889
rect 13873 8863 13874 8889
rect 13846 8857 13874 8863
rect 13902 9450 13930 9455
rect 13762 8806 13818 8834
rect 13902 8833 13930 9422
rect 13958 9281 13986 9590
rect 14182 9617 14210 9926
rect 15022 9954 15050 9959
rect 15022 9907 15050 9926
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 14182 9591 14183 9617
rect 14209 9591 14210 9617
rect 14182 9585 14210 9591
rect 14238 9617 14266 9623
rect 14238 9591 14239 9617
rect 14265 9591 14266 9617
rect 13958 9255 13959 9281
rect 13985 9255 13986 9281
rect 13958 9249 13986 9255
rect 14014 9561 14042 9567
rect 14014 9535 14015 9561
rect 14041 9535 14042 9561
rect 14014 9282 14042 9535
rect 14014 9249 14042 9254
rect 14070 9505 14098 9511
rect 14070 9479 14071 9505
rect 14097 9479 14098 9505
rect 13902 8807 13903 8833
rect 13929 8807 13930 8833
rect 13734 8787 13762 8806
rect 13902 8801 13930 8807
rect 14070 8833 14098 9479
rect 14238 9506 14266 9591
rect 14238 9473 14266 9478
rect 15358 9281 15386 9287
rect 15358 9255 15359 9281
rect 15385 9255 15386 9281
rect 15022 9226 15050 9231
rect 15022 9169 15050 9198
rect 15246 9226 15274 9231
rect 15246 9179 15274 9198
rect 15022 9143 15023 9169
rect 15049 9143 15050 9169
rect 15022 9137 15050 9143
rect 15358 9170 15386 9255
rect 15358 9137 15386 9142
rect 18774 9170 18802 9982
rect 18830 9977 18858 9982
rect 20006 9897 20034 9903
rect 20006 9871 20007 9897
rect 20033 9871 20034 9897
rect 18830 9842 18858 9847
rect 18830 9225 18858 9814
rect 20006 9786 20034 9871
rect 20006 9753 20034 9758
rect 20006 9673 20034 9679
rect 20006 9647 20007 9673
rect 20033 9647 20034 9673
rect 18830 9199 18831 9225
rect 18857 9199 18858 9225
rect 18830 9193 18858 9199
rect 18942 9617 18970 9623
rect 18942 9591 18943 9617
rect 18969 9591 18970 9617
rect 18942 9226 18970 9591
rect 20006 9450 20034 9647
rect 20006 9417 20034 9422
rect 18942 9193 18970 9198
rect 18774 9137 18802 9142
rect 20006 9114 20034 9119
rect 20006 9067 20034 9086
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 14070 8807 14071 8833
rect 14097 8807 14098 8833
rect 14070 8801 14098 8807
rect 14126 8834 14154 8839
rect 13118 8409 13146 8414
rect 14126 8554 14154 8806
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 14070 8386 14098 8391
rect 14126 8386 14154 8526
rect 14294 8442 14322 8447
rect 14294 8395 14322 8414
rect 20006 8442 20034 8863
rect 20006 8409 20034 8414
rect 14070 8385 14154 8386
rect 14070 8359 14071 8385
rect 14097 8359 14154 8385
rect 14070 8358 14154 8359
rect 14070 8353 14098 8358
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 12670 6841 12698 6846
rect 12950 7938 12978 7943
rect 12950 7321 12978 7910
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 12950 7295 12951 7321
rect 12977 7295 12978 7321
rect 12950 4214 12978 7295
rect 13174 7153 13202 7159
rect 13174 7127 13175 7153
rect 13201 7127 13202 7153
rect 13174 6874 13202 7127
rect 13174 6841 13202 6846
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 11886 2535 11887 2561
rect 11913 2535 11914 2561
rect 11886 2529 11914 2535
rect 12278 4186 12362 4214
rect 12670 4186 12978 4214
rect 12278 1777 12306 4186
rect 12390 2618 12418 2623
rect 12390 2571 12418 2590
rect 12670 2169 12698 4186
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 12670 2143 12671 2169
rect 12697 2143 12698 2169
rect 12670 2137 12698 2143
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1745 12306 1751
rect 12446 2058 12474 2063
rect 11774 462 11858 490
rect 11774 400 11802 462
rect 12446 400 12474 2030
rect 13118 2058 13146 2063
rect 13118 2011 13146 2030
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 8736 0 8792 400
rect 9744 0 9800 400
rect 10416 0 10472 400
rect 11088 0 11144 400
rect 11424 0 11480 400
rect 11760 0 11816 400
rect 12432 0 12488 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 8414 19110 8442 19138
rect 9030 19137 9058 19138
rect 9030 19111 9031 19137
rect 9031 19111 9057 19137
rect 9057 19111 9058 19137
rect 9030 19110 9058 19111
rect 8078 18718 8106 18746
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 9198 18745 9226 18746
rect 9198 18719 9199 18745
rect 9199 18719 9225 18745
rect 9225 18719 9226 18745
rect 9198 18718 9226 18719
rect 10430 19110 10458 19138
rect 11046 19137 11074 19138
rect 11046 19111 11047 19137
rect 11047 19111 11073 19137
rect 11073 19111 11074 19137
rect 11046 19110 11074 19111
rect 11774 19110 11802 19138
rect 10094 18718 10122 18746
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 7406 13790 7434 13818
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 2086 13454 2114 13482
rect 966 12249 994 12250
rect 966 12223 967 12249
rect 967 12223 993 12249
rect 993 12223 994 12249
rect 966 12222 994 12223
rect 966 11465 994 11466
rect 966 11439 967 11465
rect 967 11439 993 11465
rect 993 11439 994 11465
rect 966 11438 994 11439
rect 966 11241 994 11242
rect 966 11215 967 11241
rect 967 11215 993 11241
rect 993 11215 994 11241
rect 966 11214 994 11215
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 2142 12361 2170 12362
rect 2142 12335 2143 12361
rect 2143 12335 2169 12361
rect 2169 12335 2170 12361
rect 2142 12334 2170 12335
rect 6734 12334 6762 12362
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 6734 12025 6762 12026
rect 6734 11999 6735 12025
rect 6735 11999 6761 12025
rect 6761 11999 6762 12025
rect 6734 11998 6762 11999
rect 6454 11662 6482 11690
rect 5278 11606 5306 11634
rect 2142 11577 2170 11578
rect 2142 11551 2143 11577
rect 2143 11551 2169 11577
rect 2169 11551 2170 11577
rect 2142 11550 2170 11551
rect 6342 11521 6370 11522
rect 6342 11495 6343 11521
rect 6343 11495 6369 11521
rect 6369 11495 6370 11521
rect 6342 11494 6370 11495
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 2142 11185 2170 11186
rect 2142 11159 2143 11185
rect 2143 11159 2169 11185
rect 2169 11159 2170 11185
rect 2142 11158 2170 11159
rect 6734 11662 6762 11690
rect 7294 13089 7322 13090
rect 7294 13063 7295 13089
rect 7295 13063 7321 13089
rect 7321 13063 7322 13089
rect 7294 13062 7322 13063
rect 8022 13817 8050 13818
rect 8022 13791 8023 13817
rect 8023 13791 8049 13817
rect 8049 13791 8050 13817
rect 8022 13790 8050 13791
rect 8806 13873 8834 13874
rect 8806 13847 8807 13873
rect 8807 13847 8833 13873
rect 8833 13847 8834 13873
rect 8806 13846 8834 13847
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 10710 18745 10738 18746
rect 10710 18719 10711 18745
rect 10711 18719 10737 18745
rect 10737 18719 10738 18745
rect 10710 18718 10738 18719
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 12446 18718 12474 18746
rect 13118 18745 13146 18746
rect 13118 18719 13119 18745
rect 13119 18719 13145 18745
rect 13145 18719 13146 18745
rect 13118 18718 13146 18719
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 9086 13846 9114 13874
rect 8358 13286 8386 13314
rect 8358 13174 8386 13202
rect 7910 13062 7938 13090
rect 8078 13006 8106 13034
rect 7742 12670 7770 12698
rect 7070 11662 7098 11690
rect 7406 11886 7434 11914
rect 7574 11662 7602 11690
rect 6958 11633 6986 11634
rect 6958 11607 6959 11633
rect 6959 11607 6985 11633
rect 6985 11607 6986 11633
rect 6958 11606 6986 11607
rect 7014 11577 7042 11578
rect 7014 11551 7015 11577
rect 7015 11551 7041 11577
rect 7041 11551 7042 11577
rect 7014 11550 7042 11551
rect 7294 11550 7322 11578
rect 6790 11494 6818 11522
rect 4998 11102 5026 11130
rect 5390 10766 5418 10794
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 2086 9926 2114 9954
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 6454 10681 6482 10682
rect 6454 10655 6455 10681
rect 6455 10655 6481 10681
rect 6481 10655 6482 10681
rect 6454 10654 6482 10655
rect 7350 11521 7378 11522
rect 7350 11495 7351 11521
rect 7351 11495 7377 11521
rect 7377 11495 7378 11521
rect 7350 11494 7378 11495
rect 7686 11438 7714 11466
rect 7238 11129 7266 11130
rect 7238 11103 7239 11129
rect 7239 11103 7265 11129
rect 7265 11103 7266 11129
rect 7238 11102 7266 11103
rect 7966 11998 7994 12026
rect 7798 11913 7826 11914
rect 7798 11887 7799 11913
rect 7799 11887 7825 11913
rect 7825 11887 7826 11913
rect 7798 11886 7826 11887
rect 7854 11774 7882 11802
rect 9422 13622 9450 13650
rect 10318 13649 10346 13650
rect 10318 13623 10319 13649
rect 10319 13623 10345 13649
rect 10345 13623 10346 13649
rect 10318 13622 10346 13623
rect 8750 13201 8778 13202
rect 8750 13175 8751 13201
rect 8751 13175 8777 13201
rect 8777 13175 8778 13201
rect 8750 13174 8778 13175
rect 8806 13286 8834 13314
rect 10094 13454 10122 13482
rect 9918 13341 9946 13342
rect 9030 13230 9058 13258
rect 9254 13286 9282 13314
rect 8750 13033 8778 13034
rect 8750 13007 8751 13033
rect 8751 13007 8777 13033
rect 8777 13007 8778 13033
rect 8750 13006 8778 13007
rect 9814 13286 9842 13314
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9534 13257 9562 13258
rect 9534 13231 9535 13257
rect 9535 13231 9561 13257
rect 9561 13231 9562 13257
rect 9534 13230 9562 13231
rect 8022 11774 8050 11802
rect 8134 11830 8162 11858
rect 8134 11662 8162 11690
rect 7910 11633 7938 11634
rect 7910 11607 7911 11633
rect 7911 11607 7937 11633
rect 7937 11607 7938 11633
rect 7910 11606 7938 11607
rect 8022 11521 8050 11522
rect 8022 11495 8023 11521
rect 8023 11495 8049 11521
rect 8049 11495 8050 11521
rect 8022 11494 8050 11495
rect 8078 11438 8106 11466
rect 8190 11577 8218 11578
rect 8190 11551 8191 11577
rect 8191 11551 8217 11577
rect 8217 11551 8218 11577
rect 8190 11550 8218 11551
rect 6566 10878 6594 10906
rect 6790 10822 6818 10850
rect 7238 10878 7266 10906
rect 7126 10822 7154 10850
rect 6734 10793 6762 10794
rect 6734 10767 6735 10793
rect 6735 10767 6761 10793
rect 6761 10767 6762 10793
rect 6734 10766 6762 10767
rect 7406 10878 7434 10906
rect 7182 10766 7210 10794
rect 6734 10654 6762 10682
rect 7854 10905 7882 10906
rect 7854 10879 7855 10905
rect 7855 10879 7881 10905
rect 7881 10879 7882 10905
rect 7854 10878 7882 10879
rect 7798 10766 7826 10794
rect 7574 10430 7602 10458
rect 6454 9982 6482 10010
rect 7126 10009 7154 10010
rect 7126 9983 7127 10009
rect 7127 9983 7153 10009
rect 7153 9983 7154 10009
rect 7126 9982 7154 9983
rect 5054 9254 5082 9282
rect 5278 9254 5306 9282
rect 6566 9254 6594 9282
rect 6734 9702 6762 9730
rect 7462 10009 7490 10010
rect 7462 9983 7463 10009
rect 7463 9983 7489 10009
rect 7489 9983 7490 10009
rect 7462 9982 7490 9983
rect 7406 9617 7434 9618
rect 7406 9591 7407 9617
rect 7407 9591 7433 9617
rect 7433 9591 7434 9617
rect 7406 9590 7434 9591
rect 6678 9198 6706 9226
rect 5614 9169 5642 9170
rect 5614 9143 5615 9169
rect 5615 9143 5641 9169
rect 5641 9143 5642 9169
rect 5614 9142 5642 9143
rect 7238 9534 7266 9562
rect 7518 9534 7546 9562
rect 7742 10318 7770 10346
rect 8022 10793 8050 10794
rect 8022 10767 8023 10793
rect 8023 10767 8049 10793
rect 8049 10767 8050 10793
rect 8022 10766 8050 10767
rect 8414 11774 8442 11802
rect 9422 12278 9450 12306
rect 9366 12054 9394 12082
rect 8526 11830 8554 11858
rect 8694 11857 8722 11858
rect 8694 11831 8695 11857
rect 8695 11831 8721 11857
rect 8721 11831 8722 11857
rect 8694 11830 8722 11831
rect 9086 11689 9114 11690
rect 9086 11663 9087 11689
rect 9087 11663 9113 11689
rect 9113 11663 9114 11689
rect 9086 11662 9114 11663
rect 8918 11633 8946 11634
rect 8918 11607 8919 11633
rect 8919 11607 8945 11633
rect 8945 11607 8946 11633
rect 8918 11606 8946 11607
rect 8470 10430 8498 10458
rect 8134 10374 8162 10402
rect 8638 10401 8666 10402
rect 8638 10375 8639 10401
rect 8639 10375 8665 10401
rect 8665 10375 8666 10401
rect 8638 10374 8666 10375
rect 8806 10878 8834 10906
rect 8190 10345 8218 10346
rect 8190 10319 8191 10345
rect 8191 10319 8217 10345
rect 8217 10319 8218 10345
rect 8190 10318 8218 10319
rect 8526 10345 8554 10346
rect 8526 10319 8527 10345
rect 8527 10319 8553 10345
rect 8553 10319 8554 10345
rect 8526 10318 8554 10319
rect 8862 10401 8890 10402
rect 8862 10375 8863 10401
rect 8863 10375 8889 10401
rect 8889 10375 8890 10401
rect 8862 10374 8890 10375
rect 9142 11046 9170 11074
rect 9030 10766 9058 10794
rect 8974 10654 9002 10682
rect 8806 10009 8834 10010
rect 8806 9983 8807 10009
rect 8807 9983 8833 10009
rect 8833 9983 8834 10009
rect 8806 9982 8834 9983
rect 7910 9758 7938 9786
rect 8078 9758 8106 9786
rect 7910 9590 7938 9618
rect 6734 9142 6762 9170
rect 6902 9254 6930 9282
rect 7126 9225 7154 9226
rect 7126 9199 7127 9225
rect 7127 9199 7153 9225
rect 7153 9199 7154 9225
rect 7126 9198 7154 9199
rect 7406 9225 7434 9226
rect 7406 9199 7407 9225
rect 7407 9199 7433 9225
rect 7433 9199 7434 9225
rect 7406 9198 7434 9199
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 8190 9534 8218 9562
rect 8358 9505 8386 9506
rect 8358 9479 8359 9505
rect 8359 9479 8385 9505
rect 8385 9479 8386 9505
rect 8358 9478 8386 9479
rect 7238 8694 7266 8722
rect 7854 8721 7882 8722
rect 7854 8695 7855 8721
rect 7855 8695 7881 8721
rect 7881 8695 7882 8721
rect 7854 8694 7882 8695
rect 7798 8526 7826 8554
rect 8190 8526 8218 8554
rect 7686 8470 7714 8498
rect 6902 8441 6930 8442
rect 6902 8415 6903 8441
rect 6903 8415 6929 8441
rect 6929 8415 6930 8441
rect 6902 8414 6930 8415
rect 7350 8414 7378 8442
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 8358 8358 8386 8386
rect 9198 10289 9226 10290
rect 9198 10263 9199 10289
rect 9199 10263 9225 10289
rect 9225 10263 9226 10289
rect 9198 10262 9226 10263
rect 9366 11830 9394 11858
rect 9422 11662 9450 11690
rect 9926 13257 9954 13258
rect 9926 13231 9927 13257
rect 9927 13231 9953 13257
rect 9953 13231 9954 13257
rect 9926 13230 9954 13231
rect 10262 13481 10290 13482
rect 10262 13455 10263 13481
rect 10263 13455 10289 13481
rect 10289 13455 10290 13481
rect 10262 13454 10290 13455
rect 9870 13201 9898 13202
rect 9870 13175 9871 13201
rect 9871 13175 9897 13201
rect 9897 13175 9898 13201
rect 9870 13174 9898 13175
rect 10150 13201 10178 13202
rect 10150 13175 10151 13201
rect 10151 13175 10177 13201
rect 10177 13175 10178 13201
rect 10150 13174 10178 13175
rect 9702 13145 9730 13146
rect 9702 13119 9703 13145
rect 9703 13119 9729 13145
rect 9729 13119 9730 13145
rect 9702 13118 9730 13119
rect 10318 13145 10346 13146
rect 10318 13119 10319 13145
rect 10319 13119 10345 13145
rect 10345 13119 10346 13145
rect 10318 13118 10346 13119
rect 10710 13873 10738 13874
rect 10710 13847 10711 13873
rect 10711 13847 10737 13873
rect 10737 13847 10738 13873
rect 10710 13846 10738 13847
rect 10486 13230 10514 13258
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9814 12081 9842 12082
rect 9814 12055 9815 12081
rect 9815 12055 9841 12081
rect 9841 12055 9842 12081
rect 9814 12054 9842 12055
rect 10878 12697 10906 12698
rect 10878 12671 10879 12697
rect 10879 12671 10905 12697
rect 10905 12671 10906 12697
rect 10878 12670 10906 12671
rect 10598 12558 10626 12586
rect 9702 11689 9730 11690
rect 9702 11663 9703 11689
rect 9703 11663 9729 11689
rect 9729 11663 9730 11689
rect 9702 11662 9730 11663
rect 9422 11494 9450 11522
rect 9590 11550 9618 11578
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 9814 11662 9842 11690
rect 9534 11270 9562 11298
rect 9758 11382 9786 11410
rect 10430 11886 10458 11914
rect 10206 11606 10234 11634
rect 10318 11633 10346 11634
rect 10318 11607 10319 11633
rect 10319 11607 10345 11633
rect 10345 11607 10346 11633
rect 10318 11606 10346 11607
rect 9982 11550 10010 11578
rect 9814 11270 9842 11298
rect 9870 11494 9898 11522
rect 9646 11102 9674 11130
rect 9814 11073 9842 11074
rect 9814 11047 9815 11073
rect 9815 11047 9841 11073
rect 9841 11047 9842 11073
rect 9814 11046 9842 11047
rect 9982 11214 10010 11242
rect 10374 11550 10402 11578
rect 10934 11969 10962 11970
rect 10934 11943 10935 11969
rect 10935 11943 10961 11969
rect 10961 11943 10962 11969
rect 10934 11942 10962 11943
rect 10822 11857 10850 11858
rect 10822 11831 10823 11857
rect 10823 11831 10849 11857
rect 10849 11831 10850 11857
rect 10822 11830 10850 11831
rect 11438 13230 11466 13258
rect 11942 13566 11970 13594
rect 11158 12697 11186 12698
rect 11158 12671 11159 12697
rect 11159 12671 11185 12697
rect 11185 12671 11186 12697
rect 11158 12670 11186 12671
rect 11046 12558 11074 12586
rect 11214 12614 11242 12642
rect 11046 11913 11074 11914
rect 11046 11887 11047 11913
rect 11047 11887 11073 11913
rect 11073 11887 11074 11913
rect 11046 11886 11074 11887
rect 10990 11830 11018 11858
rect 10934 11662 10962 11690
rect 10766 11577 10794 11578
rect 10766 11551 10767 11577
rect 10767 11551 10793 11577
rect 10793 11551 10794 11577
rect 10766 11550 10794 11551
rect 10878 11550 10906 11578
rect 9926 11129 9954 11130
rect 9926 11103 9927 11129
rect 9927 11103 9953 11129
rect 9953 11103 9954 11129
rect 9926 11102 9954 11103
rect 10094 11382 10122 11410
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 10094 10766 10122 10794
rect 10150 11214 10178 11242
rect 10654 11270 10682 11298
rect 9646 10486 9674 10514
rect 9478 10289 9506 10290
rect 9478 10263 9479 10289
rect 9479 10263 9505 10289
rect 9505 10263 9506 10289
rect 9478 10262 9506 10263
rect 9310 10038 9338 10066
rect 9422 10009 9450 10010
rect 9422 9983 9423 10009
rect 9423 9983 9449 10009
rect 9449 9983 9450 10009
rect 9422 9982 9450 9983
rect 9254 9561 9282 9562
rect 9254 9535 9255 9561
rect 9255 9535 9281 9561
rect 9281 9535 9282 9561
rect 9254 9534 9282 9535
rect 9142 9142 9170 9170
rect 8414 8414 8442 8442
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 8190 7265 8218 7266
rect 8190 7239 8191 7265
rect 8191 7239 8217 7265
rect 8217 7239 8218 7265
rect 8190 7238 8218 7239
rect 8526 7574 8554 7602
rect 8414 7238 8442 7266
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 9478 9505 9506 9506
rect 9478 9479 9479 9505
rect 9479 9479 9505 9505
rect 9505 9479 9506 9505
rect 9478 9478 9506 9479
rect 9926 10542 9954 10570
rect 10094 10262 10122 10290
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9814 10094 9842 10122
rect 9758 9617 9786 9618
rect 9758 9591 9759 9617
rect 9759 9591 9785 9617
rect 9785 9591 9786 9617
rect 9758 9590 9786 9591
rect 9870 9758 9898 9786
rect 10038 9617 10066 9618
rect 10038 9591 10039 9617
rect 10039 9591 10065 9617
rect 10065 9591 10066 9617
rect 10038 9590 10066 9591
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 10094 9422 10122 9450
rect 9534 9198 9562 9226
rect 9534 9086 9562 9114
rect 9534 8889 9562 8890
rect 9534 8863 9535 8889
rect 9535 8863 9561 8889
rect 9561 8863 9562 8889
rect 9534 8862 9562 8863
rect 9366 8777 9394 8778
rect 9366 8751 9367 8777
rect 9367 8751 9393 8777
rect 9393 8751 9394 8777
rect 9366 8750 9394 8751
rect 9422 8470 9450 8498
rect 9870 9142 9898 9170
rect 9926 9198 9954 9226
rect 9646 8945 9674 8946
rect 9646 8919 9647 8945
rect 9647 8919 9673 8945
rect 9673 8919 9674 8945
rect 9646 8918 9674 8919
rect 10038 8918 10066 8946
rect 10206 10486 10234 10514
rect 10206 10094 10234 10122
rect 10262 9702 10290 9730
rect 11774 12614 11802 12642
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 20118 18185 20146 18186
rect 20118 18159 20119 18185
rect 20119 18159 20145 18185
rect 20145 18159 20146 18185
rect 20118 18158 20146 18159
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 12502 13593 12530 13594
rect 12502 13567 12503 13593
rect 12503 13567 12529 13593
rect 12529 13567 12530 13593
rect 12502 13566 12530 13567
rect 13902 13537 13930 13538
rect 13902 13511 13903 13537
rect 13903 13511 13929 13537
rect 13929 13511 13930 13537
rect 13902 13510 13930 13511
rect 14350 13510 14378 13538
rect 12558 13454 12586 13482
rect 12166 13257 12194 13258
rect 12166 13231 12167 13257
rect 12167 13231 12193 13257
rect 12193 13231 12194 13257
rect 12166 13230 12194 13231
rect 12334 12697 12362 12698
rect 12334 12671 12335 12697
rect 12335 12671 12361 12697
rect 12361 12671 12362 12697
rect 12334 12670 12362 12671
rect 12222 12558 12250 12586
rect 13846 13481 13874 13482
rect 13846 13455 13847 13481
rect 13847 13455 13873 13481
rect 13873 13455 13874 13481
rect 13846 13454 13874 13455
rect 12894 13145 12922 13146
rect 12894 13119 12895 13145
rect 12895 13119 12921 13145
rect 12921 13119 12922 13145
rect 12894 13118 12922 13119
rect 12614 13062 12642 13090
rect 12446 12446 12474 12474
rect 13286 13089 13314 13090
rect 13286 13063 13287 13089
rect 13287 13063 13313 13089
rect 13313 13063 13314 13089
rect 13286 13062 13314 13063
rect 18830 13537 18858 13538
rect 18830 13511 18831 13537
rect 18831 13511 18857 13537
rect 18857 13511 18858 13537
rect 18830 13510 18858 13511
rect 14574 13145 14602 13146
rect 14574 13119 14575 13145
rect 14575 13119 14601 13145
rect 14601 13119 14602 13145
rect 14574 13118 14602 13119
rect 14294 12809 14322 12810
rect 14294 12783 14295 12809
rect 14295 12783 14321 12809
rect 14321 12783 14322 12809
rect 14294 12782 14322 12783
rect 12726 12558 12754 12586
rect 13062 12558 13090 12586
rect 13006 12446 13034 12474
rect 12502 12334 12530 12362
rect 11494 11969 11522 11970
rect 11494 11943 11495 11969
rect 11495 11943 11521 11969
rect 11521 11943 11522 11969
rect 11494 11942 11522 11943
rect 12670 12278 12698 12306
rect 12950 12278 12978 12306
rect 11158 11633 11186 11634
rect 11158 11607 11159 11633
rect 11159 11607 11185 11633
rect 11185 11607 11186 11633
rect 11158 11606 11186 11607
rect 11326 11577 11354 11578
rect 11326 11551 11327 11577
rect 11327 11551 11353 11577
rect 11353 11551 11354 11577
rect 11326 11550 11354 11551
rect 11326 11465 11354 11466
rect 11326 11439 11327 11465
rect 11327 11439 11353 11465
rect 11353 11439 11354 11465
rect 11326 11438 11354 11439
rect 10710 11073 10738 11074
rect 10710 11047 10711 11073
rect 10711 11047 10737 11073
rect 10737 11047 10738 11073
rect 10710 11046 10738 11047
rect 10654 10990 10682 11018
rect 10934 10990 10962 11018
rect 10822 10430 10850 10458
rect 10598 9646 10626 9674
rect 10206 9590 10234 9618
rect 9534 8358 9562 8386
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 9926 8526 9954 8554
rect 9534 8022 9562 8050
rect 9870 8049 9898 8050
rect 9870 8023 9871 8049
rect 9871 8023 9897 8049
rect 9897 8023 9898 8049
rect 9870 8022 9898 8023
rect 9310 7966 9338 7994
rect 9590 7966 9618 7994
rect 9590 7601 9618 7602
rect 9590 7575 9591 7601
rect 9591 7575 9617 7601
rect 9617 7575 9618 7601
rect 9590 7574 9618 7575
rect 10990 10374 11018 10402
rect 12054 11689 12082 11690
rect 12054 11663 12055 11689
rect 12055 11663 12081 11689
rect 12081 11663 12082 11689
rect 12054 11662 12082 11663
rect 11662 11550 11690 11578
rect 11886 11577 11914 11578
rect 11886 11551 11887 11577
rect 11887 11551 11913 11577
rect 11913 11551 11914 11577
rect 11886 11550 11914 11551
rect 11326 11046 11354 11074
rect 11550 11102 11578 11130
rect 11830 11046 11858 11074
rect 11662 10710 11690 10738
rect 10934 10345 10962 10346
rect 10934 10319 10935 10345
rect 10935 10319 10961 10345
rect 10961 10319 10962 10345
rect 10934 10318 10962 10319
rect 10934 9561 10962 9562
rect 10934 9535 10935 9561
rect 10935 9535 10961 9561
rect 10961 9535 10962 9561
rect 10934 9534 10962 9535
rect 10990 9198 11018 9226
rect 10822 9142 10850 9170
rect 10710 9086 10738 9114
rect 11158 9534 11186 9562
rect 11158 9310 11186 9338
rect 11326 9281 11354 9282
rect 11326 9255 11327 9281
rect 11327 9255 11353 9281
rect 11353 9255 11354 9281
rect 11326 9254 11354 9255
rect 10374 8750 10402 8778
rect 10430 8414 10458 8442
rect 10934 8414 10962 8442
rect 9982 8358 10010 8386
rect 10206 8385 10234 8386
rect 10206 8359 10207 8385
rect 10207 8359 10233 8385
rect 10233 8359 10234 8385
rect 10206 8358 10234 8359
rect 9982 7993 10010 7994
rect 9982 7967 9983 7993
rect 9983 7967 10009 7993
rect 10009 7967 10010 7993
rect 9982 7966 10010 7967
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 9814 7657 9842 7658
rect 9814 7631 9815 7657
rect 9815 7631 9841 7657
rect 9841 7631 9842 7657
rect 9814 7630 9842 7631
rect 10206 7630 10234 7658
rect 10374 7630 10402 7658
rect 8974 7238 9002 7266
rect 10766 7657 10794 7658
rect 10766 7631 10767 7657
rect 10767 7631 10793 7657
rect 10793 7631 10794 7657
rect 10766 7630 10794 7631
rect 10654 7601 10682 7602
rect 10654 7575 10655 7601
rect 10655 7575 10681 7601
rect 10681 7575 10682 7601
rect 10654 7574 10682 7575
rect 9758 6958 9786 6986
rect 8974 6510 9002 6538
rect 9366 6790 9394 6818
rect 9646 6678 9674 6706
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 8750 2030 8778 2058
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9366 2057 9394 2058
rect 9366 2031 9367 2057
rect 9367 2031 9393 2057
rect 9393 2031 9394 2057
rect 9366 2030 9394 2031
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 9982 6985 10010 6986
rect 9982 6959 9983 6985
rect 9983 6959 10009 6985
rect 10009 6959 10010 6985
rect 9982 6958 10010 6959
rect 10038 6929 10066 6930
rect 10038 6903 10039 6929
rect 10039 6903 10065 6929
rect 10065 6903 10066 6929
rect 10038 6902 10066 6903
rect 9926 6817 9954 6818
rect 9926 6791 9927 6817
rect 9927 6791 9953 6817
rect 9953 6791 9954 6817
rect 9926 6790 9954 6791
rect 9870 6734 9898 6762
rect 10598 6902 10626 6930
rect 10486 6873 10514 6874
rect 10486 6847 10487 6873
rect 10487 6847 10513 6873
rect 10513 6847 10514 6873
rect 10486 6846 10514 6847
rect 11494 9617 11522 9618
rect 11494 9591 11495 9617
rect 11495 9591 11521 9617
rect 11521 9591 11522 9617
rect 11494 9590 11522 9591
rect 11494 9366 11522 9394
rect 11438 9310 11466 9338
rect 11774 10318 11802 10346
rect 12222 11550 12250 11578
rect 12334 11830 12362 11858
rect 11998 10878 12026 10906
rect 12222 10878 12250 10906
rect 11942 10849 11970 10850
rect 11942 10823 11943 10849
rect 11943 10823 11969 10849
rect 11969 10823 11970 10849
rect 11942 10822 11970 10823
rect 11998 10793 12026 10794
rect 11998 10767 11999 10793
rect 11999 10767 12025 10793
rect 12025 10767 12026 10793
rect 11998 10766 12026 10767
rect 11886 10094 11914 10122
rect 12110 10710 12138 10738
rect 12166 10038 12194 10066
rect 12110 9729 12138 9730
rect 12110 9703 12111 9729
rect 12111 9703 12137 9729
rect 12137 9703 12138 9729
rect 12110 9702 12138 9703
rect 12054 9534 12082 9562
rect 11942 9337 11970 9338
rect 11942 9311 11943 9337
rect 11943 9311 11969 9337
rect 11969 9311 11970 9337
rect 11942 9310 11970 9311
rect 11662 9254 11690 9282
rect 11662 9169 11690 9170
rect 11662 9143 11663 9169
rect 11663 9143 11689 9169
rect 11689 9143 11690 9169
rect 11662 9142 11690 9143
rect 11494 8889 11522 8890
rect 11494 8863 11495 8889
rect 11495 8863 11521 8889
rect 11521 8863 11522 8889
rect 11494 8862 11522 8863
rect 11606 8526 11634 8554
rect 11494 8414 11522 8442
rect 12614 11662 12642 11690
rect 13062 12361 13090 12362
rect 13062 12335 13063 12361
rect 13063 12335 13089 12361
rect 13089 12335 13090 12361
rect 13062 12334 13090 12335
rect 13174 12473 13202 12474
rect 13174 12447 13175 12473
rect 13175 12447 13201 12473
rect 13201 12447 13202 12473
rect 13174 12446 13202 12447
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 20006 13118 20034 13146
rect 18830 12782 18858 12810
rect 20006 12782 20034 12810
rect 13286 12361 13314 12362
rect 13286 12335 13287 12361
rect 13287 12335 13313 12361
rect 13313 12335 13314 12361
rect 13286 12334 13314 12335
rect 14014 12361 14042 12362
rect 14014 12335 14015 12361
rect 14015 12335 14041 12361
rect 14041 12335 14042 12361
rect 14014 12334 14042 12335
rect 13398 12278 13426 12306
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 12726 11046 12754 11074
rect 12614 10065 12642 10066
rect 12614 10039 12615 10065
rect 12615 10039 12641 10065
rect 12641 10039 12642 10065
rect 12614 10038 12642 10039
rect 13230 11158 13258 11186
rect 13118 10990 13146 11018
rect 12894 10793 12922 10794
rect 12894 10767 12895 10793
rect 12895 10767 12921 10793
rect 12921 10767 12922 10793
rect 12894 10766 12922 10767
rect 13286 11129 13314 11130
rect 13286 11103 13287 11129
rect 13287 11103 13313 11129
rect 13313 11103 13314 11129
rect 13286 11102 13314 11103
rect 13062 10737 13090 10738
rect 13062 10711 13063 10737
rect 13063 10711 13089 10737
rect 13089 10711 13090 10737
rect 13062 10710 13090 10711
rect 13510 11158 13538 11186
rect 13622 11185 13650 11186
rect 13622 11159 13623 11185
rect 13623 11159 13649 11185
rect 13649 11159 13650 11185
rect 13622 11158 13650 11159
rect 13454 11046 13482 11074
rect 14014 11046 14042 11074
rect 13790 10737 13818 10738
rect 13790 10711 13791 10737
rect 13791 10711 13817 10737
rect 13817 10711 13818 10737
rect 13790 10710 13818 10711
rect 13510 10486 13538 10514
rect 14574 10990 14602 11018
rect 14630 10934 14658 10962
rect 14574 10513 14602 10514
rect 14574 10487 14575 10513
rect 14575 10487 14601 10513
rect 14601 10487 14602 10513
rect 14574 10486 14602 10487
rect 14630 10345 14658 10346
rect 14630 10319 14631 10345
rect 14631 10319 14657 10345
rect 14657 10319 14658 10345
rect 14630 10318 14658 10319
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 14854 10934 14882 10962
rect 20006 11102 20034 11130
rect 18830 10934 18858 10962
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 14854 10318 14882 10346
rect 20006 10766 20034 10794
rect 18830 10318 18858 10346
rect 12334 9702 12362 9730
rect 12726 9702 12754 9730
rect 12670 9561 12698 9562
rect 12670 9535 12671 9561
rect 12671 9535 12697 9561
rect 12697 9535 12698 9561
rect 12670 9534 12698 9535
rect 12502 9422 12530 9450
rect 12894 10009 12922 10010
rect 12894 9983 12895 10009
rect 12895 9983 12921 10009
rect 12921 9983 12922 10009
rect 12894 9982 12922 9983
rect 13230 10009 13258 10010
rect 13230 9983 13231 10009
rect 13231 9983 13257 10009
rect 13257 9983 13258 10009
rect 13230 9982 13258 9983
rect 12894 9897 12922 9898
rect 12894 9871 12895 9897
rect 12895 9871 12921 9897
rect 12921 9871 12922 9897
rect 12894 9870 12922 9871
rect 12950 9478 12978 9506
rect 12782 9281 12810 9282
rect 12782 9255 12783 9281
rect 12783 9255 12809 9281
rect 12809 9255 12810 9281
rect 12782 9254 12810 9255
rect 11046 8358 11074 8386
rect 11494 8302 11522 8330
rect 11382 7630 11410 7658
rect 12334 8553 12362 8554
rect 12334 8527 12335 8553
rect 12335 8527 12361 8553
rect 12361 8527 12362 8553
rect 12334 8526 12362 8527
rect 13510 9870 13538 9898
rect 13174 9646 13202 9674
rect 13342 9505 13370 9506
rect 13342 9479 13343 9505
rect 13343 9479 13369 9505
rect 13369 9479 13370 9505
rect 13342 9478 13370 9479
rect 13454 9478 13482 9506
rect 13006 9310 13034 9338
rect 13286 9366 13314 9394
rect 13342 9198 13370 9226
rect 13790 9590 13818 9618
rect 13734 9561 13762 9562
rect 13734 9535 13735 9561
rect 13735 9535 13761 9561
rect 13761 9535 13762 9561
rect 13734 9534 13762 9535
rect 13622 9505 13650 9506
rect 13622 9479 13623 9505
rect 13623 9479 13649 9505
rect 13649 9479 13650 9505
rect 13622 9478 13650 9479
rect 13734 9422 13762 9450
rect 13790 9505 13818 9506
rect 13790 9479 13791 9505
rect 13791 9479 13817 9505
rect 13817 9479 13818 9505
rect 13790 9478 13818 9479
rect 12950 8833 12978 8834
rect 12950 8807 12951 8833
rect 12951 8807 12977 8833
rect 12977 8807 12978 8833
rect 12950 8806 12978 8807
rect 13118 9169 13146 9170
rect 13118 9143 13119 9169
rect 13119 9143 13145 9169
rect 13145 9143 13146 9169
rect 13118 9142 13146 9143
rect 12670 8441 12698 8442
rect 12670 8415 12671 8441
rect 12671 8415 12697 8441
rect 12697 8415 12698 8441
rect 12670 8414 12698 8415
rect 12222 8302 12250 8330
rect 12334 7937 12362 7938
rect 12334 7911 12335 7937
rect 12335 7911 12361 7937
rect 12361 7911 12362 7937
rect 12334 7910 12362 7911
rect 10822 6790 10850 6818
rect 11494 6846 11522 6874
rect 12110 6846 12138 6874
rect 10934 6734 10962 6762
rect 11606 6790 11634 6818
rect 10094 6510 10122 6538
rect 10374 6678 10402 6706
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 10710 6537 10738 6538
rect 10710 6511 10711 6537
rect 10711 6511 10737 6537
rect 10737 6511 10738 6537
rect 10710 6510 10738 6511
rect 11942 6817 11970 6818
rect 11942 6791 11943 6817
rect 11943 6791 11969 6817
rect 11969 6791 11970 6817
rect 11942 6790 11970 6791
rect 12166 6790 12194 6818
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 10430 2030 10458 2058
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 11046 2057 11074 2058
rect 11046 2031 11047 2057
rect 11047 2031 11073 2057
rect 11073 2031 11074 2057
rect 11046 2030 11074 2031
rect 11438 1806 11466 1834
rect 11830 2590 11858 2618
rect 13566 9142 13594 9170
rect 14182 9926 14210 9954
rect 13958 9590 13986 9618
rect 13902 9422 13930 9450
rect 13734 8833 13762 8834
rect 13734 8807 13735 8833
rect 13735 8807 13761 8833
rect 13761 8807 13762 8833
rect 13734 8806 13762 8807
rect 15022 9953 15050 9954
rect 15022 9927 15023 9953
rect 15023 9927 15049 9953
rect 15049 9927 15050 9953
rect 15022 9926 15050 9927
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 14014 9254 14042 9282
rect 14238 9478 14266 9506
rect 15022 9198 15050 9226
rect 15246 9225 15274 9226
rect 15246 9199 15247 9225
rect 15247 9199 15273 9225
rect 15273 9199 15274 9225
rect 15246 9198 15274 9199
rect 15358 9142 15386 9170
rect 18830 9814 18858 9842
rect 20006 9758 20034 9786
rect 20006 9422 20034 9450
rect 18942 9198 18970 9226
rect 18774 9142 18802 9170
rect 20006 9113 20034 9114
rect 20006 9087 20007 9113
rect 20007 9087 20033 9113
rect 20033 9087 20034 9113
rect 20006 9086 20034 9087
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 14126 8806 14154 8834
rect 13118 8414 13146 8442
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 14126 8526 14154 8554
rect 14294 8441 14322 8442
rect 14294 8415 14295 8441
rect 14295 8415 14321 8441
rect 14321 8415 14322 8441
rect 14294 8414 14322 8415
rect 20006 8414 20034 8442
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 12670 6846 12698 6874
rect 12950 7910 12978 7938
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 13174 6846 13202 6874
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 12390 2617 12418 2618
rect 12390 2591 12391 2617
rect 12391 2591 12417 2617
rect 12417 2591 12418 2617
rect 12390 2590 12418 2591
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 12446 2030 12474 2058
rect 13118 2057 13146 2058
rect 13118 2031 13119 2057
rect 13119 2031 13145 2057
rect 13145 2031 13146 2057
rect 13118 2030 13146 2031
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 8409 19110 8414 19138
rect 8442 19110 9030 19138
rect 9058 19110 9063 19138
rect 10425 19110 10430 19138
rect 10458 19110 11046 19138
rect 11074 19110 11079 19138
rect 11769 19110 11774 19138
rect 11802 19110 12782 19138
rect 12810 19110 12815 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 8073 18718 8078 18746
rect 8106 18718 9198 18746
rect 9226 18718 9231 18746
rect 10089 18718 10094 18746
rect 10122 18718 10710 18746
rect 10738 18718 10743 18746
rect 12441 18718 12446 18746
rect 12474 18718 13118 18746
rect 13146 18718 13151 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 20600 18186 21000 18200
rect 20113 18158 20118 18186
rect 20146 18158 21000 18186
rect 20600 18144 21000 18158
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 8801 13846 8806 13874
rect 8834 13846 9086 13874
rect 9114 13846 10710 13874
rect 10738 13846 10743 13874
rect 7401 13790 7406 13818
rect 7434 13790 8022 13818
rect 8050 13790 8055 13818
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 9417 13622 9422 13650
rect 9450 13622 10318 13650
rect 10346 13622 10351 13650
rect 11937 13566 11942 13594
rect 11970 13566 12502 13594
rect 12530 13566 12535 13594
rect 13897 13510 13902 13538
rect 13930 13510 14350 13538
rect 14378 13510 18830 13538
rect 18858 13510 18863 13538
rect 0 13482 400 13496
rect 0 13454 2086 13482
rect 2114 13454 2119 13482
rect 10089 13454 10094 13482
rect 10122 13454 10262 13482
rect 10290 13454 10295 13482
rect 12553 13454 12558 13482
rect 12586 13454 13846 13482
rect 13874 13454 13879 13482
rect 0 13440 400 13454
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 8353 13286 8358 13314
rect 8386 13286 8806 13314
rect 8834 13286 9254 13314
rect 9282 13286 9814 13314
rect 9842 13286 9847 13314
rect 9025 13230 9030 13258
rect 9058 13230 9534 13258
rect 9562 13230 9567 13258
rect 9921 13230 9926 13258
rect 9954 13230 10486 13258
rect 10514 13230 10519 13258
rect 11433 13230 11438 13258
rect 11466 13230 12166 13258
rect 12194 13230 12199 13258
rect 8353 13174 8358 13202
rect 8386 13174 8750 13202
rect 8778 13174 8783 13202
rect 9865 13174 9870 13202
rect 9898 13174 10150 13202
rect 10178 13174 10183 13202
rect 20600 13146 21000 13160
rect 9697 13118 9702 13146
rect 9730 13118 10318 13146
rect 10346 13118 10351 13146
rect 12889 13118 12894 13146
rect 12922 13118 14574 13146
rect 14602 13118 14607 13146
rect 20001 13118 20006 13146
rect 20034 13118 21000 13146
rect 20600 13104 21000 13118
rect 7289 13062 7294 13090
rect 7322 13062 7910 13090
rect 7938 13062 7943 13090
rect 12609 13062 12614 13090
rect 12642 13062 13286 13090
rect 13314 13062 13319 13090
rect 8073 13006 8078 13034
rect 8106 13006 8750 13034
rect 8778 13006 8783 13034
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 20600 12810 21000 12824
rect 14289 12782 14294 12810
rect 14322 12782 18830 12810
rect 18858 12782 18863 12810
rect 20001 12782 20006 12810
rect 20034 12782 21000 12810
rect 20600 12768 21000 12782
rect 7737 12670 7742 12698
rect 7770 12670 10878 12698
rect 10906 12670 10911 12698
rect 11153 12670 11158 12698
rect 11186 12670 12334 12698
rect 12362 12670 12367 12698
rect 11209 12614 11214 12642
rect 11242 12614 11774 12642
rect 11802 12614 11807 12642
rect 10593 12558 10598 12586
rect 10626 12558 11046 12586
rect 11074 12558 12222 12586
rect 12250 12558 12726 12586
rect 12754 12558 13062 12586
rect 13090 12558 13095 12586
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 12441 12446 12446 12474
rect 12474 12446 13006 12474
rect 13034 12446 13174 12474
rect 13202 12446 13207 12474
rect 2137 12334 2142 12362
rect 2170 12334 6734 12362
rect 6762 12334 6767 12362
rect 12497 12334 12502 12362
rect 12530 12334 13062 12362
rect 13090 12334 13095 12362
rect 13281 12334 13286 12362
rect 13314 12334 14014 12362
rect 14042 12334 14047 12362
rect 9417 12278 9422 12306
rect 9450 12278 12670 12306
rect 12698 12278 12703 12306
rect 12945 12278 12950 12306
rect 12978 12278 13398 12306
rect 13426 12278 13431 12306
rect 961 12222 966 12250
rect 994 12222 999 12250
rect 0 12138 400 12152
rect 966 12138 994 12222
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 0 12110 994 12138
rect 0 12096 400 12110
rect 9361 12054 9366 12082
rect 9394 12054 9814 12082
rect 9842 12054 9847 12082
rect 6729 11998 6734 12026
rect 6762 11998 7966 12026
rect 7994 11998 7999 12026
rect 10929 11942 10934 11970
rect 10962 11942 11494 11970
rect 11522 11942 11527 11970
rect 7401 11886 7406 11914
rect 7434 11886 7798 11914
rect 7826 11886 7831 11914
rect 10425 11886 10430 11914
rect 10458 11886 11046 11914
rect 11074 11886 11079 11914
rect 8129 11830 8134 11858
rect 8162 11830 8526 11858
rect 8554 11830 8694 11858
rect 8722 11830 9366 11858
rect 9394 11830 9399 11858
rect 10817 11830 10822 11858
rect 10850 11830 10990 11858
rect 11018 11830 12334 11858
rect 12362 11830 12367 11858
rect 7849 11774 7854 11802
rect 7882 11774 8022 11802
rect 8050 11774 8414 11802
rect 8442 11774 8447 11802
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 6449 11662 6454 11690
rect 6482 11662 6734 11690
rect 6762 11662 7070 11690
rect 7098 11662 7574 11690
rect 7602 11662 8134 11690
rect 8162 11662 8167 11690
rect 9081 11662 9086 11690
rect 9114 11662 9422 11690
rect 9450 11662 9455 11690
rect 9683 11662 9702 11690
rect 9730 11662 9735 11690
rect 9809 11662 9814 11690
rect 9842 11662 10934 11690
rect 10962 11662 10967 11690
rect 12049 11662 12054 11690
rect 12082 11662 12614 11690
rect 12642 11662 12647 11690
rect 4186 11606 5278 11634
rect 5306 11606 6958 11634
rect 6986 11606 6991 11634
rect 7546 11606 7910 11634
rect 7938 11606 8918 11634
rect 8946 11606 8951 11634
rect 9590 11606 10206 11634
rect 10234 11606 10239 11634
rect 10313 11606 10318 11634
rect 10346 11606 11158 11634
rect 11186 11606 11191 11634
rect 4186 11578 4214 11606
rect 7546 11578 7574 11606
rect 9590 11578 9618 11606
rect 2137 11550 2142 11578
rect 2170 11550 4214 11578
rect 7009 11550 7014 11578
rect 7042 11550 7294 11578
rect 7322 11550 7574 11578
rect 8185 11550 8190 11578
rect 8218 11550 9590 11578
rect 9618 11550 9623 11578
rect 9977 11550 9982 11578
rect 10010 11550 10374 11578
rect 10402 11550 10766 11578
rect 10794 11550 10799 11578
rect 10873 11550 10878 11578
rect 10906 11550 11326 11578
rect 11354 11550 11662 11578
rect 11690 11550 11695 11578
rect 11881 11550 11886 11578
rect 11914 11550 12222 11578
rect 12250 11550 12255 11578
rect 6337 11494 6342 11522
rect 6370 11494 6790 11522
rect 6818 11494 6823 11522
rect 7345 11494 7350 11522
rect 7378 11494 8022 11522
rect 8050 11494 8055 11522
rect 9417 11494 9422 11522
rect 9450 11494 9870 11522
rect 9898 11494 9903 11522
rect 0 11466 400 11480
rect 0 11438 966 11466
rect 994 11438 999 11466
rect 7681 11438 7686 11466
rect 7714 11438 8078 11466
rect 8106 11438 11326 11466
rect 11354 11438 11359 11466
rect 0 11424 400 11438
rect 9753 11382 9758 11410
rect 9786 11382 10094 11410
rect 10122 11382 10127 11410
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 9529 11270 9534 11298
rect 9562 11270 9814 11298
rect 9842 11270 10654 11298
rect 10682 11270 10687 11298
rect 961 11214 966 11242
rect 994 11214 999 11242
rect 9977 11214 9982 11242
rect 10010 11214 10150 11242
rect 10178 11214 10183 11242
rect 0 11130 400 11144
rect 966 11130 994 11214
rect 2137 11158 2142 11186
rect 2170 11158 4214 11186
rect 13225 11158 13230 11186
rect 13258 11158 13510 11186
rect 13538 11158 13622 11186
rect 13650 11158 13655 11186
rect 0 11102 994 11130
rect 4186 11130 4214 11158
rect 20600 11130 21000 11144
rect 4186 11102 4998 11130
rect 5026 11102 7238 11130
rect 7266 11102 7271 11130
rect 9641 11102 9646 11130
rect 9674 11102 9926 11130
rect 9954 11102 9959 11130
rect 11545 11102 11550 11130
rect 11578 11102 13286 11130
rect 13314 11102 13319 11130
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 0 11088 400 11102
rect 20600 11088 21000 11102
rect 9137 11046 9142 11074
rect 9170 11046 9814 11074
rect 9842 11046 10710 11074
rect 10738 11046 10743 11074
rect 11321 11046 11326 11074
rect 11354 11046 11830 11074
rect 11858 11046 11863 11074
rect 12721 11046 12726 11074
rect 12754 11046 13454 11074
rect 13482 11046 14014 11074
rect 14042 11046 14047 11074
rect 10649 10990 10654 11018
rect 10682 10990 10934 11018
rect 10962 10990 10967 11018
rect 13113 10990 13118 11018
rect 13146 10990 14574 11018
rect 14602 10990 14607 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 14625 10934 14630 10962
rect 14658 10934 14854 10962
rect 14882 10934 18830 10962
rect 18858 10934 18863 10962
rect 6561 10878 6566 10906
rect 6594 10878 7238 10906
rect 7266 10878 7406 10906
rect 7434 10878 7854 10906
rect 7882 10878 7887 10906
rect 8801 10878 8806 10906
rect 8834 10878 11998 10906
rect 12026 10878 12222 10906
rect 12250 10878 12255 10906
rect 6785 10822 6790 10850
rect 6818 10822 7126 10850
rect 7154 10822 11942 10850
rect 11970 10822 11975 10850
rect 20600 10794 21000 10808
rect 5385 10766 5390 10794
rect 5418 10766 6734 10794
rect 6762 10766 7182 10794
rect 7210 10766 7798 10794
rect 7826 10766 7831 10794
rect 8017 10766 8022 10794
rect 8050 10766 9030 10794
rect 9058 10766 10094 10794
rect 10122 10766 10127 10794
rect 11993 10766 11998 10794
rect 12026 10766 12894 10794
rect 12922 10766 12927 10794
rect 20001 10766 20006 10794
rect 20034 10766 21000 10794
rect 20600 10752 21000 10766
rect 11657 10710 11662 10738
rect 11690 10710 12110 10738
rect 12138 10710 12143 10738
rect 13057 10710 13062 10738
rect 13090 10710 13790 10738
rect 13818 10710 13823 10738
rect 6449 10654 6454 10682
rect 6482 10654 6734 10682
rect 6762 10654 8974 10682
rect 9002 10654 9007 10682
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 9921 10542 9926 10570
rect 9954 10542 10094 10570
rect 10122 10542 10127 10570
rect 9641 10486 9646 10514
rect 9674 10486 10206 10514
rect 10234 10486 10239 10514
rect 13505 10486 13510 10514
rect 13538 10486 14574 10514
rect 14602 10486 14607 10514
rect 7569 10430 7574 10458
rect 7602 10430 8470 10458
rect 8498 10430 10822 10458
rect 10850 10430 10855 10458
rect 8129 10374 8134 10402
rect 8162 10374 8638 10402
rect 8666 10374 8862 10402
rect 8890 10374 10990 10402
rect 11018 10374 11023 10402
rect 7737 10318 7742 10346
rect 7770 10318 8190 10346
rect 8218 10318 8526 10346
rect 8554 10318 10934 10346
rect 10962 10318 11774 10346
rect 11802 10318 11807 10346
rect 14625 10318 14630 10346
rect 14658 10318 14854 10346
rect 14882 10318 18830 10346
rect 18858 10318 18863 10346
rect 9193 10262 9198 10290
rect 9226 10262 9478 10290
rect 9506 10262 10094 10290
rect 10122 10262 10127 10290
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 9809 10094 9814 10122
rect 9842 10094 10206 10122
rect 10234 10094 11886 10122
rect 11914 10094 11919 10122
rect 9305 10038 9310 10066
rect 9338 10038 12082 10066
rect 12161 10038 12166 10066
rect 12194 10038 12614 10066
rect 12642 10038 12647 10066
rect 12054 10010 12082 10038
rect 6449 9982 6454 10010
rect 6482 9982 7126 10010
rect 7154 9982 7462 10010
rect 7490 9982 7495 10010
rect 7546 9982 8806 10010
rect 8834 9982 9422 10010
rect 9450 9982 9455 10010
rect 12054 9982 12894 10010
rect 12922 9982 13230 10010
rect 13258 9982 13263 10010
rect 7546 9954 7574 9982
rect 2081 9926 2086 9954
rect 2114 9926 7574 9954
rect 14177 9926 14182 9954
rect 14210 9926 15022 9954
rect 15050 9926 18858 9954
rect 12889 9870 12894 9898
rect 12922 9870 13510 9898
rect 13538 9870 13543 9898
rect 18830 9842 18858 9926
rect 18825 9814 18830 9842
rect 18858 9814 18863 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 20600 9786 21000 9800
rect 7905 9758 7910 9786
rect 7938 9758 8078 9786
rect 8106 9758 9870 9786
rect 9898 9758 9903 9786
rect 20001 9758 20006 9786
rect 20034 9758 21000 9786
rect 20600 9744 21000 9758
rect 6729 9702 6734 9730
rect 6762 9702 10262 9730
rect 10290 9702 10295 9730
rect 12105 9702 12110 9730
rect 12138 9702 12334 9730
rect 12362 9702 12726 9730
rect 12754 9702 12759 9730
rect 10593 9646 10598 9674
rect 10626 9646 13174 9674
rect 13202 9646 13207 9674
rect 7401 9590 7406 9618
rect 7434 9590 7910 9618
rect 7938 9590 7943 9618
rect 9753 9590 9758 9618
rect 9786 9590 10038 9618
rect 10066 9590 10206 9618
rect 10234 9590 11494 9618
rect 11522 9590 11527 9618
rect 13785 9590 13790 9618
rect 13818 9590 13958 9618
rect 13986 9590 13991 9618
rect 7233 9534 7238 9562
rect 7266 9534 7518 9562
rect 7546 9534 8190 9562
rect 8218 9534 8223 9562
rect 9249 9534 9254 9562
rect 9282 9534 10934 9562
rect 10962 9534 11158 9562
rect 11186 9534 11191 9562
rect 12049 9534 12054 9562
rect 12082 9534 12670 9562
rect 12698 9534 13734 9562
rect 13762 9534 13767 9562
rect 8353 9478 8358 9506
rect 8386 9478 9478 9506
rect 9506 9478 9511 9506
rect 12945 9478 12950 9506
rect 12978 9478 13342 9506
rect 13370 9478 13375 9506
rect 13449 9478 13454 9506
rect 13482 9478 13622 9506
rect 13650 9478 13655 9506
rect 13785 9478 13790 9506
rect 13818 9478 14238 9506
rect 14266 9478 14271 9506
rect 20600 9450 21000 9464
rect 10089 9422 10094 9450
rect 10122 9422 12502 9450
rect 12530 9422 12535 9450
rect 13729 9422 13734 9450
rect 13762 9422 13902 9450
rect 13930 9422 13935 9450
rect 20001 9422 20006 9450
rect 20034 9422 21000 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 20600 9408 21000 9422
rect 11489 9366 11494 9394
rect 11522 9366 13286 9394
rect 13314 9366 13454 9394
rect 11153 9310 11158 9338
rect 11186 9310 11438 9338
rect 11466 9310 11471 9338
rect 11937 9310 11942 9338
rect 11970 9310 13006 9338
rect 13034 9310 13039 9338
rect 13426 9282 13454 9366
rect 5049 9254 5054 9282
rect 5082 9254 5278 9282
rect 5306 9254 6566 9282
rect 6594 9254 6902 9282
rect 6930 9254 6935 9282
rect 11321 9254 11326 9282
rect 11354 9254 11662 9282
rect 11690 9254 12782 9282
rect 12810 9254 12815 9282
rect 13426 9254 14014 9282
rect 14042 9254 14047 9282
rect 6673 9198 6678 9226
rect 6706 9198 7126 9226
rect 7154 9198 7406 9226
rect 7434 9198 7439 9226
rect 9529 9198 9534 9226
rect 9562 9198 9926 9226
rect 9954 9198 10990 9226
rect 11018 9198 11023 9226
rect 13337 9198 13342 9226
rect 13370 9198 15022 9226
rect 15050 9198 15246 9226
rect 15274 9198 18942 9226
rect 18970 9198 18975 9226
rect 5609 9142 5614 9170
rect 5642 9142 6734 9170
rect 6762 9142 6767 9170
rect 9137 9142 9142 9170
rect 9170 9142 9870 9170
rect 9898 9142 9903 9170
rect 10817 9142 10822 9170
rect 10850 9142 11662 9170
rect 11690 9142 11695 9170
rect 13113 9142 13118 9170
rect 13146 9142 13566 9170
rect 13594 9142 13599 9170
rect 15353 9142 15358 9170
rect 15386 9142 18774 9170
rect 18802 9142 18807 9170
rect 20600 9114 21000 9128
rect 9529 9086 9534 9114
rect 9562 9086 10094 9114
rect 10122 9086 10710 9114
rect 10738 9086 10743 9114
rect 20001 9086 20006 9114
rect 20034 9086 21000 9114
rect 20600 9072 21000 9086
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 9641 8918 9646 8946
rect 9674 8918 10038 8946
rect 10066 8918 10071 8946
rect 9529 8862 9534 8890
rect 9562 8862 11494 8890
rect 11522 8862 11527 8890
rect 12945 8806 12950 8834
rect 12978 8806 13734 8834
rect 13762 8806 13767 8834
rect 14121 8806 14126 8834
rect 14154 8806 18830 8834
rect 18858 8806 18863 8834
rect 9361 8750 9366 8778
rect 9394 8750 10374 8778
rect 10402 8750 10407 8778
rect 7233 8694 7238 8722
rect 7266 8694 7854 8722
rect 7882 8694 7887 8722
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 7793 8526 7798 8554
rect 7826 8526 8190 8554
rect 8218 8526 9926 8554
rect 9954 8526 11606 8554
rect 11634 8526 11639 8554
rect 12329 8526 12334 8554
rect 12362 8526 14126 8554
rect 14154 8526 14159 8554
rect 7681 8470 7686 8498
rect 7714 8470 9422 8498
rect 9450 8470 9455 8498
rect 20600 8442 21000 8456
rect 6897 8414 6902 8442
rect 6930 8414 7350 8442
rect 7378 8414 8414 8442
rect 8442 8414 8447 8442
rect 10425 8414 10430 8442
rect 10458 8414 10934 8442
rect 10962 8414 11494 8442
rect 11522 8414 11527 8442
rect 12665 8414 12670 8442
rect 12698 8414 13118 8442
rect 13146 8414 14294 8442
rect 14322 8414 14327 8442
rect 20001 8414 20006 8442
rect 20034 8414 21000 8442
rect 20600 8400 21000 8414
rect 8353 8358 8358 8386
rect 8386 8358 9534 8386
rect 9562 8358 9567 8386
rect 9977 8358 9982 8386
rect 10010 8358 10206 8386
rect 10234 8358 11046 8386
rect 11074 8358 11079 8386
rect 11489 8302 11494 8330
rect 11522 8302 12222 8330
rect 12250 8302 12255 8330
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 9529 8022 9534 8050
rect 9562 8022 9870 8050
rect 9898 8022 9903 8050
rect 9305 7966 9310 7994
rect 9338 7966 9590 7994
rect 9618 7966 9982 7994
rect 10010 7966 10015 7994
rect 12329 7910 12334 7938
rect 12362 7910 12950 7938
rect 12978 7910 12983 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 9809 7630 9814 7658
rect 9842 7630 10206 7658
rect 10234 7630 10239 7658
rect 10369 7630 10374 7658
rect 10402 7630 10766 7658
rect 10794 7630 11382 7658
rect 11410 7630 11415 7658
rect 10206 7602 10234 7630
rect 8521 7574 8526 7602
rect 8554 7574 9590 7602
rect 9618 7574 9623 7602
rect 10206 7574 10654 7602
rect 10682 7574 10687 7602
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 8185 7238 8190 7266
rect 8218 7238 8414 7266
rect 8442 7238 8974 7266
rect 9002 7238 9007 7266
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 9753 6958 9758 6986
rect 9786 6958 9982 6986
rect 10010 6958 10015 6986
rect 9697 6902 9702 6930
rect 9730 6902 10038 6930
rect 10066 6902 10598 6930
rect 10626 6902 10631 6930
rect 10481 6846 10486 6874
rect 10514 6846 11494 6874
rect 11522 6846 12110 6874
rect 12138 6846 12670 6874
rect 12698 6846 13174 6874
rect 13202 6846 13207 6874
rect 9361 6790 9366 6818
rect 9394 6790 9926 6818
rect 9954 6790 9959 6818
rect 10817 6790 10822 6818
rect 10850 6790 11606 6818
rect 11634 6790 11942 6818
rect 11970 6790 12166 6818
rect 12194 6790 12199 6818
rect 9865 6734 9870 6762
rect 9898 6734 10934 6762
rect 10962 6734 10967 6762
rect 9641 6678 9646 6706
rect 9674 6678 10374 6706
rect 10402 6678 10407 6706
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 8969 6510 8974 6538
rect 9002 6510 10094 6538
rect 10122 6510 10710 6538
rect 10738 6510 10743 6538
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 11825 2590 11830 2618
rect 11858 2590 12390 2618
rect 12418 2590 12423 2618
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 8745 2030 8750 2058
rect 8778 2030 9366 2058
rect 9394 2030 9399 2058
rect 10425 2030 10430 2058
rect 10458 2030 11046 2058
rect 11074 2030 11079 2058
rect 12441 2030 12446 2058
rect 12474 2030 13118 2058
rect 13146 2030 13151 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 11433 1806 11438 1834
rect 11466 1806 12782 1834
rect 12810 1806 12815 1834
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 9702 11662 9730 11690
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 10094 10542 10122 10570
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 10094 9086 10122 9114
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 9702 6902 9730 6930
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 9702 11690 9730 11695
rect 9702 6930 9730 11662
rect 9702 6897 9730 6902
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 10094 10570 10122 10575
rect 10094 9114 10122 10542
rect 10094 9081 10122 9086
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7056 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7840 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1698175906
transform 1 0 12432 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_
timestamp 1698175906
transform 1 0 7336 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9352 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _116_
timestamp 1698175906
transform 1 0 9744 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11368 0 -1 9408
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12712 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform 1 0 9744 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698175906
transform 1 0 10640 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform 1 0 11760 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _122_
timestamp 1698175906
transform 1 0 7000 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8232 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _124_
timestamp 1698175906
transform 1 0 9520 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10360 0 1 10192
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform 1 0 11816 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12040 0 -1 8624
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _128_
timestamp 1698175906
transform 1 0 9408 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11032 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _130_
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _131_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12600 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform 1 0 10080 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _133_
timestamp 1698175906
transform 1 0 7392 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _134_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8400 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _135_
timestamp 1698175906
transform 1 0 10080 0 1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _136_
timestamp 1698175906
transform -1 0 10024 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1698175906
transform -1 0 9520 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform 1 0 9800 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _139_
timestamp 1698175906
transform 1 0 10192 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _140_
timestamp 1698175906
transform -1 0 7952 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _141_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7672 0 1 9408
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _142_
timestamp 1698175906
transform -1 0 7000 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _143_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8512 0 -1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _144_
timestamp 1698175906
transform 1 0 8400 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _145_
timestamp 1698175906
transform -1 0 9632 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _146_
timestamp 1698175906
transform -1 0 9296 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _147_
timestamp 1698175906
transform 1 0 7952 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _148_
timestamp 1698175906
transform -1 0 8008 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _149_
timestamp 1698175906
transform -1 0 7672 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _150_
timestamp 1698175906
transform 1 0 11088 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _151_
timestamp 1698175906
transform 1 0 7616 0 1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _152_
timestamp 1698175906
transform -1 0 8960 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _153_
timestamp 1698175906
transform -1 0 8568 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _154_
timestamp 1698175906
transform -1 0 8904 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _155_
timestamp 1698175906
transform -1 0 8176 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _156_
timestamp 1698175906
transform -1 0 7336 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _157_
timestamp 1698175906
transform -1 0 9408 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _158_
timestamp 1698175906
transform -1 0 9184 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _159_
timestamp 1698175906
transform -1 0 7112 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _160_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _161_
timestamp 1698175906
transform -1 0 7392 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _162_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 6944 0 -1 10976
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _163_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8288 0 -1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _164_
timestamp 1698175906
transform 1 0 7280 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _165_
timestamp 1698175906
transform -1 0 9912 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _166_
timestamp 1698175906
transform -1 0 10472 0 1 8624
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _167_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9464 0 -1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _168_
timestamp 1698175906
transform -1 0 8064 0 -1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _169_
timestamp 1698175906
transform -1 0 8456 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _170_
timestamp 1698175906
transform -1 0 8176 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _171_
timestamp 1698175906
transform 1 0 9408 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _172_
timestamp 1698175906
transform 1 0 10136 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _173_
timestamp 1698175906
transform 1 0 9464 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _174_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9856 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _175_
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _176_
timestamp 1698175906
transform 1 0 10472 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform 1 0 10080 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _178_
timestamp 1698175906
transform -1 0 9800 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _179_
timestamp 1698175906
transform -1 0 11872 0 1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _180_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12432 0 1 9408
box -43 -43 1891 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _181_
timestamp 1698175906
transform 1 0 10024 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _182_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10640 0 1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _183_
timestamp 1698175906
transform 1 0 11312 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _184_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11032 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _185_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10808 0 1 10976
box -43 -43 995 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _186_
timestamp 1698175906
transform 1 0 11312 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _187_
timestamp 1698175906
transform 1 0 12040 0 1 7840
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _188_
timestamp 1698175906
transform -1 0 11984 0 1 7840
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _189_
timestamp 1698175906
transform 1 0 9576 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _190_
timestamp 1698175906
transform 1 0 10136 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _191_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9800 0 -1 7056
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _192_
timestamp 1698175906
transform -1 0 11704 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _193_
timestamp 1698175906
transform 1 0 13944 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _194_
timestamp 1698175906
transform 1 0 13720 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _195_
timestamp 1698175906
transform 1 0 11592 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _196_
timestamp 1698175906
transform -1 0 13104 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _197_
timestamp 1698175906
transform 1 0 11704 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _198_
timestamp 1698175906
transform 1 0 12040 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _199_
timestamp 1698175906
transform 1 0 13216 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _200_
timestamp 1698175906
transform 1 0 9688 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _201_
timestamp 1698175906
transform -1 0 13048 0 -1 10192
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _202_
timestamp 1698175906
transform 1 0 13440 0 1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _203_
timestamp 1698175906
transform -1 0 14000 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _204_
timestamp 1698175906
transform 1 0 12600 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _205_
timestamp 1698175906
transform 1 0 10696 0 1 12544
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _206_
timestamp 1698175906
transform 1 0 12264 0 1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _207_
timestamp 1698175906
transform -1 0 14168 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _208_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12152 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _209_
timestamp 1698175906
transform 1 0 12992 0 -1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _210_
timestamp 1698175906
transform -1 0 14728 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _211_
timestamp 1698175906
transform 1 0 13048 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _212_
timestamp 1698175906
transform 1 0 11760 0 -1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _213_
timestamp 1698175906
transform 1 0 12824 0 -1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _214_
timestamp 1698175906
transform -1 0 14728 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _215_
timestamp 1698175906
transform 1 0 11424 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _216_
timestamp 1698175906
transform 1 0 13216 0 1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _217_
timestamp 1698175906
transform 1 0 9800 0 -1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _218_
timestamp 1698175906
transform 1 0 8792 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _219_
timestamp 1698175906
transform 1 0 9184 0 1 8624
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 8960 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 4928 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 5152 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 6776 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 8008 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 6832 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform -1 0 6832 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform -1 0 6552 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform -1 0 8288 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 8064 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 6944 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _232_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10360 0 -1 7056
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform 1 0 8568 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 10472 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform 1 0 11424 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform 1 0 8848 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 13496 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698175906
transform 1 0 10976 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform 1 0 13496 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _240_
timestamp 1698175906
transform 1 0 12824 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _241_
timestamp 1698175906
transform 1 0 12768 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _242_
timestamp 1698175906
transform 1 0 13328 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _243_
timestamp 1698175906
transform 1 0 13328 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _244_
timestamp 1698175906
transform 1 0 7224 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _247_
timestamp 1698175906
transform 1 0 15120 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _248_
timestamp 1698175906
transform 1 0 12096 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _249_
timestamp 1698175906
transform 1 0 11480 0 1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14280 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 10696 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 6552 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 6888 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 8400 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 9352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 8456 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 7616 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 7504 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 8680 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 10024 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform -1 0 8848 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform -1 0 12208 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 10696 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 12208 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 13160 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform 1 0 10696 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 14000 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform 1 0 12712 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform 1 0 13104 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__CLK
timestamp 1698175906
transform 1 0 14560 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__CLK
timestamp 1698175906
transform 1 0 14616 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__CLK
timestamp 1698175906
transform 1 0 12712 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__CLK
timestamp 1698175906
transform 1 0 13216 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__CLK
timestamp 1698175906
transform 1 0 8960 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 8792 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9352 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 11424 0 -1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 11088 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_144
timestamp 1698175906
transform 1 0 8736 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_171
timestamp 1698175906
transform 1 0 10248 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_201 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11928 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 14000 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 15792 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 16240 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_177 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_193
timestamp 1698175906
transform 1 0 11480 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_197
timestamp 1698175906
transform 1 0 11704 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_225
timestamp 1698175906
transform 1 0 13272 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_139
timestamp 1698175906
transform 1 0 8456 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_143
timestamp 1698175906
transform 1 0 8680 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_145
timestamp 1698175906
transform 1 0 8792 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_181
timestamp 1698175906
transform 1 0 10808 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_189
timestamp 1698175906
transform 1 0 11256 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_199
timestamp 1698175906
transform 1 0 11816 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_203
timestamp 1698175906
transform 1 0 12040 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_206
timestamp 1698175906
transform 1 0 12208 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_238
timestamp 1698175906
transform 1 0 14000 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_242
timestamp 1698175906
transform 1 0 14224 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698175906
transform 1 0 14336 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_158
timestamp 1698175906
transform 1 0 9520 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_123
timestamp 1698175906
transform 1 0 7560 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_131
timestamp 1698175906
transform 1 0 8008 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_165
timestamp 1698175906
transform 1 0 9912 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_185
timestamp 1698175906
transform 1 0 11032 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_189
timestamp 1698175906
transform 1 0 11256 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_191
timestamp 1698175906
transform 1 0 11368 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_221
timestamp 1698175906
transform 1 0 13048 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_225
timestamp 1698175906
transform 1 0 13272 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 14168 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 8288 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_150
timestamp 1698175906
transform 1 0 9072 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_154
timestamp 1698175906
transform 1 0 9296 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_156
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_167
timestamp 1698175906
transform 1 0 10024 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_183
timestamp 1698175906
transform 1 0 10920 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_199
timestamp 1698175906
transform 1 0 11816 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698175906
transform 1 0 12264 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 12376 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 16128 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_115
timestamp 1698175906
transform 1 0 7112 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_146
timestamp 1698175906
transform 1 0 8848 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_150
timestamp 1698175906
transform 1 0 9072 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_158
timestamp 1698175906
transform 1 0 9520 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_168
timestamp 1698175906
transform 1 0 10080 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698175906
transform 1 0 10304 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 10416 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_185
timestamp 1698175906
transform 1 0 11032 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_189
timestamp 1698175906
transform 1 0 11256 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_202
timestamp 1698175906
transform 1 0 11984 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_210
timestamp 1698175906
transform 1 0 12432 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698175906
transform 1 0 14224 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 14336 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_104
timestamp 1698175906
transform 1 0 6496 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_108
timestamp 1698175906
transform 1 0 6720 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698175906
transform 1 0 8400 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_144
timestamp 1698175906
transform 1 0 8736 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_150
timestamp 1698175906
transform 1 0 9072 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_154
timestamp 1698175906
transform 1 0 9296 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_164
timestamp 1698175906
transform 1 0 9856 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_168
timestamp 1698175906
transform 1 0 10080 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_175
timestamp 1698175906
transform 1 0 10472 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_183
timestamp 1698175906
transform 1 0 10920 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_187
timestamp 1698175906
transform 1 0 11144 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_189
timestamp 1698175906
transform 1 0 11256 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_196
timestamp 1698175906
transform 1 0 11648 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_200
timestamp 1698175906
transform 1 0 11872 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_202
timestamp 1698175906
transform 1 0 11984 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_241
timestamp 1698175906
transform 1 0 14168 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_245
timestamp 1698175906
transform 1 0 14392 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698175906
transform 1 0 16184 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 16296 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 20048 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 20160 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_123
timestamp 1698175906
transform 1 0 7560 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_131
timestamp 1698175906
transform 1 0 8008 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_135
timestamp 1698175906
transform 1 0 8232 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_137
timestamp 1698175906
transform 1 0 8344 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_140
timestamp 1698175906
transform 1 0 8512 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_148
timestamp 1698175906
transform 1 0 8960 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_185
timestamp 1698175906
transform 1 0 11032 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_189
timestamp 1698175906
transform 1 0 11256 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_197
timestamp 1698175906
transform 1 0 11704 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_221
timestamp 1698175906
transform 1 0 13048 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_229
timestamp 1698175906
transform 1 0 13496 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698175906
transform 1 0 14168 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_109
timestamp 1698175906
transform 1 0 6776 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_125
timestamp 1698175906
transform 1 0 7672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_162
timestamp 1698175906
transform 1 0 9744 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_172
timestamp 1698175906
transform 1 0 10304 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_176
timestamp 1698175906
transform 1 0 10528 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_191
timestamp 1698175906
transform 1 0 11368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_203
timestamp 1698175906
transform 1 0 12040 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698175906
transform 1 0 12264 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 12376 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_214
timestamp 1698175906
transform 1 0 12656 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_220
timestamp 1698175906
transform 1 0 12992 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_264
timestamp 1698175906
transform 1 0 15456 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 18256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 18704 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 4536 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698175906
transform 1 0 4760 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_75
timestamp 1698175906
transform 1 0 4872 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_125
timestamp 1698175906
transform 1 0 7672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_127
timestamp 1698175906
transform 1 0 7784 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_134
timestamp 1698175906
transform 1 0 8176 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_139
timestamp 1698175906
transform 1 0 8456 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_147
timestamp 1698175906
transform 1 0 8904 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698175906
transform 1 0 10416 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_104
timestamp 1698175906
transform 1 0 6496 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_107
timestamp 1698175906
transform 1 0 6664 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_111
timestamp 1698175906
transform 1 0 6888 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_113
timestamp 1698175906
transform 1 0 7000 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_128
timestamp 1698175906
transform 1 0 7840 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698175906
transform 1 0 8288 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_144
timestamp 1698175906
transform 1 0 8736 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_205
timestamp 1698175906
transform 1 0 12152 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 12376 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_258
timestamp 1698175906
transform 1 0 15120 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_274
timestamp 1698175906
transform 1 0 16016 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 16240 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 18256 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 18704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_115
timestamp 1698175906
transform 1 0 7112 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_125
timestamp 1698175906
transform 1 0 7672 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_130
timestamp 1698175906
transform 1 0 7952 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698175906
transform 1 0 10360 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_185
timestamp 1698175906
transform 1 0 11032 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_236
timestamp 1698175906
transform 1 0 13888 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_240
timestamp 1698175906
transform 1 0 14112 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 14336 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_251
timestamp 1698175906
transform 1 0 14728 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_88
timestamp 1698175906
transform 1 0 5600 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_96
timestamp 1698175906
transform 1 0 6048 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_100
timestamp 1698175906
transform 1 0 6272 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_112
timestamp 1698175906
transform 1 0 6944 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_119
timestamp 1698175906
transform 1 0 7336 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_123
timestamp 1698175906
transform 1 0 7560 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_132
timestamp 1698175906
transform 1 0 8064 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_207
timestamp 1698175906
transform 1 0 12264 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 12376 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_214
timestamp 1698175906
transform 1 0 12656 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_255
timestamp 1698175906
transform 1 0 14952 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_271
timestamp 1698175906
transform 1 0 15848 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 16296 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 2240 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 2464 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_69
timestamp 1698175906
transform 1 0 4536 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_73
timestamp 1698175906
transform 1 0 4760 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_75
timestamp 1698175906
transform 1 0 4872 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_120
timestamp 1698175906
transform 1 0 7392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_160
timestamp 1698175906
transform 1 0 9632 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_204
timestamp 1698175906
transform 1 0 12096 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_220
timestamp 1698175906
transform 1 0 12992 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_233
timestamp 1698175906
transform 1 0 13720 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_241
timestamp 1698175906
transform 1 0 14168 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_251
timestamp 1698175906
transform 1 0 14728 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 2240 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 4032 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 4480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_80
timestamp 1698175906
transform 1 0 5152 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_115
timestamp 1698175906
transform 1 0 7112 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_117
timestamp 1698175906
transform 1 0 7224 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_122
timestamp 1698175906
transform 1 0 7504 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_126
timestamp 1698175906
transform 1 0 7728 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698175906
transform 1 0 8288 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_152
timestamp 1698175906
transform 1 0 9184 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_154
timestamp 1698175906
transform 1 0 9296 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_174
timestamp 1698175906
transform 1 0 10416 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_184
timestamp 1698175906
transform 1 0 10976 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_192
timestamp 1698175906
transform 1 0 11424 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_196
timestamp 1698175906
transform 1 0 11648 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_198
timestamp 1698175906
transform 1 0 11760 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_205
timestamp 1698175906
transform 1 0 12152 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_220
timestamp 1698175906
transform 1 0 12992 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_255
timestamp 1698175906
transform 1 0 14952 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_271
timestamp 1698175906
transform 1 0 15848 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 16296 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 20048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 20160 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_141
timestamp 1698175906
transform 1 0 8568 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_145
timestamp 1698175906
transform 1 0 8792 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_166
timestamp 1698175906
transform 1 0 9968 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_187
timestamp 1698175906
transform 1 0 11144 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_191
timestamp 1698175906
transform 1 0 11368 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_200
timestamp 1698175906
transform 1 0 11872 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_204
timestamp 1698175906
transform 1 0 12096 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_213
timestamp 1698175906
transform 1 0 12600 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 2240 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 4032 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 4480 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698175906
transform 1 0 8288 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_174
timestamp 1698175906
transform 1 0 10416 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_204
timestamp 1698175906
transform 1 0 12096 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698175906
transform 1 0 12320 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_219
timestamp 1698175906
transform 1 0 12936 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_229
timestamp 1698175906
transform 1 0 13496 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_241
timestamp 1698175906
transform 1 0 14168 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_273
timestamp 1698175906
transform 1 0 15960 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698175906
transform 1 0 16184 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 16296 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_123
timestamp 1698175906
transform 1 0 7560 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_127
timestamp 1698175906
transform 1 0 7784 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_134
timestamp 1698175906
transform 1 0 8176 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_138
timestamp 1698175906
transform 1 0 8400 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_141
timestamp 1698175906
transform 1 0 8568 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_149
timestamp 1698175906
transform 1 0 9016 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_151
timestamp 1698175906
transform 1 0 9128 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_158
timestamp 1698175906
transform 1 0 9520 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 10416 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_189
timestamp 1698175906
transform 1 0 11256 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_205
timestamp 1698175906
transform 1 0 12152 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_251
timestamp 1698175906
transform 1 0 14728 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_104
timestamp 1698175906
transform 1 0 6496 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_108
timestamp 1698175906
transform 1 0 6720 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 8456 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_147
timestamp 1698175906
transform 1 0 8904 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_155
timestamp 1698175906
transform 1 0 9352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_157
timestamp 1698175906
transform 1 0 9464 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_173
timestamp 1698175906
transform 1 0 10360 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_189
timestamp 1698175906
transform 1 0 11256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 12376 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_212
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_216
timestamp 1698175906
transform 1 0 12768 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_246
timestamp 1698175906
transform 1 0 14448 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_250
timestamp 1698175906
transform 1 0 14672 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_266
timestamp 1698175906
transform 1 0 15568 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_274
timestamp 1698175906
transform 1 0 16016 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698175906
transform 1 0 16240 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_111
timestamp 1698175906
transform 1 0 6888 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_181
timestamp 1698175906
transform 1 0 10808 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_183
timestamp 1698175906
transform 1 0 10920 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_213
timestamp 1698175906
transform 1 0 12600 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_217
timestamp 1698175906
transform 1 0 12824 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_233
timestamp 1698175906
transform 1 0 13720 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698175906
transform 1 0 14000 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 14224 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 18648 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_104
timestamp 1698175906
transform 1 0 6496 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_120
timestamp 1698175906
transform 1 0 7392 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_128
timestamp 1698175906
transform 1 0 7840 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698175906
transform 1 0 8456 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_146
timestamp 1698175906
transform 1 0 8848 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_177
timestamp 1698175906
transform 1 0 10584 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_181
timestamp 1698175906
transform 1 0 10808 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_197
timestamp 1698175906
transform 1 0 11704 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_205
timestamp 1698175906
transform 1 0 12152 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 12376 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_333
timestamp 1698175906
transform 1 0 19320 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_341
timestamp 1698175906
transform 1 0 19768 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_168
timestamp 1698175906
transform 1 0 10080 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_195
timestamp 1698175906
transform 1 0 11592 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698175906
transform 1 0 12040 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 14000 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 15792 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 16240 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_40
timestamp 1698175906
transform 1 0 2912 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_42
timestamp 1698175906
transform 1 0 3024 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_47
timestamp 1698175906
transform 1 0 3304 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_63
timestamp 1698175906
transform 1 0 4200 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_67
timestamp 1698175906
transform 1 0 4424 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_165
timestamp 1698175906
transform 1 0 9912 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_169
timestamp 1698175906
transform 1 0 10136 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698175906
transform 1 0 10416 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_201
timestamp 1698175906
transform 1 0 11928 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_203
timestamp 1698175906
transform 1 0 12040 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita10_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 3304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita10_26
timestamp 1698175906
transform 1 0 19992 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8792 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 10472 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 18760 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 12096 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 18760 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 10136 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 18760 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 11816 0 1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 8456 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform -1 0 10192 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 2240 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform -1 0 2240 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 2240 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 10472 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13440 400 13496 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 3024 20600 3080 21000 0 FreeSans 224 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 8736 0 8792 400 0 FreeSans 224 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 11760 20600 11816 21000 0 FreeSans 224 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 12432 0 12488 400 0 FreeSans 224 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 10416 0 10472 400 0 FreeSans 224 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 20600 9744 21000 9800 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 11424 0 11480 400 0 FreeSans 224 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 20600 18144 21000 18200 0 FreeSans 224 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 20600 9408 21000 9464 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 11088 0 11144 400 0 FreeSans 224 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 20600 10752 21000 10808 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 10080 20600 10136 21000 0 FreeSans 224 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 20600 9072 21000 9128 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 12432 20600 12488 21000 0 FreeSans 224 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 11760 0 11816 400 0 FreeSans 224 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 8400 20600 8456 21000 0 FreeSans 224 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 9744 0 9800 400 0 FreeSans 224 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 0 12096 400 12152 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 11088 400 11144 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 0 11424 400 11480 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 8064 20600 8120 21000 0 FreeSans 224 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 10416 20600 10472 21000 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 20600 8400 21000 8456 0 FreeSans 224 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 13020 8512 13020 8512 0 _000_
rlabel metal2 9436 13748 9436 13748 0 _001_
rlabel metal3 6076 10780 6076 10780 0 _002_
rlabel metal2 6748 9632 6748 9632 0 _003_
rlabel metal2 7252 8596 7252 8596 0 _004_
rlabel metal2 8428 11228 8428 11228 0 _005_
rlabel metal2 7924 12908 7924 12908 0 _006_
rlabel metal2 6804 11368 6804 11368 0 _007_
rlabel metal2 6412 11004 6412 11004 0 _008_
rlabel metal2 7420 11788 7420 11788 0 _009_
rlabel metal3 9072 7588 9072 7588 0 _010_
rlabel metal2 7420 13692 7420 13692 0 _011_
rlabel metal2 10864 6916 10864 6916 0 _012_
rlabel metal3 9296 13244 9296 13244 0 _013_
rlabel metal2 10864 12068 10864 12068 0 _014_
rlabel metal2 11900 7420 11900 7420 0 _015_
rlabel metal2 9324 6664 9324 6664 0 _016_
rlabel metal2 13860 9408 13860 9408 0 _017_
rlabel metal3 11816 13244 11816 13244 0 _018_
rlabel metal2 13972 9436 13972 9436 0 _019_
rlabel metal2 12628 12936 12628 12936 0 _020_
rlabel metal2 13244 12572 13244 12572 0 _021_
rlabel metal3 13440 10724 13440 10724 0 _022_
rlabel metal2 13580 11368 13580 11368 0 _023_
rlabel metal2 9436 8624 9436 8624 0 _024_
rlabel metal2 6972 11284 6972 11284 0 _025_
rlabel metal2 6860 10864 6860 10864 0 _026_
rlabel metal3 7700 11508 7700 11508 0 _027_
rlabel metal2 9744 7364 9744 7364 0 _028_
rlabel metal2 9800 7644 9800 7644 0 _029_
rlabel metal2 8036 13944 8036 13944 0 _030_
rlabel metal2 8148 13916 8148 13916 0 _031_
rlabel metal3 10780 9604 10780 9604 0 _032_
rlabel metal3 10584 7644 10584 7644 0 _033_
rlabel metal2 9688 11676 9688 11676 0 _034_
rlabel metal2 10948 7000 10948 7000 0 _035_
rlabel metal2 10668 7308 10668 7308 0 _036_
rlabel metal3 10024 13132 10024 13132 0 _037_
rlabel metal3 11228 11956 11228 11956 0 _038_
rlabel metal2 12740 9856 12740 9856 0 _039_
rlabel metal2 10220 11256 10220 11256 0 _040_
rlabel metal2 11676 8008 11676 8008 0 _041_
rlabel metal2 10948 11396 10948 11396 0 _042_
rlabel metal2 11508 10332 11508 10332 0 _043_
rlabel metal2 11788 8176 11788 8176 0 _044_
rlabel metal2 11956 7952 11956 7952 0 _045_
rlabel metal2 9716 6944 9716 6944 0 _046_
rlabel metal2 10276 7000 10276 7000 0 _047_
rlabel metal2 14028 9408 14028 9408 0 _048_
rlabel metal2 14084 9156 14084 9156 0 _049_
rlabel metal2 13020 9408 13020 9408 0 _050_
rlabel metal2 12460 12936 12460 12936 0 _051_
rlabel metal2 12040 13020 12040 13020 0 _052_
rlabel metal2 13468 9408 13468 9408 0 _053_
rlabel metal3 12488 9996 12488 9996 0 _054_
rlabel metal2 13524 9744 13524 9744 0 _055_
rlabel metal3 13216 13468 13216 13468 0 _056_
rlabel metal3 13580 11172 13580 11172 0 _057_
rlabel metal3 11760 12684 11760 12684 0 _058_
rlabel metal3 13664 12348 13664 12348 0 _059_
rlabel metal2 12516 12208 12516 12208 0 _060_
rlabel metal2 14588 11032 14588 11032 0 _061_
rlabel metal2 13412 10584 13412 10584 0 _062_
rlabel metal3 12460 10780 12460 10780 0 _063_
rlabel metal3 14056 10500 14056 10500 0 _064_
rlabel metal2 11564 11004 11564 11004 0 _065_
rlabel metal3 9856 8932 9856 8932 0 _066_
rlabel metal2 9044 8652 9044 8652 0 _067_
rlabel metal2 7924 9408 7924 9408 0 _068_
rlabel metal2 12516 9464 12516 9464 0 _069_
rlabel metal2 13916 9128 13916 9128 0 _070_
rlabel metal2 10864 10388 10864 10388 0 _071_
rlabel metal2 10836 9044 10836 9044 0 _072_
rlabel metal2 9240 9548 9240 9548 0 _073_
rlabel metal3 10640 8372 10640 8372 0 _074_
rlabel metal3 12068 9268 12068 9268 0 _075_
rlabel metal2 12852 8960 12852 8960 0 _076_
rlabel metal2 9996 11424 9996 11424 0 _077_
rlabel metal2 11760 11172 11760 11172 0 _078_
rlabel metal2 12012 10976 12012 10976 0 _079_
rlabel metal2 7532 9576 7532 9576 0 _080_
rlabel metal2 9492 9296 9492 9296 0 _081_
rlabel metal2 10220 10444 10220 10444 0 _082_
rlabel metal2 10220 10192 10220 10192 0 _083_
rlabel metal2 11844 11858 11844 11858 0 _084_
rlabel metal2 12404 8596 12404 8596 0 _085_
rlabel metal2 9940 9016 9940 9016 0 _086_
rlabel metal2 10640 8932 10640 8932 0 _087_
rlabel metal2 13804 9156 13804 9156 0 _088_
rlabel metal2 11200 11620 11200 11620 0 _089_
rlabel metal3 11368 10332 11368 10332 0 _090_
rlabel metal2 8204 11004 8204 11004 0 _091_
rlabel metal2 10780 12768 10780 12768 0 _092_
rlabel metal2 9436 12460 9436 12460 0 _093_
rlabel metal2 8820 13244 8820 13244 0 _094_
rlabel metal3 10192 13468 10192 13468 0 _095_
rlabel metal2 7000 9548 7000 9548 0 _096_
rlabel metal2 9856 7532 9856 7532 0 _097_
rlabel metal3 9940 10388 9940 10388 0 _098_
rlabel metal3 9800 10276 9800 10276 0 _099_
rlabel metal2 10108 11284 10108 11284 0 _100_
rlabel metal2 7952 8932 7952 8932 0 _101_
rlabel metal2 7252 10864 7252 10864 0 _102_
rlabel metal2 11340 11256 11340 11256 0 _103_
rlabel metal2 8428 11816 8428 11816 0 _104_
rlabel metal2 8708 10864 8708 10864 0 _105_
rlabel metal2 8092 12880 8092 12880 0 _106_
rlabel metal2 7112 10780 7112 10780 0 _107_
rlabel metal2 6748 10976 6748 10976 0 _108_
rlabel metal2 7308 11368 7308 11368 0 _109_
rlabel metal3 1239 13468 1239 13468 0 clk
rlabel metal2 11172 10220 11172 10220 0 clknet_0_clk
rlabel metal2 10724 13720 10724 13720 0 clknet_1_0__leaf_clk
rlabel metal2 13468 11172 13468 11172 0 clknet_1_1__leaf_clk
rlabel metal3 6804 9996 6804 9996 0 dut10.count\[0\]
rlabel metal3 7280 9212 7280 9212 0 dut10.count\[1\]
rlabel metal2 9548 8232 9548 8232 0 dut10.count\[2\]
rlabel metal2 9492 11228 9492 11228 0 dut10.count\[3\]
rlabel metal2 8876 3178 8876 3178 0 net1
rlabel metal2 14084 12600 14084 12600 0 net10
rlabel metal2 14868 10836 14868 10836 0 net11
rlabel metal2 14840 11508 14840 11508 0 net12
rlabel metal2 10164 13580 10164 13580 0 net13
rlabel metal2 14196 9772 14196 9772 0 net14
rlabel metal2 12572 13580 12572 13580 0 net15
rlabel metal2 11816 6356 11816 6356 0 net16
rlabel metal2 8316 14140 8316 14140 0 net17
rlabel metal2 9856 1764 9856 1764 0 net18
rlabel metal2 6748 12180 6748 12180 0 net19
rlabel metal2 12096 15960 12096 15960 0 net2
rlabel metal3 3178 11172 3178 11172 0 net20
rlabel metal3 3178 11564 3178 11564 0 net21
rlabel metal2 8820 13748 8820 13748 0 net22
rlabel metal2 10500 14910 10500 14910 0 net23
rlabel metal2 14112 8372 14112 8372 0 net24
rlabel metal2 3108 18956 3108 18956 0 net25
rlabel metal3 20377 18172 20377 18172 0 net26
rlabel metal2 12684 3178 12684 3178 0 net3
rlabel metal2 10556 3178 10556 3178 0 net4
rlabel metal2 15372 9212 15372 9212 0 net5
rlabel metal2 12292 2982 12292 2982 0 net6
rlabel metal2 15036 9184 15036 9184 0 net7
rlabel metal2 11620 6160 11620 6160 0 net8
rlabel metal2 14364 13300 14364 13300 0 net9
rlabel metal2 8764 1211 8764 1211 0 segm[10]
rlabel metal2 11788 19873 11788 19873 0 segm[11]
rlabel metal2 12460 1211 12460 1211 0 segm[12]
rlabel metal2 10444 1211 10444 1211 0 segm[13]
rlabel metal2 20020 9828 20020 9828 0 segm[1]
rlabel metal2 11452 1099 11452 1099 0 segm[2]
rlabel metal2 20020 9548 20020 9548 0 segm[4]
rlabel metal2 11116 1043 11116 1043 0 segm[5]
rlabel metal2 20020 13356 20020 13356 0 segm[6]
rlabel metal2 20020 12908 20020 12908 0 segm[7]
rlabel metal2 20020 11172 20020 11172 0 segm[8]
rlabel metal2 20020 10752 20020 10752 0 segm[9]
rlabel metal2 10108 19677 10108 19677 0 sel[0]
rlabel metal3 20321 9100 20321 9100 0 sel[10]
rlabel metal2 12460 19677 12460 19677 0 sel[11]
rlabel metal2 11788 427 11788 427 0 sel[1]
rlabel metal2 8428 19873 8428 19873 0 sel[2]
rlabel metal2 9772 1015 9772 1015 0 sel[3]
rlabel metal3 679 12124 679 12124 0 sel[4]
rlabel metal3 679 11116 679 11116 0 sel[5]
rlabel metal3 679 11452 679 11452 0 sel[6]
rlabel metal2 8092 19677 8092 19677 0 sel[7]
rlabel metal2 10444 19873 10444 19873 0 sel[8]
rlabel metal2 20020 8652 20020 8652 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
