magic
tech gf180mcuD
magscale 1 5
timestamp 1699642722
<< obsm1 >>
rect 672 1538 20328 19305
<< metal2 >>
rect 8064 20600 8120 21000
rect 9408 20600 9464 21000
rect 9744 20600 9800 21000
rect 10080 20600 10136 21000
rect 10752 20600 10808 21000
rect 12096 20600 12152 21000
rect 12768 20600 12824 21000
rect 13104 20600 13160 21000
rect 13440 20600 13496 21000
rect 8064 0 8120 400
rect 9072 0 9128 400
rect 9744 0 9800 400
rect 10080 0 10136 400
rect 10416 0 10472 400
<< obsm2 >>
rect 966 20570 8034 20600
rect 8150 20570 9378 20600
rect 9494 20570 9714 20600
rect 9830 20570 10050 20600
rect 10166 20570 10722 20600
rect 10838 20570 12066 20600
rect 12182 20570 12738 20600
rect 12854 20570 13074 20600
rect 13190 20570 13410 20600
rect 13526 20570 20146 20600
rect 966 430 20146 20570
rect 966 400 8034 430
rect 8150 400 9042 430
rect 9158 400 9714 430
rect 9830 400 10050 430
rect 10166 400 10386 430
rect 10502 400 20146 430
<< metal3 >>
rect 0 14112 400 14168
rect 0 12768 400 12824
rect 20600 12432 21000 12488
rect 0 12096 400 12152
rect 20600 11088 21000 11144
rect 20600 10752 21000 10808
rect 20600 10416 21000 10472
rect 0 9072 400 9128
rect 20600 9072 21000 9128
rect 0 8736 400 8792
rect 20600 8400 21000 8456
rect 0 8064 400 8120
rect 20600 5376 21000 5432
<< obsm3 >>
rect 400 14198 20600 19250
rect 430 14082 20600 14198
rect 400 12854 20600 14082
rect 430 12738 20600 12854
rect 400 12518 20600 12738
rect 400 12402 20570 12518
rect 400 12182 20600 12402
rect 430 12066 20600 12182
rect 400 11174 20600 12066
rect 400 11058 20570 11174
rect 400 10838 20600 11058
rect 400 10722 20570 10838
rect 400 10502 20600 10722
rect 400 10386 20570 10502
rect 400 9158 20600 10386
rect 430 9042 20570 9158
rect 400 8822 20600 9042
rect 430 8706 20600 8822
rect 400 8486 20600 8706
rect 400 8370 20570 8486
rect 400 8150 20600 8370
rect 430 8034 20600 8150
rect 400 5462 20600 8034
rect 400 5346 20570 5462
rect 400 1554 20600 5346
<< metal4 >>
rect 2224 1538 2384 19238
rect 9904 1538 10064 19238
rect 17584 1538 17744 19238
<< labels >>
rlabel metal3 s 0 14112 400 14168 6 clk
port 1 nsew signal input
rlabel metal2 s 13440 20600 13496 21000 6 segm[0]
port 2 nsew signal output
rlabel metal3 s 20600 10416 21000 10472 6 segm[10]
port 3 nsew signal output
rlabel metal2 s 9744 20600 9800 21000 6 segm[11]
port 4 nsew signal output
rlabel metal3 s 0 8064 400 8120 6 segm[12]
port 5 nsew signal output
rlabel metal3 s 20600 10752 21000 10808 6 segm[13]
port 6 nsew signal output
rlabel metal2 s 10416 0 10472 400 6 segm[1]
port 7 nsew signal output
rlabel metal3 s 0 9072 400 9128 6 segm[2]
port 8 nsew signal output
rlabel metal3 s 20600 5376 21000 5432 6 segm[3]
port 9 nsew signal output
rlabel metal2 s 9744 0 9800 400 6 segm[4]
port 10 nsew signal output
rlabel metal2 s 13104 20600 13160 21000 6 segm[5]
port 11 nsew signal output
rlabel metal3 s 0 12096 400 12152 6 segm[6]
port 12 nsew signal output
rlabel metal3 s 20600 8400 21000 8456 6 segm[7]
port 13 nsew signal output
rlabel metal3 s 20600 9072 21000 9128 6 segm[8]
port 14 nsew signal output
rlabel metal2 s 12768 20600 12824 21000 6 segm[9]
port 15 nsew signal output
rlabel metal2 s 10752 20600 10808 21000 6 sel[0]
port 16 nsew signal output
rlabel metal3 s 20600 12432 21000 12488 6 sel[10]
port 17 nsew signal output
rlabel metal2 s 12096 20600 12152 21000 6 sel[11]
port 18 nsew signal output
rlabel metal2 s 10080 20600 10136 21000 6 sel[1]
port 19 nsew signal output
rlabel metal3 s 0 12768 400 12824 6 sel[2]
port 20 nsew signal output
rlabel metal2 s 9408 20600 9464 21000 6 sel[3]
port 21 nsew signal output
rlabel metal2 s 8064 20600 8120 21000 6 sel[4]
port 22 nsew signal output
rlabel metal2 s 10080 0 10136 400 6 sel[5]
port 23 nsew signal output
rlabel metal2 s 9072 0 9128 400 6 sel[6]
port 24 nsew signal output
rlabel metal3 s 0 8736 400 8792 6 sel[7]
port 25 nsew signal output
rlabel metal2 s 8064 0 8120 400 6 sel[8]
port 26 nsew signal output
rlabel metal3 s 20600 11088 21000 11144 6 sel[9]
port 27 nsew signal output
rlabel metal4 s 2224 1538 2384 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 19238 6 vss
port 29 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 21000 21000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 485802
string GDS_FILE /home/urielcho/Proyectos_caravel/ITA23_GFMPW1b/openlane/ita57/runs/23_11_10_12_56/results/signoff/ita57.magic.gds
string GDS_START 164258
<< end >>

