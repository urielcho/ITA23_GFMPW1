magic
tech gf180mcuD
magscale 1 5
timestamp 1699643673
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 8975 19137 9001 19143
rect 8975 19105 9001 19111
rect 11215 19137 11241 19143
rect 11215 19105 11241 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 14687 19137 14713 19143
rect 14687 19105 14713 19111
rect 8465 18999 8471 19025
rect 8497 18999 8503 19025
rect 10817 18999 10823 19025
rect 10849 18999 10855 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 14289 18999 14295 19025
rect 14321 18999 14327 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 11047 18745 11073 18751
rect 11047 18713 11073 18719
rect 13119 18745 13145 18751
rect 13119 18713 13145 18719
rect 10537 18607 10543 18633
rect 10569 18607 10575 18633
rect 12721 18607 12727 18633
rect 12753 18607 12759 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 11159 18353 11185 18359
rect 11159 18321 11185 18327
rect 13399 18353 13425 18359
rect 13399 18321 13425 18327
rect 10649 18215 10655 18241
rect 10681 18215 10687 18241
rect 12889 18215 12895 18241
rect 12921 18215 12927 18241
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 11943 14041 11969 14047
rect 11943 14009 11969 14015
rect 11999 13929 12025 13935
rect 11999 13897 12025 13903
rect 11943 13817 11969 13823
rect 11943 13785 11969 13791
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 10369 13567 10375 13593
rect 10401 13567 10407 13593
rect 12329 13567 12335 13593
rect 12361 13567 12367 13593
rect 12559 13537 12585 13543
rect 8913 13511 8919 13537
rect 8945 13511 8951 13537
rect 10929 13511 10935 13537
rect 10961 13511 10967 13537
rect 12559 13505 12585 13511
rect 12727 13537 12753 13543
rect 12727 13505 12753 13511
rect 9305 13455 9311 13481
rect 9337 13455 9343 13481
rect 11265 13455 11271 13481
rect 11297 13455 11303 13481
rect 12889 13455 12895 13481
rect 12921 13455 12927 13481
rect 13225 13455 13231 13481
rect 13257 13455 13263 13481
rect 8751 13425 8777 13431
rect 8751 13393 8777 13399
rect 13063 13425 13089 13431
rect 13063 13393 13089 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 8079 13257 8105 13263
rect 8079 13225 8105 13231
rect 10375 13257 10401 13263
rect 10375 13225 10401 13231
rect 11327 13257 11353 13263
rect 11327 13225 11353 13231
rect 11943 13257 11969 13263
rect 11943 13225 11969 13231
rect 13175 13257 13201 13263
rect 13175 13225 13201 13231
rect 11439 13201 11465 13207
rect 11439 13169 11465 13175
rect 11495 13201 11521 13207
rect 11495 13169 11521 13175
rect 12671 13201 12697 13207
rect 12671 13169 12697 13175
rect 12727 13201 12753 13207
rect 12727 13169 12753 13175
rect 8135 13145 8161 13151
rect 10319 13145 10345 13151
rect 6449 13119 6455 13145
rect 6481 13119 6487 13145
rect 8689 13119 8695 13145
rect 8721 13119 8727 13145
rect 8135 13113 8161 13119
rect 10319 13113 10345 13119
rect 11999 13145 12025 13151
rect 11999 13113 12025 13119
rect 12559 13145 12585 13151
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 12559 13113 12585 13119
rect 8359 13089 8385 13095
rect 10655 13089 10681 13095
rect 6785 13063 6791 13089
rect 6817 13063 6823 13089
rect 7849 13063 7855 13089
rect 7881 13063 7887 13089
rect 9081 13063 9087 13089
rect 9113 13063 9119 13089
rect 10145 13063 10151 13089
rect 10177 13063 10183 13089
rect 8359 13057 8385 13063
rect 10655 13057 10681 13063
rect 8079 13033 8105 13039
rect 8079 13001 8105 13007
rect 10375 13033 10401 13039
rect 10375 13001 10401 13007
rect 11943 13033 11969 13039
rect 11943 13001 11969 13007
rect 20007 13033 20033 13039
rect 20007 13001 20033 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 967 12809 993 12815
rect 967 12777 993 12783
rect 7127 12809 7153 12815
rect 7127 12777 7153 12783
rect 9759 12809 9785 12815
rect 11881 12783 11887 12809
rect 11913 12783 11919 12809
rect 13001 12783 13007 12809
rect 13033 12783 13039 12809
rect 9759 12777 9785 12783
rect 7407 12753 7433 12759
rect 2137 12727 2143 12753
rect 2169 12727 2175 12753
rect 7407 12721 7433 12727
rect 9535 12753 9561 12759
rect 9535 12721 9561 12727
rect 10039 12753 10065 12759
rect 13231 12753 13257 12759
rect 11545 12727 11551 12753
rect 11577 12727 11583 12753
rect 10039 12721 10065 12727
rect 13231 12721 13257 12727
rect 13399 12753 13425 12759
rect 13399 12721 13425 12727
rect 6175 12697 6201 12703
rect 6175 12665 6201 12671
rect 6231 12697 6257 12703
rect 9479 12697 9505 12703
rect 8129 12671 8135 12697
rect 8161 12671 8167 12697
rect 8633 12671 8639 12697
rect 8665 12671 8671 12697
rect 6231 12665 6257 12671
rect 9479 12665 9505 12671
rect 13287 12697 13313 12703
rect 13287 12665 13313 12671
rect 13567 12697 13593 12703
rect 13567 12665 13593 12671
rect 13623 12697 13649 12703
rect 13623 12665 13649 12671
rect 6063 12641 6089 12647
rect 6063 12609 6089 12615
rect 7071 12641 7097 12647
rect 7071 12609 7097 12615
rect 7183 12641 7209 12647
rect 7183 12609 7209 12615
rect 8303 12641 8329 12647
rect 8303 12609 8329 12615
rect 8471 12641 8497 12647
rect 8471 12609 8497 12615
rect 9367 12641 9393 12647
rect 9367 12609 9393 12615
rect 9703 12641 9729 12647
rect 9703 12609 9729 12615
rect 9815 12641 9841 12647
rect 9815 12609 9841 12615
rect 13455 12641 13481 12647
rect 13455 12609 13481 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 13281 12391 13287 12417
rect 13313 12391 13319 12417
rect 2137 12335 2143 12361
rect 2169 12335 2175 12361
rect 6505 12335 6511 12361
rect 6537 12335 6543 12361
rect 8409 12335 8415 12361
rect 8441 12335 8447 12361
rect 9417 12335 9423 12361
rect 9449 12335 9455 12361
rect 12945 12335 12951 12361
rect 12977 12335 12983 12361
rect 6735 12305 6761 12311
rect 8751 12305 8777 12311
rect 5049 12279 5055 12305
rect 5081 12279 5087 12305
rect 6113 12279 6119 12305
rect 6145 12279 6151 12305
rect 6953 12279 6959 12305
rect 6985 12279 6991 12305
rect 8017 12279 8023 12305
rect 8049 12279 8055 12305
rect 6735 12273 6761 12279
rect 8751 12273 8777 12279
rect 9199 12305 9225 12311
rect 14575 12305 14601 12311
rect 9753 12279 9759 12305
rect 9785 12279 9791 12305
rect 10817 12279 10823 12305
rect 10849 12279 10855 12305
rect 14345 12279 14351 12305
rect 14377 12279 14383 12305
rect 9199 12273 9225 12279
rect 14575 12273 14601 12279
rect 967 12249 993 12255
rect 967 12217 993 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 8023 12081 8049 12087
rect 8023 12049 8049 12055
rect 8247 12081 8273 12087
rect 8247 12049 8273 12055
rect 9367 12081 9393 12087
rect 9367 12049 9393 12055
rect 9423 12081 9449 12087
rect 9423 12049 9449 12055
rect 6399 12025 6425 12031
rect 6399 11993 6425 11999
rect 20007 12025 20033 12031
rect 20007 11993 20033 11999
rect 6119 11969 6145 11975
rect 6119 11937 6145 11943
rect 8527 11969 8553 11975
rect 8527 11937 8553 11943
rect 8639 11969 8665 11975
rect 8639 11937 8665 11943
rect 9647 11969 9673 11975
rect 9647 11937 9673 11943
rect 9759 11969 9785 11975
rect 18825 11943 18831 11969
rect 18857 11943 18863 11969
rect 9759 11937 9785 11943
rect 8023 11913 8049 11919
rect 8023 11881 8049 11887
rect 8079 11913 8105 11919
rect 8079 11881 8105 11887
rect 8359 11913 8385 11919
rect 8359 11881 8385 11887
rect 9479 11913 9505 11919
rect 9479 11881 9505 11887
rect 9983 11913 10009 11919
rect 9983 11881 10009 11887
rect 10039 11913 10065 11919
rect 10039 11881 10065 11887
rect 6343 11857 6369 11863
rect 6343 11825 6369 11831
rect 6455 11857 6481 11863
rect 7463 11857 7489 11863
rect 7289 11831 7295 11857
rect 7321 11831 7327 11857
rect 6455 11825 6481 11831
rect 7463 11825 7489 11831
rect 8695 11857 8721 11863
rect 8695 11825 8721 11831
rect 10151 11857 10177 11863
rect 10151 11825 10177 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 9983 11689 10009 11695
rect 9983 11657 10009 11663
rect 6567 11633 6593 11639
rect 6567 11601 6593 11607
rect 6623 11633 6649 11639
rect 6623 11601 6649 11607
rect 8303 11633 8329 11639
rect 8303 11601 8329 11607
rect 20119 11633 20145 11639
rect 20119 11601 20145 11607
rect 8247 11577 8273 11583
rect 2137 11551 2143 11577
rect 2169 11551 2175 11577
rect 6281 11551 6287 11577
rect 6313 11551 6319 11577
rect 8247 11545 8273 11551
rect 9927 11577 9953 11583
rect 9927 11545 9953 11551
rect 10039 11577 10065 11583
rect 10039 11545 10065 11551
rect 10151 11577 10177 11583
rect 12671 11577 12697 11583
rect 14575 11577 14601 11583
rect 10929 11551 10935 11577
rect 10961 11551 10967 11577
rect 12945 11551 12951 11577
rect 12977 11551 12983 11577
rect 10151 11545 10177 11551
rect 12671 11545 12697 11551
rect 14575 11545 14601 11551
rect 6847 11521 6873 11527
rect 4825 11495 4831 11521
rect 4857 11495 4863 11521
rect 5889 11495 5895 11521
rect 5921 11495 5927 11521
rect 11265 11495 11271 11521
rect 11297 11495 11303 11521
rect 12329 11495 12335 11521
rect 12361 11495 12367 11521
rect 13281 11495 13287 11521
rect 13313 11495 13319 11521
rect 14345 11495 14351 11521
rect 14377 11495 14383 11521
rect 6847 11489 6873 11495
rect 967 11465 993 11471
rect 967 11433 993 11439
rect 6567 11465 6593 11471
rect 6567 11433 6593 11439
rect 8303 11465 8329 11471
rect 8303 11433 8329 11439
rect 10263 11465 10289 11471
rect 10263 11433 10289 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 11103 11297 11129 11303
rect 11103 11265 11129 11271
rect 12223 11297 12249 11303
rect 12223 11265 12249 11271
rect 5951 11241 5977 11247
rect 5951 11209 5977 11215
rect 8527 11241 8553 11247
rect 8527 11209 8553 11215
rect 13007 11241 13033 11247
rect 13007 11209 13033 11215
rect 13455 11241 13481 11247
rect 13455 11209 13481 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 8079 11185 8105 11191
rect 8079 11153 8105 11159
rect 8415 11185 8441 11191
rect 8415 11153 8441 11159
rect 8695 11185 8721 11191
rect 8695 11153 8721 11159
rect 10711 11185 10737 11191
rect 10711 11153 10737 11159
rect 10823 11185 10849 11191
rect 10823 11153 10849 11159
rect 10991 11185 11017 11191
rect 10991 11153 11017 11159
rect 11999 11185 12025 11191
rect 11999 11153 12025 11159
rect 12391 11185 12417 11191
rect 12391 11153 12417 11159
rect 13063 11185 13089 11191
rect 13063 11153 13089 11159
rect 13287 11185 13313 11191
rect 13287 11153 13313 11159
rect 13343 11185 13369 11191
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 13343 11153 13369 11159
rect 5783 11129 5809 11135
rect 5783 11097 5809 11103
rect 6903 11129 6929 11135
rect 6903 11097 6929 11103
rect 8751 11129 8777 11135
rect 12055 11129 12081 11135
rect 11545 11103 11551 11129
rect 11577 11103 11583 11129
rect 11825 11103 11831 11129
rect 11857 11103 11863 11129
rect 8751 11097 8777 11103
rect 12055 11097 12081 11103
rect 12167 11129 12193 11135
rect 12167 11097 12193 11103
rect 12503 11129 12529 11135
rect 12503 11097 12529 11103
rect 13623 11129 13649 11135
rect 13623 11097 13649 11103
rect 5895 11073 5921 11079
rect 5895 11041 5921 11047
rect 6007 11073 6033 11079
rect 6007 11041 6033 11047
rect 6735 11073 6761 11079
rect 6735 11041 6761 11047
rect 6847 11073 6873 11079
rect 10655 11073 10681 11079
rect 7905 11047 7911 11073
rect 7937 11047 7943 11073
rect 8241 11047 8247 11073
rect 8273 11047 8279 11073
rect 6847 11041 6873 11047
rect 10655 11041 10681 11047
rect 12279 11073 12305 11079
rect 12279 11041 12305 11047
rect 12951 11073 12977 11079
rect 12951 11041 12977 11047
rect 13511 11073 13537 11079
rect 13511 11041 13537 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 10375 10905 10401 10911
rect 10375 10873 10401 10879
rect 10823 10905 10849 10911
rect 10823 10873 10849 10879
rect 10935 10905 10961 10911
rect 10935 10873 10961 10879
rect 13287 10905 13313 10911
rect 14177 10879 14183 10905
rect 14209 10879 14215 10905
rect 13287 10873 13313 10879
rect 8863 10849 8889 10855
rect 6673 10823 6679 10849
rect 6705 10823 6711 10849
rect 8863 10817 8889 10823
rect 10487 10849 10513 10855
rect 10487 10817 10513 10823
rect 11383 10849 11409 10855
rect 12055 10849 12081 10855
rect 11545 10823 11551 10849
rect 11577 10823 11583 10849
rect 11383 10817 11409 10823
rect 12055 10817 12081 10823
rect 12615 10849 12641 10855
rect 12615 10817 12641 10823
rect 12839 10849 12865 10855
rect 14351 10849 14377 10855
rect 13673 10823 13679 10849
rect 13705 10823 13711 10849
rect 12839 10817 12865 10823
rect 14351 10817 14377 10823
rect 14407 10849 14433 10855
rect 14407 10817 14433 10823
rect 8695 10793 8721 10799
rect 6337 10767 6343 10793
rect 6369 10767 6375 10793
rect 8695 10761 8721 10767
rect 10543 10793 10569 10799
rect 10543 10761 10569 10767
rect 10655 10793 10681 10799
rect 10655 10761 10681 10767
rect 11271 10793 11297 10799
rect 13399 10793 13425 10799
rect 14015 10793 14041 10799
rect 11489 10767 11495 10793
rect 11521 10767 11527 10793
rect 11825 10767 11831 10793
rect 11857 10767 11863 10793
rect 11937 10767 11943 10793
rect 11969 10767 11975 10793
rect 12721 10767 12727 10793
rect 12753 10767 12759 10793
rect 13169 10767 13175 10793
rect 13201 10767 13207 10793
rect 13505 10767 13511 10793
rect 13537 10767 13543 10793
rect 13785 10767 13791 10793
rect 13817 10767 13823 10793
rect 11271 10761 11297 10767
rect 13399 10761 13425 10767
rect 14015 10761 14041 10767
rect 14519 10793 14545 10799
rect 18825 10767 18831 10793
rect 18857 10767 18863 10793
rect 14519 10761 14545 10767
rect 7967 10737 7993 10743
rect 7737 10711 7743 10737
rect 7769 10711 7775 10737
rect 7967 10705 7993 10711
rect 9143 10737 9169 10743
rect 9143 10705 9169 10711
rect 9759 10737 9785 10743
rect 11887 10737 11913 10743
rect 10873 10711 10879 10737
rect 10905 10711 10911 10737
rect 11657 10711 11663 10737
rect 11689 10711 11695 10737
rect 9759 10705 9785 10711
rect 11887 10705 11913 10711
rect 12783 10737 12809 10743
rect 12783 10705 12809 10711
rect 13343 10737 13369 10743
rect 13343 10705 13369 10711
rect 9255 10681 9281 10687
rect 9255 10649 9281 10655
rect 9367 10681 9393 10687
rect 9367 10649 9393 10655
rect 9591 10681 9617 10687
rect 9591 10649 9617 10655
rect 20007 10681 20033 10687
rect 20007 10649 20033 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 10767 10513 10793 10519
rect 10767 10481 10793 10487
rect 12889 10431 12895 10457
rect 12921 10431 12927 10457
rect 10655 10401 10681 10407
rect 10033 10375 10039 10401
rect 10065 10375 10071 10401
rect 11769 10375 11775 10401
rect 11801 10375 11807 10401
rect 10655 10369 10681 10375
rect 7961 10319 7967 10345
rect 7993 10319 7999 10345
rect 11103 10289 11129 10295
rect 10929 10263 10935 10289
rect 10961 10263 10967 10289
rect 11265 10263 11271 10289
rect 11297 10263 11303 10289
rect 11103 10257 11129 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 12839 10121 12865 10127
rect 12839 10089 12865 10095
rect 8079 10065 8105 10071
rect 8079 10033 8105 10039
rect 8247 10065 8273 10071
rect 8247 10033 8273 10039
rect 8415 10065 8441 10071
rect 8415 10033 8441 10039
rect 8975 10065 9001 10071
rect 12895 10065 12921 10071
rect 9361 10039 9367 10065
rect 9393 10039 9399 10065
rect 11713 10039 11719 10065
rect 11745 10039 11751 10065
rect 8975 10033 9001 10039
rect 12895 10033 12921 10039
rect 7911 10009 7937 10015
rect 5497 9983 5503 10009
rect 5529 9983 5535 10009
rect 5833 9983 5839 10009
rect 5865 9983 5871 10009
rect 7911 9977 7937 9983
rect 8695 10009 8721 10015
rect 12671 10009 12697 10015
rect 9249 9983 9255 10009
rect 9281 9983 9287 10009
rect 9753 9983 9759 10009
rect 9785 9983 9791 10009
rect 8695 9977 8721 9983
rect 12671 9977 12697 9983
rect 13007 10009 13033 10015
rect 13337 9983 13343 10009
rect 13369 9983 13375 10009
rect 13729 9983 13735 10009
rect 13761 9983 13767 10009
rect 13007 9977 13033 9983
rect 7127 9953 7153 9959
rect 6897 9927 6903 9953
rect 6929 9927 6935 9953
rect 14793 9927 14799 9953
rect 14825 9927 14831 9953
rect 7127 9921 7153 9927
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 8863 9729 8889 9735
rect 8863 9697 8889 9703
rect 12503 9729 12529 9735
rect 12503 9697 12529 9703
rect 8751 9673 8777 9679
rect 7849 9647 7855 9673
rect 7881 9647 7887 9673
rect 8297 9647 8303 9673
rect 8329 9647 8335 9673
rect 8751 9641 8777 9647
rect 12447 9673 12473 9679
rect 12447 9641 12473 9647
rect 7407 9617 7433 9623
rect 7407 9585 7433 9591
rect 7743 9617 7769 9623
rect 9535 9617 9561 9623
rect 7905 9591 7911 9617
rect 7937 9591 7943 9617
rect 7743 9585 7769 9591
rect 9535 9585 9561 9591
rect 9703 9617 9729 9623
rect 11607 9617 11633 9623
rect 11943 9617 11969 9623
rect 9865 9591 9871 9617
rect 9897 9591 9903 9617
rect 10201 9591 10207 9617
rect 10233 9591 10239 9617
rect 10817 9591 10823 9617
rect 10849 9591 10855 9617
rect 11769 9591 11775 9617
rect 11801 9591 11807 9617
rect 12329 9591 12335 9617
rect 12361 9591 12367 9617
rect 13281 9591 13287 9617
rect 13313 9591 13319 9617
rect 9703 9585 9729 9591
rect 11607 9585 11633 9591
rect 11943 9585 11969 9591
rect 7575 9561 7601 9567
rect 7575 9529 7601 9535
rect 9199 9561 9225 9567
rect 9199 9529 9225 9535
rect 9591 9561 9617 9567
rect 11887 9561 11913 9567
rect 9977 9535 9983 9561
rect 10009 9535 10015 9561
rect 10705 9535 10711 9561
rect 10737 9535 10743 9561
rect 11153 9535 11159 9561
rect 11185 9535 11191 9561
rect 11321 9535 11327 9561
rect 11353 9535 11359 9561
rect 9591 9529 9617 9535
rect 11887 9529 11913 9535
rect 13063 9561 13089 9567
rect 13063 9529 13089 9535
rect 13119 9561 13145 9567
rect 13119 9529 13145 9535
rect 8079 9505 8105 9511
rect 12951 9505 12977 9511
rect 9025 9479 9031 9505
rect 9057 9479 9063 9505
rect 9361 9479 9367 9505
rect 9393 9479 9399 9505
rect 10313 9479 10319 9505
rect 10345 9479 10351 9505
rect 11545 9479 11551 9505
rect 11577 9479 11583 9505
rect 12161 9479 12167 9505
rect 12193 9479 12199 9505
rect 8079 9473 8105 9479
rect 12951 9473 12977 9479
rect 13007 9505 13033 9511
rect 13007 9473 13033 9479
rect 13567 9505 13593 9511
rect 13567 9473 13593 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 8863 9337 8889 9343
rect 11943 9337 11969 9343
rect 10089 9311 10095 9337
rect 10121 9311 10127 9337
rect 8863 9305 8889 9311
rect 11943 9305 11969 9311
rect 10767 9281 10793 9287
rect 10767 9249 10793 9255
rect 10823 9281 10849 9287
rect 11601 9255 11607 9281
rect 11633 9255 11639 9281
rect 11769 9255 11775 9281
rect 11801 9255 11807 9281
rect 10823 9249 10849 9255
rect 9927 9225 9953 9231
rect 5721 9199 5727 9225
rect 5753 9199 5759 9225
rect 7513 9199 7519 9225
rect 7545 9199 7551 9225
rect 8745 9199 8751 9225
rect 8777 9199 8783 9225
rect 9137 9199 9143 9225
rect 9169 9199 9175 9225
rect 9249 9199 9255 9225
rect 9281 9199 9287 9225
rect 9585 9199 9591 9225
rect 9617 9199 9623 9225
rect 9927 9193 9953 9199
rect 10487 9225 10513 9231
rect 10487 9193 10513 9199
rect 10655 9225 10681 9231
rect 10655 9193 10681 9199
rect 11439 9225 11465 9231
rect 13113 9199 13119 9225
rect 13145 9199 13151 9225
rect 18825 9199 18831 9225
rect 18857 9199 18863 9225
rect 11439 9193 11465 9199
rect 7407 9169 7433 9175
rect 6113 9143 6119 9169
rect 6145 9143 6151 9169
rect 7177 9143 7183 9169
rect 7209 9143 7215 9169
rect 7407 9137 7433 9143
rect 7743 9169 7769 9175
rect 7743 9137 7769 9143
rect 10991 9169 11017 9175
rect 14799 9169 14825 9175
rect 13505 9143 13511 9169
rect 13537 9143 13543 9169
rect 14569 9143 14575 9169
rect 14601 9143 14607 9169
rect 10991 9137 11017 9143
rect 14799 9137 14825 9143
rect 7351 9113 7377 9119
rect 7351 9081 7377 9087
rect 9703 9113 9729 9119
rect 9703 9081 9729 9087
rect 10543 9113 10569 9119
rect 10543 9081 10569 9087
rect 11047 9113 11073 9119
rect 11047 9081 11073 9087
rect 20007 9113 20033 9119
rect 20007 9081 20033 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 9143 8945 9169 8951
rect 9143 8913 9169 8919
rect 967 8889 993 8895
rect 20007 8889 20033 8895
rect 6281 8863 6287 8889
rect 6313 8863 6319 8889
rect 9305 8863 9311 8889
rect 9337 8863 9343 8889
rect 12385 8863 12391 8889
rect 12417 8863 12423 8889
rect 13169 8863 13175 8889
rect 13201 8863 13207 8889
rect 13393 8863 13399 8889
rect 13425 8863 13431 8889
rect 967 8857 993 8863
rect 20007 8857 20033 8863
rect 6735 8833 6761 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 6735 8801 6761 8807
rect 6847 8833 6873 8839
rect 6847 8801 6873 8807
rect 7631 8833 7657 8839
rect 7631 8801 7657 8807
rect 8471 8833 8497 8839
rect 8471 8801 8497 8807
rect 8919 8833 8945 8839
rect 8919 8801 8945 8807
rect 9479 8833 9505 8839
rect 9479 8801 9505 8807
rect 12783 8833 12809 8839
rect 13455 8833 13481 8839
rect 13113 8807 13119 8833
rect 13145 8807 13151 8833
rect 12783 8801 12809 8807
rect 13455 8801 13481 8807
rect 13623 8833 13649 8839
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 13623 8801 13649 8807
rect 6343 8777 6369 8783
rect 6343 8745 6369 8751
rect 6455 8777 6481 8783
rect 6455 8745 6481 8751
rect 7015 8777 7041 8783
rect 7015 8745 7041 8751
rect 7351 8777 7377 8783
rect 7351 8745 7377 8751
rect 8527 8777 8553 8783
rect 9255 8777 9281 8783
rect 8745 8751 8751 8777
rect 8777 8751 8783 8777
rect 8527 8745 8553 8751
rect 9255 8745 9281 8751
rect 12223 8777 12249 8783
rect 12223 8745 12249 8751
rect 12335 8777 12361 8783
rect 12335 8745 12361 8751
rect 12895 8777 12921 8783
rect 12895 8745 12921 8751
rect 12951 8777 12977 8783
rect 12951 8745 12977 8751
rect 6903 8721 6929 8727
rect 6903 8689 6929 8695
rect 7295 8721 7321 8727
rect 7295 8689 7321 8695
rect 7407 8721 7433 8727
rect 7407 8689 7433 8695
rect 8639 8721 8665 8727
rect 13399 8721 13425 8727
rect 9641 8695 9647 8721
rect 9673 8695 9679 8721
rect 8639 8689 8665 8695
rect 13399 8689 13425 8695
rect 13567 8721 13593 8727
rect 13567 8689 13593 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 7407 8553 7433 8559
rect 7407 8521 7433 8527
rect 10599 8553 10625 8559
rect 10599 8521 10625 8527
rect 9087 8497 9113 8503
rect 10711 8497 10737 8503
rect 6113 8471 6119 8497
rect 6145 8471 6151 8497
rect 9193 8471 9199 8497
rect 9225 8471 9231 8497
rect 9087 8465 9113 8471
rect 10711 8465 10737 8471
rect 11271 8497 11297 8503
rect 13281 8471 13287 8497
rect 13313 8471 13319 8497
rect 11271 8465 11297 8471
rect 11047 8441 11073 8447
rect 5721 8415 5727 8441
rect 5753 8415 5759 8441
rect 9473 8415 9479 8441
rect 9505 8415 9511 8441
rect 10929 8415 10935 8441
rect 10961 8415 10967 8441
rect 11047 8409 11073 8415
rect 11103 8441 11129 8447
rect 12945 8415 12951 8441
rect 12977 8415 12983 8441
rect 11103 8409 11129 8415
rect 9143 8385 9169 8391
rect 7177 8359 7183 8385
rect 7209 8359 7215 8385
rect 9143 8353 9169 8359
rect 9311 8385 9337 8391
rect 9311 8353 9337 8359
rect 10655 8385 10681 8391
rect 10655 8353 10681 8359
rect 11215 8385 11241 8391
rect 14575 8385 14601 8391
rect 14345 8359 14351 8385
rect 14377 8359 14383 8385
rect 11215 8353 11241 8359
rect 14575 8353 14601 8359
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 10823 8161 10849 8167
rect 10823 8129 10849 8135
rect 10935 8161 10961 8167
rect 10935 8129 10961 8135
rect 11047 8105 11073 8111
rect 11047 8073 11073 8079
rect 20007 8105 20033 8111
rect 20007 8073 20033 8079
rect 8807 8049 8833 8055
rect 8807 8017 8833 8023
rect 8975 8049 9001 8055
rect 8975 8017 9001 8023
rect 9031 8049 9057 8055
rect 9367 8049 9393 8055
rect 9871 8049 9897 8055
rect 9137 8023 9143 8049
rect 9169 8023 9175 8049
rect 9641 8023 9647 8049
rect 9673 8023 9679 8049
rect 9031 8017 9057 8023
rect 9367 8017 9393 8023
rect 9871 8017 9897 8023
rect 10207 8049 10233 8055
rect 10207 8017 10233 8023
rect 13007 8049 13033 8055
rect 13007 8017 13033 8023
rect 13175 8049 13201 8055
rect 13175 8017 13201 8023
rect 13623 8049 13649 8055
rect 13623 8017 13649 8023
rect 13791 8049 13817 8055
rect 13791 8017 13817 8023
rect 14071 8049 14097 8055
rect 18825 8023 18831 8049
rect 18857 8023 18863 8049
rect 14071 8017 14097 8023
rect 13287 7993 13313 7999
rect 13287 7961 13313 7967
rect 13735 7993 13761 7999
rect 13735 7961 13761 7967
rect 8863 7937 8889 7943
rect 8863 7905 8889 7911
rect 9423 7937 9449 7943
rect 9423 7905 9449 7911
rect 9479 7937 9505 7943
rect 9479 7905 9505 7911
rect 10095 7937 10121 7943
rect 10095 7905 10121 7911
rect 10151 7937 10177 7943
rect 10151 7905 10177 7911
rect 11159 7937 11185 7943
rect 11159 7905 11185 7911
rect 11215 7937 11241 7943
rect 11215 7905 11241 7911
rect 11271 7937 11297 7943
rect 11271 7905 11297 7911
rect 13175 7937 13201 7943
rect 13175 7905 13201 7911
rect 13903 7937 13929 7943
rect 13903 7905 13929 7911
rect 14015 7937 14041 7943
rect 14015 7905 14041 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 11383 7769 11409 7775
rect 8969 7743 8975 7769
rect 9001 7743 9007 7769
rect 9305 7743 9311 7769
rect 9337 7743 9343 7769
rect 11383 7737 11409 7743
rect 14407 7769 14433 7775
rect 14407 7737 14433 7743
rect 6561 7687 6567 7713
rect 6593 7687 6599 7713
rect 9809 7687 9815 7713
rect 9841 7687 9847 7713
rect 13113 7687 13119 7713
rect 13145 7687 13151 7713
rect 8751 7657 8777 7663
rect 9647 7657 9673 7663
rect 6169 7631 6175 7657
rect 6201 7631 6207 7657
rect 9081 7631 9087 7657
rect 9113 7631 9119 7657
rect 9417 7631 9423 7657
rect 9449 7631 9455 7657
rect 8751 7625 8777 7631
rect 9647 7625 9673 7631
rect 11159 7657 11185 7663
rect 11495 7657 11521 7663
rect 11321 7631 11327 7657
rect 11353 7631 11359 7657
rect 12721 7631 12727 7657
rect 12753 7631 12759 7657
rect 11159 7625 11185 7631
rect 11495 7625 11521 7631
rect 7855 7601 7881 7607
rect 7625 7575 7631 7601
rect 7657 7575 7663 7601
rect 7855 7569 7881 7575
rect 8695 7601 8721 7607
rect 8695 7569 8721 7575
rect 11439 7601 11465 7607
rect 14177 7575 14183 7601
rect 14209 7575 14215 7601
rect 11439 7569 11465 7575
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 11551 7321 11577 7327
rect 8185 7295 8191 7321
rect 8217 7295 8223 7321
rect 9249 7295 9255 7321
rect 9281 7295 9287 7321
rect 11551 7289 11577 7295
rect 11887 7321 11913 7327
rect 11887 7289 11913 7295
rect 7849 7239 7855 7265
rect 7881 7239 7887 7265
rect 11657 7239 11663 7265
rect 11689 7239 11695 7265
rect 11993 7239 11999 7265
rect 12025 7239 12031 7265
rect 11495 7209 11521 7215
rect 11495 7177 11521 7183
rect 11831 7209 11857 7215
rect 11831 7177 11857 7183
rect 9479 7153 9505 7159
rect 9479 7121 9505 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 8919 6985 8945 6991
rect 8919 6953 8945 6959
rect 9871 6985 9897 6991
rect 9871 6953 9897 6959
rect 9983 6985 10009 6991
rect 9983 6953 10009 6959
rect 10207 6929 10233 6935
rect 11265 6903 11271 6929
rect 11297 6903 11303 6929
rect 10207 6897 10233 6903
rect 9759 6873 9785 6879
rect 9759 6841 9785 6847
rect 10263 6873 10289 6879
rect 10369 6847 10375 6873
rect 10401 6847 10407 6873
rect 10929 6847 10935 6873
rect 10961 6847 10967 6873
rect 10263 6841 10289 6847
rect 9255 6817 9281 6823
rect 9255 6785 9281 6791
rect 9815 6817 9841 6823
rect 12671 6817 12697 6823
rect 12329 6791 12335 6817
rect 12361 6791 12367 6817
rect 9815 6785 9841 6791
rect 12671 6785 12697 6791
rect 8863 6761 8889 6767
rect 8863 6729 8889 6735
rect 9031 6761 9057 6767
rect 9031 6729 9057 6735
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 12503 6537 12529 6543
rect 7681 6511 7687 6537
rect 7713 6511 7719 6537
rect 8745 6511 8751 6537
rect 8777 6511 8783 6537
rect 10369 6511 10375 6537
rect 10401 6511 10407 6537
rect 11153 6511 11159 6537
rect 11185 6511 11191 6537
rect 12217 6511 12223 6537
rect 12249 6511 12255 6537
rect 12503 6505 12529 6511
rect 7345 6455 7351 6481
rect 7377 6455 7383 6481
rect 8913 6455 8919 6481
rect 8945 6455 8951 6481
rect 10817 6455 10823 6481
rect 10849 6455 10855 6481
rect 9305 6399 9311 6425
rect 9337 6399 9343 6425
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 8807 6201 8833 6207
rect 8807 6169 8833 6175
rect 9087 6201 9113 6207
rect 9087 6169 9113 6175
rect 9143 6089 9169 6095
rect 8969 6063 8975 6089
rect 9001 6063 9007 6089
rect 9143 6057 9169 6063
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 9529 2143 9535 2169
rect 9561 2143 9567 2169
rect 12609 2143 12615 2169
rect 12641 2143 12647 2169
rect 10039 2057 10065 2063
rect 10039 2025 10065 2031
rect 13119 2057 13145 2063
rect 13119 2025 13145 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 9311 1833 9337 1839
rect 9311 1801 9337 1807
rect 11047 1833 11073 1839
rect 11047 1801 11073 1807
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 8801 1751 8807 1777
rect 8833 1751 8839 1777
rect 10537 1751 10543 1777
rect 10569 1751 10575 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 7519 1665 7545 1671
rect 7519 1633 7545 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 8975 19111 9001 19137
rect 11215 19111 11241 19137
rect 12783 19111 12809 19137
rect 14687 19111 14713 19137
rect 8471 18999 8497 19025
rect 10823 18999 10849 19025
rect 12279 18999 12305 19025
rect 14295 18999 14321 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 11047 18719 11073 18745
rect 13119 18719 13145 18745
rect 10543 18607 10569 18633
rect 12727 18607 12753 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 11159 18327 11185 18353
rect 13399 18327 13425 18353
rect 10655 18215 10681 18241
rect 12895 18215 12921 18241
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 11943 14015 11969 14041
rect 11999 13903 12025 13929
rect 11943 13791 11969 13817
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 10375 13567 10401 13593
rect 12335 13567 12361 13593
rect 8919 13511 8945 13537
rect 10935 13511 10961 13537
rect 12559 13511 12585 13537
rect 12727 13511 12753 13537
rect 9311 13455 9337 13481
rect 11271 13455 11297 13481
rect 12895 13455 12921 13481
rect 13231 13455 13257 13481
rect 8751 13399 8777 13425
rect 13063 13399 13089 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 8079 13231 8105 13257
rect 10375 13231 10401 13257
rect 11327 13231 11353 13257
rect 11943 13231 11969 13257
rect 13175 13231 13201 13257
rect 11439 13175 11465 13201
rect 11495 13175 11521 13201
rect 12671 13175 12697 13201
rect 12727 13175 12753 13201
rect 6455 13119 6481 13145
rect 8135 13119 8161 13145
rect 8695 13119 8721 13145
rect 10319 13119 10345 13145
rect 11999 13119 12025 13145
rect 12559 13119 12585 13145
rect 18831 13119 18857 13145
rect 6791 13063 6817 13089
rect 7855 13063 7881 13089
rect 8359 13063 8385 13089
rect 9087 13063 9113 13089
rect 10151 13063 10177 13089
rect 10655 13063 10681 13089
rect 8079 13007 8105 13033
rect 10375 13007 10401 13033
rect 11943 13007 11969 13033
rect 20007 13007 20033 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 967 12783 993 12809
rect 7127 12783 7153 12809
rect 9759 12783 9785 12809
rect 11887 12783 11913 12809
rect 13007 12783 13033 12809
rect 2143 12727 2169 12753
rect 7407 12727 7433 12753
rect 9535 12727 9561 12753
rect 10039 12727 10065 12753
rect 11551 12727 11577 12753
rect 13231 12727 13257 12753
rect 13399 12727 13425 12753
rect 6175 12671 6201 12697
rect 6231 12671 6257 12697
rect 8135 12671 8161 12697
rect 8639 12671 8665 12697
rect 9479 12671 9505 12697
rect 13287 12671 13313 12697
rect 13567 12671 13593 12697
rect 13623 12671 13649 12697
rect 6063 12615 6089 12641
rect 7071 12615 7097 12641
rect 7183 12615 7209 12641
rect 8303 12615 8329 12641
rect 8471 12615 8497 12641
rect 9367 12615 9393 12641
rect 9703 12615 9729 12641
rect 9815 12615 9841 12641
rect 13455 12615 13481 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 13287 12391 13313 12417
rect 2143 12335 2169 12361
rect 6511 12335 6537 12361
rect 8415 12335 8441 12361
rect 9423 12335 9449 12361
rect 12951 12335 12977 12361
rect 5055 12279 5081 12305
rect 6119 12279 6145 12305
rect 6735 12279 6761 12305
rect 6959 12279 6985 12305
rect 8023 12279 8049 12305
rect 8751 12279 8777 12305
rect 9199 12279 9225 12305
rect 9759 12279 9785 12305
rect 10823 12279 10849 12305
rect 14351 12279 14377 12305
rect 14575 12279 14601 12305
rect 967 12223 993 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 8023 12055 8049 12081
rect 8247 12055 8273 12081
rect 9367 12055 9393 12081
rect 9423 12055 9449 12081
rect 6399 11999 6425 12025
rect 20007 11999 20033 12025
rect 6119 11943 6145 11969
rect 8527 11943 8553 11969
rect 8639 11943 8665 11969
rect 9647 11943 9673 11969
rect 9759 11943 9785 11969
rect 18831 11943 18857 11969
rect 8023 11887 8049 11913
rect 8079 11887 8105 11913
rect 8359 11887 8385 11913
rect 9479 11887 9505 11913
rect 9983 11887 10009 11913
rect 10039 11887 10065 11913
rect 6343 11831 6369 11857
rect 6455 11831 6481 11857
rect 7295 11831 7321 11857
rect 7463 11831 7489 11857
rect 8695 11831 8721 11857
rect 10151 11831 10177 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 9983 11663 10009 11689
rect 6567 11607 6593 11633
rect 6623 11607 6649 11633
rect 8303 11607 8329 11633
rect 20119 11607 20145 11633
rect 2143 11551 2169 11577
rect 6287 11551 6313 11577
rect 8247 11551 8273 11577
rect 9927 11551 9953 11577
rect 10039 11551 10065 11577
rect 10151 11551 10177 11577
rect 10935 11551 10961 11577
rect 12671 11551 12697 11577
rect 12951 11551 12977 11577
rect 14575 11551 14601 11577
rect 4831 11495 4857 11521
rect 5895 11495 5921 11521
rect 6847 11495 6873 11521
rect 11271 11495 11297 11521
rect 12335 11495 12361 11521
rect 13287 11495 13313 11521
rect 14351 11495 14377 11521
rect 967 11439 993 11465
rect 6567 11439 6593 11465
rect 8303 11439 8329 11465
rect 10263 11439 10289 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 11103 11271 11129 11297
rect 12223 11271 12249 11297
rect 5951 11215 5977 11241
rect 8527 11215 8553 11241
rect 13007 11215 13033 11241
rect 13455 11215 13481 11241
rect 20007 11215 20033 11241
rect 8079 11159 8105 11185
rect 8415 11159 8441 11185
rect 8695 11159 8721 11185
rect 10711 11159 10737 11185
rect 10823 11159 10849 11185
rect 10991 11159 11017 11185
rect 11999 11159 12025 11185
rect 12391 11159 12417 11185
rect 13063 11159 13089 11185
rect 13287 11159 13313 11185
rect 13343 11159 13369 11185
rect 18831 11159 18857 11185
rect 5783 11103 5809 11129
rect 6903 11103 6929 11129
rect 8751 11103 8777 11129
rect 11551 11103 11577 11129
rect 11831 11103 11857 11129
rect 12055 11103 12081 11129
rect 12167 11103 12193 11129
rect 12503 11103 12529 11129
rect 13623 11103 13649 11129
rect 5895 11047 5921 11073
rect 6007 11047 6033 11073
rect 6735 11047 6761 11073
rect 6847 11047 6873 11073
rect 7911 11047 7937 11073
rect 8247 11047 8273 11073
rect 10655 11047 10681 11073
rect 12279 11047 12305 11073
rect 12951 11047 12977 11073
rect 13511 11047 13537 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 10375 10879 10401 10905
rect 10823 10879 10849 10905
rect 10935 10879 10961 10905
rect 13287 10879 13313 10905
rect 14183 10879 14209 10905
rect 6679 10823 6705 10849
rect 8863 10823 8889 10849
rect 10487 10823 10513 10849
rect 11383 10823 11409 10849
rect 11551 10823 11577 10849
rect 12055 10823 12081 10849
rect 12615 10823 12641 10849
rect 12839 10823 12865 10849
rect 13679 10823 13705 10849
rect 14351 10823 14377 10849
rect 14407 10823 14433 10849
rect 6343 10767 6369 10793
rect 8695 10767 8721 10793
rect 10543 10767 10569 10793
rect 10655 10767 10681 10793
rect 11271 10767 11297 10793
rect 11495 10767 11521 10793
rect 11831 10767 11857 10793
rect 11943 10767 11969 10793
rect 12727 10767 12753 10793
rect 13175 10767 13201 10793
rect 13399 10767 13425 10793
rect 13511 10767 13537 10793
rect 13791 10767 13817 10793
rect 14015 10767 14041 10793
rect 14519 10767 14545 10793
rect 18831 10767 18857 10793
rect 7743 10711 7769 10737
rect 7967 10711 7993 10737
rect 9143 10711 9169 10737
rect 9759 10711 9785 10737
rect 10879 10711 10905 10737
rect 11663 10711 11689 10737
rect 11887 10711 11913 10737
rect 12783 10711 12809 10737
rect 13343 10711 13369 10737
rect 9255 10655 9281 10681
rect 9367 10655 9393 10681
rect 9591 10655 9617 10681
rect 20007 10655 20033 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 10767 10487 10793 10513
rect 12895 10431 12921 10457
rect 10039 10375 10065 10401
rect 10655 10375 10681 10401
rect 11775 10375 11801 10401
rect 7967 10319 7993 10345
rect 10935 10263 10961 10289
rect 11103 10263 11129 10289
rect 11271 10263 11297 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 12839 10095 12865 10121
rect 8079 10039 8105 10065
rect 8247 10039 8273 10065
rect 8415 10039 8441 10065
rect 8975 10039 9001 10065
rect 9367 10039 9393 10065
rect 11719 10039 11745 10065
rect 12895 10039 12921 10065
rect 5503 9983 5529 10009
rect 5839 9983 5865 10009
rect 7911 9983 7937 10009
rect 8695 9983 8721 10009
rect 9255 9983 9281 10009
rect 9759 9983 9785 10009
rect 12671 9983 12697 10009
rect 13007 9983 13033 10009
rect 13343 9983 13369 10009
rect 13735 9983 13761 10009
rect 6903 9927 6929 9953
rect 7127 9927 7153 9953
rect 14799 9927 14825 9953
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 8863 9703 8889 9729
rect 12503 9703 12529 9729
rect 7855 9647 7881 9673
rect 8303 9647 8329 9673
rect 8751 9647 8777 9673
rect 12447 9647 12473 9673
rect 7407 9591 7433 9617
rect 7743 9591 7769 9617
rect 7911 9591 7937 9617
rect 9535 9591 9561 9617
rect 9703 9591 9729 9617
rect 9871 9591 9897 9617
rect 10207 9591 10233 9617
rect 10823 9591 10849 9617
rect 11607 9591 11633 9617
rect 11775 9591 11801 9617
rect 11943 9591 11969 9617
rect 12335 9591 12361 9617
rect 13287 9591 13313 9617
rect 7575 9535 7601 9561
rect 9199 9535 9225 9561
rect 9591 9535 9617 9561
rect 9983 9535 10009 9561
rect 10711 9535 10737 9561
rect 11159 9535 11185 9561
rect 11327 9535 11353 9561
rect 11887 9535 11913 9561
rect 13063 9535 13089 9561
rect 13119 9535 13145 9561
rect 8079 9479 8105 9505
rect 9031 9479 9057 9505
rect 9367 9479 9393 9505
rect 10319 9479 10345 9505
rect 11551 9479 11577 9505
rect 12167 9479 12193 9505
rect 12951 9479 12977 9505
rect 13007 9479 13033 9505
rect 13567 9479 13593 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 8863 9311 8889 9337
rect 10095 9311 10121 9337
rect 11943 9311 11969 9337
rect 10767 9255 10793 9281
rect 10823 9255 10849 9281
rect 11607 9255 11633 9281
rect 11775 9255 11801 9281
rect 5727 9199 5753 9225
rect 7519 9199 7545 9225
rect 8751 9199 8777 9225
rect 9143 9199 9169 9225
rect 9255 9199 9281 9225
rect 9591 9199 9617 9225
rect 9927 9199 9953 9225
rect 10487 9199 10513 9225
rect 10655 9199 10681 9225
rect 11439 9199 11465 9225
rect 13119 9199 13145 9225
rect 18831 9199 18857 9225
rect 6119 9143 6145 9169
rect 7183 9143 7209 9169
rect 7407 9143 7433 9169
rect 7743 9143 7769 9169
rect 10991 9143 11017 9169
rect 13511 9143 13537 9169
rect 14575 9143 14601 9169
rect 14799 9143 14825 9169
rect 7351 9087 7377 9113
rect 9703 9087 9729 9113
rect 10543 9087 10569 9113
rect 11047 9087 11073 9113
rect 20007 9087 20033 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 9143 8919 9169 8945
rect 967 8863 993 8889
rect 6287 8863 6313 8889
rect 9311 8863 9337 8889
rect 12391 8863 12417 8889
rect 13175 8863 13201 8889
rect 13399 8863 13425 8889
rect 20007 8863 20033 8889
rect 2143 8807 2169 8833
rect 6735 8807 6761 8833
rect 6847 8807 6873 8833
rect 7631 8807 7657 8833
rect 8471 8807 8497 8833
rect 8919 8807 8945 8833
rect 9479 8807 9505 8833
rect 12783 8807 12809 8833
rect 13119 8807 13145 8833
rect 13455 8807 13481 8833
rect 13623 8807 13649 8833
rect 18831 8807 18857 8833
rect 6343 8751 6369 8777
rect 6455 8751 6481 8777
rect 7015 8751 7041 8777
rect 7351 8751 7377 8777
rect 8527 8751 8553 8777
rect 8751 8751 8777 8777
rect 9255 8751 9281 8777
rect 12223 8751 12249 8777
rect 12335 8751 12361 8777
rect 12895 8751 12921 8777
rect 12951 8751 12977 8777
rect 6903 8695 6929 8721
rect 7295 8695 7321 8721
rect 7407 8695 7433 8721
rect 8639 8695 8665 8721
rect 9647 8695 9673 8721
rect 13399 8695 13425 8721
rect 13567 8695 13593 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7407 8527 7433 8553
rect 10599 8527 10625 8553
rect 6119 8471 6145 8497
rect 9087 8471 9113 8497
rect 9199 8471 9225 8497
rect 10711 8471 10737 8497
rect 11271 8471 11297 8497
rect 13287 8471 13313 8497
rect 5727 8415 5753 8441
rect 9479 8415 9505 8441
rect 10935 8415 10961 8441
rect 11047 8415 11073 8441
rect 11103 8415 11129 8441
rect 12951 8415 12977 8441
rect 7183 8359 7209 8385
rect 9143 8359 9169 8385
rect 9311 8359 9337 8385
rect 10655 8359 10681 8385
rect 11215 8359 11241 8385
rect 14351 8359 14377 8385
rect 14575 8359 14601 8385
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 10823 8135 10849 8161
rect 10935 8135 10961 8161
rect 11047 8079 11073 8105
rect 20007 8079 20033 8105
rect 8807 8023 8833 8049
rect 8975 8023 9001 8049
rect 9031 8023 9057 8049
rect 9143 8023 9169 8049
rect 9367 8023 9393 8049
rect 9647 8023 9673 8049
rect 9871 8023 9897 8049
rect 10207 8023 10233 8049
rect 13007 8023 13033 8049
rect 13175 8023 13201 8049
rect 13623 8023 13649 8049
rect 13791 8023 13817 8049
rect 14071 8023 14097 8049
rect 18831 8023 18857 8049
rect 13287 7967 13313 7993
rect 13735 7967 13761 7993
rect 8863 7911 8889 7937
rect 9423 7911 9449 7937
rect 9479 7911 9505 7937
rect 10095 7911 10121 7937
rect 10151 7911 10177 7937
rect 11159 7911 11185 7937
rect 11215 7911 11241 7937
rect 11271 7911 11297 7937
rect 13175 7911 13201 7937
rect 13903 7911 13929 7937
rect 14015 7911 14041 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 8975 7743 9001 7769
rect 9311 7743 9337 7769
rect 11383 7743 11409 7769
rect 14407 7743 14433 7769
rect 6567 7687 6593 7713
rect 9815 7687 9841 7713
rect 13119 7687 13145 7713
rect 6175 7631 6201 7657
rect 8751 7631 8777 7657
rect 9087 7631 9113 7657
rect 9423 7631 9449 7657
rect 9647 7631 9673 7657
rect 11159 7631 11185 7657
rect 11327 7631 11353 7657
rect 11495 7631 11521 7657
rect 12727 7631 12753 7657
rect 7631 7575 7657 7601
rect 7855 7575 7881 7601
rect 8695 7575 8721 7601
rect 11439 7575 11465 7601
rect 14183 7575 14209 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 8191 7295 8217 7321
rect 9255 7295 9281 7321
rect 11551 7295 11577 7321
rect 11887 7295 11913 7321
rect 7855 7239 7881 7265
rect 11663 7239 11689 7265
rect 11999 7239 12025 7265
rect 11495 7183 11521 7209
rect 11831 7183 11857 7209
rect 9479 7127 9505 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 8919 6959 8945 6985
rect 9871 6959 9897 6985
rect 9983 6959 10009 6985
rect 10207 6903 10233 6929
rect 11271 6903 11297 6929
rect 9759 6847 9785 6873
rect 10263 6847 10289 6873
rect 10375 6847 10401 6873
rect 10935 6847 10961 6873
rect 9255 6791 9281 6817
rect 9815 6791 9841 6817
rect 12335 6791 12361 6817
rect 12671 6791 12697 6817
rect 8863 6735 8889 6761
rect 9031 6735 9057 6761
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 7687 6511 7713 6537
rect 8751 6511 8777 6537
rect 10375 6511 10401 6537
rect 11159 6511 11185 6537
rect 12223 6511 12249 6537
rect 12503 6511 12529 6537
rect 7351 6455 7377 6481
rect 8919 6455 8945 6481
rect 10823 6455 10849 6481
rect 9311 6399 9337 6425
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 8807 6175 8833 6201
rect 9087 6175 9113 6201
rect 8975 6063 9001 6089
rect 9143 6063 9169 6089
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 9535 2143 9561 2169
rect 12615 2143 12641 2169
rect 10039 2031 10065 2057
rect 13119 2031 13145 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 9311 1807 9337 1833
rect 11047 1807 11073 1833
rect 12783 1807 12809 1833
rect 8807 1751 8833 1777
rect 10543 1751 10569 1777
rect 12279 1751 12305 1777
rect 7519 1639 7545 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 7728 20600 7784 21000
rect 10080 20600 10136 21000
rect 10416 20600 10472 21000
rect 10752 20600 10808 21000
rect 12096 20600 12152 21000
rect 12432 20600 12488 21000
rect 12768 20600 12824 21000
rect 13104 20600 13160 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 7742 19138 7770 20600
rect 7742 19105 7770 19110
rect 8974 19138 9002 19143
rect 8974 19091 9002 19110
rect 8470 19025 8498 19031
rect 8470 18999 8471 19025
rect 8497 18999 8498 19025
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 7854 13258 7882 13263
rect 2086 13146 2114 13151
rect 966 12809 994 12815
rect 966 12783 967 12809
rect 993 12783 994 12809
rect 966 12474 994 12783
rect 966 12441 994 12446
rect 966 12250 994 12255
rect 966 12203 994 12222
rect 966 11466 994 11471
rect 966 11419 994 11438
rect 2086 10738 2114 13118
rect 6454 13146 6482 13151
rect 6454 13145 6538 13146
rect 6454 13119 6455 13145
rect 6481 13119 6538 13145
rect 6454 13118 6538 13119
rect 6454 13113 6482 13118
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 2142 12754 2170 12759
rect 2142 12707 2170 12726
rect 5054 12754 5082 12759
rect 2142 12362 2170 12367
rect 2142 12315 2170 12334
rect 5054 12305 5082 12726
rect 6174 12754 6202 12759
rect 6174 12697 6202 12726
rect 6174 12671 6175 12697
rect 6201 12671 6202 12697
rect 6174 12665 6202 12671
rect 6230 12698 6258 12703
rect 6230 12651 6258 12670
rect 6454 12698 6482 12703
rect 5054 12279 5055 12305
rect 5081 12279 5082 12305
rect 5054 12273 5082 12279
rect 6062 12641 6090 12647
rect 6062 12615 6063 12641
rect 6089 12615 6090 12641
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 6062 11970 6090 12615
rect 6118 12306 6146 12311
rect 6118 12305 6426 12306
rect 6118 12279 6119 12305
rect 6145 12279 6426 12305
rect 6118 12278 6426 12279
rect 6118 12273 6146 12278
rect 6398 12025 6426 12278
rect 6454 12250 6482 12670
rect 6510 12361 6538 13118
rect 6790 13090 6818 13095
rect 6790 13089 7154 13090
rect 6790 13063 6791 13089
rect 6817 13063 7154 13089
rect 6790 13062 7154 13063
rect 6790 13057 6818 13062
rect 7126 12809 7154 13062
rect 7854 13089 7882 13230
rect 8078 13258 8106 13263
rect 8078 13211 8106 13230
rect 8470 13258 8498 18999
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 10094 18354 10122 20600
rect 10430 18746 10458 20600
rect 10766 19138 10794 20600
rect 10766 19105 10794 19110
rect 11214 19138 11242 19143
rect 11214 19091 11242 19110
rect 12110 19138 12138 20600
rect 12110 19105 12138 19110
rect 10430 18713 10458 18718
rect 10822 19025 10850 19031
rect 10822 18999 10823 19025
rect 10849 18999 10850 19025
rect 10094 18321 10122 18326
rect 10542 18633 10570 18639
rect 10542 18607 10543 18633
rect 10569 18607 10570 18633
rect 10150 18242 10178 18247
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 8918 13537 8946 13543
rect 8918 13511 8919 13537
rect 8945 13511 8946 13537
rect 8470 13225 8498 13230
rect 8750 13426 8778 13431
rect 8918 13426 8946 13511
rect 9310 13482 9338 13487
rect 9310 13481 9786 13482
rect 9310 13455 9311 13481
rect 9337 13455 9786 13481
rect 9310 13454 9786 13455
rect 9310 13449 9338 13454
rect 8750 13425 8946 13426
rect 8750 13399 8751 13425
rect 8777 13399 8946 13425
rect 8750 13398 8946 13399
rect 8134 13146 8162 13151
rect 8134 13099 8162 13118
rect 8638 13146 8666 13151
rect 7854 13063 7855 13089
rect 7881 13063 7882 13089
rect 7854 13057 7882 13063
rect 8358 13090 8386 13095
rect 8358 13089 8442 13090
rect 8358 13063 8359 13089
rect 8385 13063 8442 13089
rect 8358 13062 8442 13063
rect 8358 13057 8386 13062
rect 7126 12783 7127 12809
rect 7153 12783 7154 12809
rect 7126 12777 7154 12783
rect 7406 13034 7434 13039
rect 7406 12753 7434 13006
rect 8078 13034 8106 13039
rect 8078 12987 8106 13006
rect 7406 12727 7407 12753
rect 7433 12727 7434 12753
rect 7406 12721 7434 12727
rect 8134 12754 8162 12759
rect 8134 12697 8162 12726
rect 8134 12671 8135 12697
rect 8161 12671 8162 12697
rect 8134 12665 8162 12671
rect 7070 12641 7098 12647
rect 7070 12615 7071 12641
rect 7097 12615 7098 12641
rect 6510 12335 6511 12361
rect 6537 12335 6538 12361
rect 6510 12306 6538 12335
rect 6958 12362 6986 12367
rect 6734 12306 6762 12311
rect 6510 12305 6762 12306
rect 6510 12279 6735 12305
rect 6761 12279 6762 12305
rect 6510 12278 6762 12279
rect 6454 12222 6650 12250
rect 6398 11999 6399 12025
rect 6425 11999 6426 12025
rect 6398 11993 6426 11999
rect 6118 11970 6146 11975
rect 6062 11969 6146 11970
rect 6062 11943 6119 11969
rect 6145 11943 6146 11969
rect 6062 11942 6146 11943
rect 6118 11937 6146 11942
rect 6342 11858 6370 11863
rect 4830 11634 4858 11639
rect 2142 11578 2170 11583
rect 2142 11531 2170 11550
rect 4830 11521 4858 11606
rect 6286 11577 6314 11583
rect 6286 11551 6287 11577
rect 6313 11551 6314 11577
rect 4830 11495 4831 11521
rect 4857 11495 4858 11521
rect 4830 11489 4858 11495
rect 5894 11521 5922 11527
rect 5894 11495 5895 11521
rect 5921 11495 5922 11521
rect 5782 11466 5810 11471
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 5782 11129 5810 11438
rect 5894 11242 5922 11495
rect 5950 11242 5978 11247
rect 5894 11241 5978 11242
rect 5894 11215 5951 11241
rect 5977 11215 5978 11241
rect 5894 11214 5978 11215
rect 5950 11209 5978 11214
rect 5782 11103 5783 11129
rect 5809 11103 5810 11129
rect 5782 11097 5810 11103
rect 2086 10705 2114 10710
rect 5894 11073 5922 11079
rect 5894 11047 5895 11073
rect 5921 11047 5922 11073
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 5502 10010 5530 10015
rect 5838 10010 5866 10015
rect 5894 10010 5922 11047
rect 6006 11074 6034 11079
rect 6006 11027 6034 11046
rect 6286 10962 6314 11551
rect 6342 11074 6370 11830
rect 6454 11857 6482 11863
rect 6454 11831 6455 11857
rect 6481 11831 6482 11857
rect 6454 11130 6482 11831
rect 6566 11634 6594 11639
rect 6566 11587 6594 11606
rect 6622 11633 6650 12222
rect 6622 11607 6623 11633
rect 6649 11607 6650 11633
rect 6622 11601 6650 11607
rect 6734 11522 6762 12278
rect 6958 12305 6986 12334
rect 6958 12279 6959 12305
rect 6985 12279 6986 12305
rect 6958 12273 6986 12279
rect 7070 11858 7098 12615
rect 7070 11825 7098 11830
rect 7182 12641 7210 12647
rect 7182 12615 7183 12641
rect 7209 12615 7210 12641
rect 6846 11522 6874 11527
rect 6734 11521 6874 11522
rect 6734 11495 6847 11521
rect 6873 11495 6874 11521
rect 6734 11494 6874 11495
rect 6566 11466 6594 11471
rect 6846 11466 6874 11494
rect 6846 11438 6986 11466
rect 6566 11419 6594 11438
rect 6454 11097 6482 11102
rect 6902 11130 6930 11135
rect 6902 11083 6930 11102
rect 6734 11074 6762 11079
rect 6342 11041 6370 11046
rect 6678 11073 6762 11074
rect 6678 11047 6735 11073
rect 6761 11047 6762 11073
rect 6678 11046 6762 11047
rect 6342 10962 6370 10967
rect 6286 10934 6342 10962
rect 6342 10793 6370 10934
rect 6678 10849 6706 11046
rect 6734 11041 6762 11046
rect 6790 11074 6818 11079
rect 6678 10823 6679 10849
rect 6705 10823 6706 10849
rect 6678 10817 6706 10823
rect 6342 10767 6343 10793
rect 6369 10767 6370 10793
rect 6342 10761 6370 10767
rect 5502 10009 5754 10010
rect 5502 9983 5503 10009
rect 5529 9983 5754 10009
rect 5502 9982 5754 9983
rect 5502 9977 5530 9982
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 5726 9226 5754 9982
rect 5838 10009 5922 10010
rect 5838 9983 5839 10009
rect 5865 9983 5922 10009
rect 5838 9982 5922 9983
rect 5838 9977 5866 9982
rect 5894 9954 5922 9982
rect 5894 9921 5922 9926
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 966 8889 994 8895
rect 966 8863 967 8889
rect 993 8863 994 8889
rect 966 8442 994 8863
rect 2142 8834 2170 8839
rect 2142 8787 2170 8806
rect 966 8409 994 8414
rect 5726 8442 5754 9198
rect 6118 9170 6146 9175
rect 6118 9123 6146 9142
rect 6286 8890 6314 8895
rect 6118 8889 6314 8890
rect 6118 8863 6287 8889
rect 6313 8863 6314 8889
rect 6118 8862 6314 8863
rect 6118 8497 6146 8862
rect 6286 8857 6314 8862
rect 6342 8834 6370 8839
rect 6342 8777 6370 8806
rect 6734 8834 6762 8839
rect 6790 8834 6818 11046
rect 6846 11073 6874 11079
rect 6846 11047 6847 11073
rect 6873 11047 6874 11073
rect 6846 11018 6874 11047
rect 6846 10985 6874 10990
rect 6958 10962 6986 11438
rect 7182 11018 7210 12615
rect 8302 12642 8330 12647
rect 8358 12642 8386 12647
rect 8302 12641 8358 12642
rect 8302 12615 8303 12641
rect 8329 12615 8358 12641
rect 8302 12614 8358 12615
rect 8302 12609 8330 12614
rect 7910 12362 7938 12367
rect 7938 12334 7994 12362
rect 7910 12329 7938 12334
rect 7966 11914 7994 12334
rect 8022 12305 8050 12311
rect 8022 12279 8023 12305
rect 8049 12279 8050 12305
rect 8022 12194 8050 12279
rect 8022 12161 8050 12166
rect 8022 12082 8050 12087
rect 8246 12082 8274 12087
rect 8022 12081 8274 12082
rect 8022 12055 8023 12081
rect 8049 12055 8247 12081
rect 8273 12055 8274 12081
rect 8022 12054 8274 12055
rect 8022 12049 8050 12054
rect 8246 12049 8274 12054
rect 8358 12026 8386 12614
rect 8414 12362 8442 13062
rect 8638 12697 8666 13118
rect 8638 12671 8639 12697
rect 8665 12671 8666 12697
rect 8638 12665 8666 12671
rect 8694 13146 8722 13151
rect 8750 13146 8778 13398
rect 8694 13145 8778 13146
rect 8694 13119 8695 13145
rect 8721 13119 8778 13145
rect 8694 13118 8778 13119
rect 9534 13146 9562 13151
rect 8470 12642 8498 12647
rect 8470 12595 8498 12614
rect 8414 12361 8498 12362
rect 8414 12335 8415 12361
rect 8441 12335 8498 12361
rect 8414 12334 8498 12335
rect 8414 12329 8442 12334
rect 8302 11998 8386 12026
rect 8470 12306 8498 12334
rect 8694 12306 8722 13118
rect 9086 13089 9114 13095
rect 9086 13063 9087 13089
rect 9113 13063 9114 13089
rect 8750 12306 8778 12311
rect 8470 12278 8750 12306
rect 8302 11970 8330 11998
rect 8190 11942 8330 11970
rect 8022 11914 8050 11919
rect 7966 11913 8050 11914
rect 7966 11887 8023 11913
rect 8049 11887 8050 11913
rect 7966 11886 8050 11887
rect 8022 11881 8050 11886
rect 8078 11914 8106 11919
rect 8190 11914 8218 11942
rect 8078 11913 8218 11914
rect 8078 11887 8079 11913
rect 8105 11887 8218 11913
rect 8078 11886 8218 11887
rect 8358 11914 8386 11919
rect 8078 11881 8106 11886
rect 7294 11858 7322 11863
rect 7294 11811 7322 11830
rect 7462 11858 7490 11863
rect 7462 11811 7490 11830
rect 8078 11186 8106 11191
rect 8078 11139 8106 11158
rect 7910 11074 7938 11079
rect 7182 10985 7210 10990
rect 7798 11046 7910 11074
rect 8134 11074 8162 11886
rect 8358 11867 8386 11886
rect 8302 11858 8330 11863
rect 8302 11746 8330 11830
rect 8302 11718 8386 11746
rect 8302 11633 8330 11639
rect 8302 11607 8303 11633
rect 8329 11607 8330 11633
rect 8246 11577 8274 11583
rect 8246 11551 8247 11577
rect 8273 11551 8274 11577
rect 8246 11186 8274 11551
rect 8302 11578 8330 11607
rect 8302 11545 8330 11550
rect 8302 11466 8330 11471
rect 8358 11466 8386 11718
rect 8302 11465 8386 11466
rect 8302 11439 8303 11465
rect 8329 11439 8386 11465
rect 8302 11438 8386 11439
rect 8302 11433 8330 11438
rect 8246 11153 8274 11158
rect 8302 11354 8330 11359
rect 8246 11074 8274 11079
rect 8134 11073 8274 11074
rect 8134 11047 8247 11073
rect 8273 11047 8274 11073
rect 8134 11046 8274 11047
rect 6958 10929 6986 10934
rect 7742 10794 7770 10799
rect 7742 10737 7770 10766
rect 7742 10711 7743 10737
rect 7769 10711 7770 10737
rect 7742 10705 7770 10711
rect 6902 9953 6930 9959
rect 6902 9927 6903 9953
rect 6929 9927 6930 9953
rect 6902 9730 6930 9927
rect 6902 9697 6930 9702
rect 7126 9953 7154 9959
rect 7126 9927 7127 9953
rect 7153 9927 7154 9953
rect 7126 9226 7154 9927
rect 7406 9618 7434 9623
rect 7126 9193 7154 9198
rect 7182 9590 7406 9618
rect 6902 9170 6930 9175
rect 6846 8834 6874 8839
rect 6790 8833 6874 8834
rect 6790 8807 6847 8833
rect 6873 8807 6874 8833
rect 6790 8806 6874 8807
rect 6734 8787 6762 8806
rect 6846 8801 6874 8806
rect 6342 8751 6343 8777
rect 6369 8751 6370 8777
rect 6342 8745 6370 8751
rect 6454 8778 6482 8783
rect 6454 8731 6482 8750
rect 6902 8721 6930 9142
rect 7182 9169 7210 9590
rect 7406 9571 7434 9590
rect 7742 9618 7770 9623
rect 7742 9571 7770 9590
rect 7574 9562 7602 9567
rect 7574 9515 7602 9534
rect 7462 9226 7490 9231
rect 7182 9143 7183 9169
rect 7209 9143 7210 9169
rect 7182 9137 7210 9143
rect 7406 9169 7434 9175
rect 7406 9143 7407 9169
rect 7433 9143 7434 9169
rect 7350 9114 7378 9119
rect 7238 9113 7378 9114
rect 7238 9087 7351 9113
rect 7377 9087 7378 9113
rect 7238 9086 7378 9087
rect 6902 8695 6903 8721
rect 6929 8695 6930 8721
rect 6902 8689 6930 8695
rect 7014 8777 7042 8783
rect 7014 8751 7015 8777
rect 7041 8751 7042 8777
rect 7014 8666 7042 8751
rect 7014 8633 7042 8638
rect 7070 8722 7098 8727
rect 6118 8471 6119 8497
rect 6145 8471 6146 8497
rect 6118 8465 6146 8471
rect 5726 8395 5754 8414
rect 6174 8386 6202 8391
rect 7070 8386 7098 8694
rect 7238 8666 7266 9086
rect 7350 9081 7378 9086
rect 7406 8834 7434 9143
rect 7406 8801 7434 8806
rect 7350 8778 7378 8783
rect 7350 8731 7378 8750
rect 7238 8633 7266 8638
rect 7294 8721 7322 8727
rect 7294 8695 7295 8721
rect 7321 8695 7322 8721
rect 7294 8442 7322 8695
rect 7406 8722 7434 8727
rect 7406 8675 7434 8694
rect 7406 8554 7434 8559
rect 7462 8554 7490 9198
rect 7518 9225 7546 9231
rect 7518 9199 7519 9225
rect 7545 9199 7546 9225
rect 7518 9170 7546 9199
rect 7518 9137 7546 9142
rect 7742 9226 7770 9231
rect 7742 9169 7770 9198
rect 7742 9143 7743 9169
rect 7769 9143 7770 9169
rect 7630 8946 7658 8951
rect 7630 8833 7658 8918
rect 7630 8807 7631 8833
rect 7657 8807 7658 8833
rect 7630 8801 7658 8807
rect 7406 8553 7490 8554
rect 7406 8527 7407 8553
rect 7433 8527 7490 8553
rect 7406 8526 7490 8527
rect 7406 8521 7434 8526
rect 7294 8409 7322 8414
rect 7182 8386 7210 8391
rect 7070 8385 7210 8386
rect 7070 8359 7183 8385
rect 7209 8359 7210 8385
rect 7070 8358 7210 8359
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 6174 7657 6202 8358
rect 7182 8353 7210 8358
rect 6566 7770 6594 7775
rect 6566 7713 6594 7742
rect 6566 7687 6567 7713
rect 6593 7687 6594 7713
rect 6566 7681 6594 7687
rect 6174 7631 6175 7657
rect 6201 7631 6202 7657
rect 6174 7625 6202 7631
rect 7630 7602 7658 7621
rect 7742 7602 7770 9143
rect 7798 8386 7826 11046
rect 7910 11027 7938 11046
rect 8246 11041 8274 11046
rect 7966 10962 7994 10967
rect 7966 10737 7994 10934
rect 7966 10711 7967 10737
rect 7993 10711 7994 10737
rect 7966 10345 7994 10711
rect 8246 10794 8274 10799
rect 7966 10319 7967 10345
rect 7993 10319 7994 10345
rect 7910 10009 7938 10015
rect 7910 9983 7911 10009
rect 7937 9983 7938 10009
rect 7854 9674 7882 9679
rect 7854 9627 7882 9646
rect 7910 9617 7938 9983
rect 7910 9591 7911 9617
rect 7937 9591 7938 9617
rect 7910 9114 7938 9591
rect 7966 9226 7994 10319
rect 8078 10570 8106 10575
rect 8078 10065 8106 10542
rect 8078 10039 8079 10065
rect 8105 10039 8106 10065
rect 8078 10033 8106 10039
rect 8246 10065 8274 10766
rect 8246 10039 8247 10065
rect 8273 10039 8274 10065
rect 8246 10033 8274 10039
rect 8302 9673 8330 11326
rect 8470 11298 8498 12278
rect 8750 12259 8778 12278
rect 8694 12194 8722 12199
rect 8526 11970 8554 11975
rect 8526 11923 8554 11942
rect 8638 11969 8666 11975
rect 8638 11943 8639 11969
rect 8665 11943 8666 11969
rect 8638 11858 8666 11943
rect 8638 11825 8666 11830
rect 8694 11857 8722 12166
rect 9086 12082 9114 13063
rect 9534 12754 9562 13118
rect 9758 12809 9786 13454
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 10150 13089 10178 18214
rect 10542 15974 10570 18607
rect 10654 18242 10682 18247
rect 10654 18195 10682 18214
rect 10374 15946 10570 15974
rect 10374 13593 10402 15946
rect 10374 13567 10375 13593
rect 10401 13567 10402 13593
rect 10374 13257 10402 13567
rect 10374 13231 10375 13257
rect 10401 13231 10402 13257
rect 10374 13225 10402 13231
rect 10318 13146 10346 13151
rect 10318 13099 10346 13118
rect 10150 13063 10151 13089
rect 10177 13063 10178 13089
rect 9758 12783 9759 12809
rect 9785 12783 9786 12809
rect 9758 12777 9786 12783
rect 10038 13034 10066 13039
rect 9534 12707 9562 12726
rect 10038 12753 10066 13006
rect 10038 12727 10039 12753
rect 10065 12727 10066 12753
rect 10038 12721 10066 12727
rect 9478 12698 9506 12703
rect 9478 12651 9506 12670
rect 10150 12698 10178 13063
rect 10654 13089 10682 13095
rect 10654 13063 10655 13089
rect 10681 13063 10682 13089
rect 10374 13034 10402 13039
rect 10374 12987 10402 13006
rect 10150 12665 10178 12670
rect 9366 12641 9394 12647
rect 9366 12615 9367 12641
rect 9393 12615 9394 12641
rect 9198 12306 9226 12311
rect 9198 12259 9226 12278
rect 9086 12049 9114 12054
rect 9366 12081 9394 12615
rect 9702 12641 9730 12647
rect 9702 12615 9703 12641
rect 9729 12615 9730 12641
rect 9702 12418 9730 12615
rect 9814 12641 9842 12647
rect 9814 12615 9815 12641
rect 9841 12615 9842 12641
rect 9814 12474 9842 12615
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9814 12446 10066 12474
rect 9702 12390 9842 12418
rect 9422 12361 9450 12367
rect 9422 12335 9423 12361
rect 9449 12335 9450 12361
rect 9422 12306 9450 12335
rect 9758 12306 9786 12311
rect 9422 12273 9450 12278
rect 9702 12305 9786 12306
rect 9702 12279 9759 12305
rect 9785 12279 9786 12305
rect 9702 12278 9786 12279
rect 9366 12055 9367 12081
rect 9393 12055 9394 12081
rect 9366 12049 9394 12055
rect 9422 12082 9450 12087
rect 9422 12035 9450 12054
rect 9646 11970 9674 11975
rect 8694 11831 8695 11857
rect 8721 11831 8722 11857
rect 8694 11825 8722 11831
rect 9478 11914 9506 11919
rect 8358 11270 8498 11298
rect 8526 11270 8834 11298
rect 8358 10962 8386 11270
rect 8526 11241 8554 11270
rect 8526 11215 8527 11241
rect 8553 11215 8554 11241
rect 8526 11209 8554 11215
rect 8414 11185 8442 11191
rect 8414 11159 8415 11185
rect 8441 11159 8442 11185
rect 8414 11074 8442 11159
rect 8694 11186 8722 11191
rect 8694 11139 8722 11158
rect 8750 11129 8778 11135
rect 8750 11103 8751 11129
rect 8777 11103 8778 11129
rect 8750 11074 8778 11103
rect 8414 11046 8778 11074
rect 8694 10962 8722 10967
rect 8358 10929 8386 10934
rect 8638 10934 8694 10962
rect 8414 10906 8442 10911
rect 8414 10178 8442 10878
rect 8414 10150 8498 10178
rect 8302 9647 8303 9673
rect 8329 9647 8330 9673
rect 7966 9193 7994 9198
rect 8078 9505 8106 9511
rect 8078 9479 8079 9505
rect 8105 9479 8106 9505
rect 8078 9114 8106 9479
rect 8302 9450 8330 9647
rect 8302 9417 8330 9422
rect 8414 10065 8442 10071
rect 8414 10039 8415 10065
rect 8441 10039 8442 10065
rect 7910 9086 8106 9114
rect 8414 9114 8442 10039
rect 7854 8386 7882 8391
rect 7798 8358 7854 8386
rect 7854 8353 7882 8358
rect 7854 7602 7882 7607
rect 7742 7601 7882 7602
rect 7742 7575 7855 7601
rect 7881 7575 7882 7601
rect 7742 7574 7882 7575
rect 7630 7569 7658 7574
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 7854 7265 7882 7574
rect 7910 7602 7938 9086
rect 8414 8834 8442 9086
rect 8470 9058 8498 10150
rect 8638 10010 8666 10934
rect 8694 10929 8722 10934
rect 8694 10794 8722 10799
rect 8694 10747 8722 10766
rect 8694 10010 8722 10015
rect 8638 10009 8722 10010
rect 8638 9983 8695 10009
rect 8721 9983 8722 10009
rect 8638 9982 8722 9983
rect 8694 9977 8722 9982
rect 8750 9898 8778 11046
rect 8806 10570 8834 11270
rect 9478 11242 9506 11886
rect 9478 10962 9506 11214
rect 9478 10929 9506 10934
rect 9590 11858 9618 11863
rect 8806 10537 8834 10542
rect 8862 10849 8890 10855
rect 8862 10823 8863 10849
rect 8889 10823 8890 10849
rect 8694 9870 8778 9898
rect 8862 10290 8890 10823
rect 9142 10737 9170 10743
rect 9142 10711 9143 10737
rect 9169 10711 9170 10737
rect 9142 10570 9170 10711
rect 9254 10682 9282 10687
rect 9142 10537 9170 10542
rect 9198 10681 9282 10682
rect 9198 10655 9255 10681
rect 9281 10655 9282 10681
rect 9198 10654 9282 10655
rect 8694 9562 8722 9870
rect 8694 9529 8722 9534
rect 8750 9730 8778 9735
rect 8750 9673 8778 9702
rect 8862 9729 8890 10262
rect 9198 10178 9226 10654
rect 9254 10649 9282 10654
rect 9366 10681 9394 10687
rect 9366 10655 9367 10681
rect 9393 10655 9394 10681
rect 9366 10290 9394 10655
rect 9590 10681 9618 11830
rect 9590 10655 9591 10681
rect 9617 10655 9618 10681
rect 9590 10514 9618 10655
rect 9590 10481 9618 10486
rect 9366 10257 9394 10262
rect 8974 10150 9226 10178
rect 8974 10066 9002 10150
rect 8862 9703 8863 9729
rect 8889 9703 8890 9729
rect 8862 9697 8890 9703
rect 8918 10065 9002 10066
rect 8918 10039 8975 10065
rect 9001 10039 9002 10065
rect 8918 10038 9002 10039
rect 8750 9647 8751 9673
rect 8777 9647 8778 9673
rect 8750 9225 8778 9647
rect 8750 9199 8751 9225
rect 8777 9199 8778 9225
rect 8750 9193 8778 9199
rect 8862 9338 8890 9343
rect 8918 9338 8946 10038
rect 8974 10033 9002 10038
rect 9366 10065 9394 10071
rect 9366 10039 9367 10065
rect 9393 10039 9394 10065
rect 9254 10009 9282 10015
rect 9254 9983 9255 10009
rect 9281 9983 9282 10009
rect 9198 9562 9226 9567
rect 9254 9562 9282 9983
rect 9366 9618 9394 10039
rect 9534 9618 9562 9623
rect 9366 9590 9534 9618
rect 9534 9571 9562 9590
rect 9226 9534 9282 9562
rect 9310 9562 9338 9567
rect 9198 9515 9226 9534
rect 9030 9506 9058 9511
rect 9030 9505 9170 9506
rect 9030 9479 9031 9505
rect 9057 9479 9170 9505
rect 9030 9478 9170 9479
rect 9030 9473 9058 9478
rect 8862 9337 9114 9338
rect 8862 9311 8863 9337
rect 8889 9311 9114 9337
rect 8862 9310 9114 9311
rect 8470 8946 8498 9030
rect 8694 9170 8722 9175
rect 8470 8918 8610 8946
rect 8470 8834 8498 8839
rect 8414 8833 8498 8834
rect 8414 8807 8471 8833
rect 8497 8807 8498 8833
rect 8414 8806 8498 8807
rect 8470 8801 8498 8806
rect 8526 8778 8554 8783
rect 8526 8731 8554 8750
rect 8582 8498 8610 8918
rect 8694 8778 8722 9142
rect 8750 8778 8778 8783
rect 8694 8777 8778 8778
rect 8694 8751 8751 8777
rect 8777 8751 8778 8777
rect 8694 8750 8778 8751
rect 8750 8745 8778 8750
rect 8862 8778 8890 9310
rect 9086 8946 9114 9310
rect 9142 9226 9170 9478
rect 9142 9179 9170 9198
rect 9254 9450 9282 9455
rect 9254 9225 9282 9422
rect 9254 9199 9255 9225
rect 9281 9199 9282 9225
rect 9254 9193 9282 9199
rect 9310 9002 9338 9534
rect 9590 9562 9618 9567
rect 9590 9515 9618 9534
rect 9366 9505 9394 9511
rect 9366 9479 9367 9505
rect 9393 9479 9394 9505
rect 9366 9338 9394 9479
rect 9366 9310 9562 9338
rect 9198 8974 9338 9002
rect 9478 9226 9506 9231
rect 9534 9226 9562 9310
rect 9590 9226 9618 9231
rect 9534 9198 9590 9226
rect 9142 8946 9170 8951
rect 9086 8945 9170 8946
rect 9086 8919 9143 8945
rect 9169 8919 9170 8945
rect 9086 8918 9170 8919
rect 9142 8913 9170 8918
rect 8918 8834 8946 8839
rect 8918 8787 8946 8806
rect 8862 8745 8890 8750
rect 8638 8722 8666 8727
rect 8638 8721 8722 8722
rect 8638 8695 8639 8721
rect 8665 8695 8722 8721
rect 8638 8694 8722 8695
rect 8638 8689 8666 8694
rect 8694 8554 8722 8694
rect 8694 8526 9114 8554
rect 8582 8470 8834 8498
rect 8806 8049 8834 8470
rect 9086 8497 9114 8526
rect 9086 8471 9087 8497
rect 9113 8471 9114 8497
rect 9086 8465 9114 8471
rect 9198 8498 9226 8974
rect 9310 8889 9338 8895
rect 9310 8863 9311 8889
rect 9337 8863 9338 8889
rect 9254 8834 9282 8839
rect 9254 8777 9282 8806
rect 9254 8751 9255 8777
rect 9281 8751 9282 8777
rect 9254 8745 9282 8751
rect 9310 8778 9338 8863
rect 9478 8833 9506 9198
rect 9478 8807 9479 8833
rect 9505 8807 9506 8833
rect 9478 8801 9506 8807
rect 9590 8834 9618 9198
rect 9646 9002 9674 11942
rect 9702 11746 9730 12278
rect 9758 12273 9786 12278
rect 9702 11713 9730 11718
rect 9758 11969 9786 11975
rect 9758 11943 9759 11969
rect 9785 11943 9786 11969
rect 9758 11074 9786 11943
rect 9814 11858 9842 12390
rect 9982 11913 10010 11919
rect 9982 11887 9983 11913
rect 10009 11887 10010 11913
rect 9982 11858 10010 11887
rect 9842 11830 10010 11858
rect 10038 11913 10066 12446
rect 10654 12306 10682 13063
rect 10654 12273 10682 12278
rect 10822 12305 10850 18999
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 11046 18746 11074 18751
rect 11046 18699 11074 18718
rect 11158 18354 11186 18359
rect 11158 18307 11186 18326
rect 12278 15974 12306 18999
rect 12446 18746 12474 20600
rect 12782 20538 12810 20600
rect 12782 20510 12922 20538
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 12446 18713 12474 18718
rect 11942 15946 12306 15974
rect 12726 18633 12754 18639
rect 12726 18607 12727 18633
rect 12753 18607 12754 18633
rect 11942 14042 11970 15946
rect 11942 14041 12362 14042
rect 11942 14015 11943 14041
rect 11969 14015 12362 14041
rect 11942 14014 12362 14015
rect 11942 14009 11970 14014
rect 11998 13929 12026 13935
rect 11998 13903 11999 13929
rect 12025 13903 12026 13929
rect 11494 13818 11522 13823
rect 11438 13790 11494 13818
rect 10934 13538 10962 13543
rect 10934 13491 10962 13510
rect 11270 13482 11298 13487
rect 11270 13481 11354 13482
rect 11270 13455 11271 13481
rect 11297 13455 11354 13481
rect 11270 13454 11354 13455
rect 11270 13449 11298 13454
rect 11326 13257 11354 13454
rect 11438 13454 11466 13790
rect 11494 13785 11522 13790
rect 11942 13818 11970 13823
rect 11942 13771 11970 13790
rect 11494 13538 11522 13543
rect 11522 13510 11578 13538
rect 11494 13505 11522 13510
rect 11438 13426 11522 13454
rect 11326 13231 11327 13257
rect 11353 13231 11354 13257
rect 11326 13225 11354 13231
rect 10822 12279 10823 12305
rect 10849 12279 10850 12305
rect 10822 12250 10850 12279
rect 11438 13201 11466 13207
rect 11438 13175 11439 13201
rect 11465 13175 11466 13201
rect 10822 12222 11018 12250
rect 10038 11887 10039 11913
rect 10065 11887 10066 11913
rect 10038 11858 10066 11887
rect 10038 11830 10122 11858
rect 9814 11825 9842 11830
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9870 11690 9898 11695
rect 9982 11690 10010 11695
rect 9898 11689 10010 11690
rect 9898 11663 9983 11689
rect 10009 11663 10010 11689
rect 9898 11662 10010 11663
rect 9870 11657 9898 11662
rect 9982 11657 10010 11662
rect 9926 11577 9954 11583
rect 9926 11551 9927 11577
rect 9953 11551 9954 11577
rect 9926 11186 9954 11551
rect 9926 11153 9954 11158
rect 10038 11577 10066 11583
rect 10038 11551 10039 11577
rect 10065 11551 10066 11577
rect 10038 11074 10066 11551
rect 9758 11046 10066 11074
rect 10094 11298 10122 11830
rect 10150 11857 10178 11863
rect 10150 11831 10151 11857
rect 10177 11831 10178 11857
rect 10150 11577 10178 11831
rect 10150 11551 10151 11577
rect 10177 11551 10178 11577
rect 10150 11545 10178 11551
rect 10934 11578 10962 11583
rect 10934 11531 10962 11550
rect 9758 10738 9786 10743
rect 9758 10009 9786 10710
rect 9758 9983 9759 10009
rect 9785 9983 9786 10009
rect 9758 9977 9786 9983
rect 9702 9618 9730 9623
rect 9814 9618 9842 11046
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 10038 10402 10066 10407
rect 10038 10355 10066 10374
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9982 10122 10010 10127
rect 9702 9617 9842 9618
rect 9702 9591 9703 9617
rect 9729 9591 9842 9617
rect 9702 9590 9842 9591
rect 9870 9730 9898 9735
rect 9870 9617 9898 9702
rect 9870 9591 9871 9617
rect 9897 9591 9898 9617
rect 9702 9585 9730 9590
rect 9870 9506 9898 9591
rect 9982 9561 10010 10094
rect 9982 9535 9983 9561
rect 10009 9535 10010 9561
rect 9982 9529 10010 9535
rect 9814 9478 9898 9506
rect 9814 9170 9842 9478
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 10094 9337 10122 11270
rect 10262 11465 10290 11471
rect 10262 11439 10263 11465
rect 10289 11439 10290 11465
rect 10262 11074 10290 11439
rect 10934 11354 10962 11359
rect 10710 11186 10738 11191
rect 10598 11185 10738 11186
rect 10598 11159 10711 11185
rect 10737 11159 10738 11185
rect 10598 11158 10738 11159
rect 10262 11041 10290 11046
rect 10374 11130 10402 11135
rect 10374 10905 10402 11102
rect 10374 10879 10375 10905
rect 10401 10879 10402 10905
rect 10374 10873 10402 10879
rect 10486 10849 10514 10855
rect 10486 10823 10487 10849
rect 10513 10823 10514 10849
rect 10206 10290 10234 10295
rect 10206 9617 10234 10262
rect 10486 10122 10514 10823
rect 10486 10089 10514 10094
rect 10542 10794 10570 10799
rect 10598 10794 10626 11158
rect 10710 11153 10738 11158
rect 10822 11185 10850 11191
rect 10822 11159 10823 11185
rect 10849 11159 10850 11185
rect 10654 11074 10682 11079
rect 10654 11027 10682 11046
rect 10822 11018 10850 11159
rect 10934 11186 10962 11326
rect 10990 11298 11018 12222
rect 11438 11802 11466 13175
rect 11494 13201 11522 13426
rect 11494 13175 11495 13201
rect 11521 13175 11522 13201
rect 11494 13169 11522 13175
rect 11550 12753 11578 13510
rect 11998 13454 12026 13903
rect 12334 13593 12362 14014
rect 12334 13567 12335 13593
rect 12361 13567 12362 13593
rect 12334 13561 12362 13567
rect 12558 13538 12586 13543
rect 12558 13491 12586 13510
rect 12726 13537 12754 18607
rect 12894 18354 12922 20510
rect 13118 19138 13146 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 13118 19105 13146 19110
rect 14686 19138 14714 19143
rect 14686 19091 14714 19110
rect 14294 19025 14322 19031
rect 14294 18999 14295 19025
rect 14321 18999 14322 19025
rect 13118 18746 13146 18751
rect 13118 18699 13146 18718
rect 12894 18321 12922 18326
rect 13398 18354 13426 18359
rect 13398 18307 13426 18326
rect 12726 13511 12727 13537
rect 12753 13511 12754 13537
rect 12726 13454 12754 13511
rect 11886 13426 12026 13454
rect 12670 13426 12754 13454
rect 12894 18241 12922 18247
rect 12894 18215 12895 18241
rect 12921 18215 12922 18241
rect 12894 13481 12922 18215
rect 12894 13455 12895 13481
rect 12921 13455 12922 13481
rect 12894 13449 12922 13455
rect 13174 13538 13202 13543
rect 11886 13202 11914 13426
rect 11942 13258 11970 13263
rect 11942 13257 12082 13258
rect 11942 13231 11943 13257
rect 11969 13231 12082 13257
rect 11942 13230 12082 13231
rect 11942 13225 11970 13230
rect 11886 13169 11914 13174
rect 11998 13146 12026 13151
rect 11998 13099 12026 13118
rect 11942 13033 11970 13039
rect 11942 13007 11943 13033
rect 11969 13007 11970 13033
rect 11886 12810 11914 12815
rect 11942 12810 11970 13007
rect 11886 12809 11970 12810
rect 11886 12783 11887 12809
rect 11913 12783 11970 12809
rect 11886 12782 11970 12783
rect 11886 12777 11914 12782
rect 11550 12727 11551 12753
rect 11577 12727 11578 12753
rect 11550 12721 11578 12727
rect 11438 11769 11466 11774
rect 11886 11802 11914 11807
rect 11270 11522 11298 11527
rect 11270 11475 11298 11494
rect 11102 11298 11130 11303
rect 10990 11297 11130 11298
rect 10990 11271 11103 11297
rect 11129 11271 11130 11297
rect 10990 11270 11130 11271
rect 11102 11265 11130 11270
rect 10990 11186 11018 11191
rect 10934 11185 11018 11186
rect 10934 11159 10991 11185
rect 11017 11159 11018 11185
rect 10934 11158 11018 11159
rect 10822 10905 10850 10990
rect 10822 10879 10823 10905
rect 10849 10879 10850 10905
rect 10822 10873 10850 10879
rect 10878 11130 10906 11135
rect 10542 10793 10598 10794
rect 10542 10767 10543 10793
rect 10569 10767 10598 10793
rect 10542 10766 10598 10767
rect 10206 9591 10207 9617
rect 10233 9591 10234 9617
rect 10206 9585 10234 9591
rect 10318 9506 10346 9511
rect 10318 9459 10346 9478
rect 10094 9311 10095 9337
rect 10121 9311 10122 9337
rect 9926 9226 9954 9231
rect 9926 9179 9954 9198
rect 9814 9137 9842 9142
rect 9646 8969 9674 8974
rect 9702 9113 9730 9119
rect 9702 9087 9703 9113
rect 9729 9087 9730 9113
rect 9590 8801 9618 8806
rect 9310 8745 9338 8750
rect 9646 8721 9674 8727
rect 9646 8695 9647 8721
rect 9673 8695 9674 8721
rect 9366 8666 9394 8671
rect 9198 8497 9282 8498
rect 9198 8471 9199 8497
rect 9225 8471 9282 8497
rect 9198 8470 9282 8471
rect 9198 8465 9226 8470
rect 9142 8385 9170 8391
rect 9142 8359 9143 8385
rect 9169 8359 9170 8385
rect 8806 8023 8807 8049
rect 8833 8023 8834 8049
rect 8806 8017 8834 8023
rect 8974 8049 9002 8055
rect 8974 8023 8975 8049
rect 9001 8023 9002 8049
rect 7910 7569 7938 7574
rect 8190 7938 8218 7943
rect 8190 7321 8218 7910
rect 8862 7938 8890 7943
rect 8862 7891 8890 7910
rect 8974 7938 9002 8023
rect 9030 8050 9058 8055
rect 9030 8003 9058 8022
rect 9142 8049 9170 8359
rect 9142 8023 9143 8049
rect 9169 8023 9170 8049
rect 9142 8017 9170 8023
rect 8974 7769 9002 7910
rect 8974 7743 8975 7769
rect 9001 7743 9002 7769
rect 8750 7658 8778 7663
rect 8694 7602 8722 7621
rect 8750 7611 8778 7630
rect 8694 7569 8722 7574
rect 8190 7295 8191 7321
rect 8217 7295 8218 7321
rect 8190 7289 8218 7295
rect 7854 7239 7855 7265
rect 7881 7239 7882 7265
rect 7686 6762 7714 6767
rect 7350 6706 7378 6711
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 7350 6481 7378 6678
rect 7686 6537 7714 6734
rect 7854 6706 7882 7239
rect 8918 6986 8946 6991
rect 8918 6939 8946 6958
rect 8862 6762 8890 6767
rect 8862 6715 8890 6734
rect 7854 6673 7882 6678
rect 8918 6706 8946 6711
rect 7686 6511 7687 6537
rect 7713 6511 7714 6537
rect 7686 6505 7714 6511
rect 8750 6537 8778 6543
rect 8750 6511 8751 6537
rect 8777 6511 8778 6537
rect 7350 6455 7351 6481
rect 7377 6455 7378 6481
rect 7350 6449 7378 6455
rect 8750 6090 8778 6511
rect 8918 6482 8946 6678
rect 8974 6650 9002 7743
rect 9254 7770 9282 8470
rect 9310 8386 9338 8391
rect 9310 8339 9338 8358
rect 9366 8162 9394 8638
rect 9646 8666 9674 8695
rect 9646 8633 9674 8638
rect 9478 8442 9506 8447
rect 9478 8441 9562 8442
rect 9478 8415 9479 8441
rect 9505 8415 9562 8441
rect 9478 8414 9562 8415
rect 9478 8409 9506 8414
rect 9366 8049 9394 8134
rect 9366 8023 9367 8049
rect 9393 8023 9394 8049
rect 9366 8017 9394 8023
rect 9422 7937 9450 7943
rect 9422 7911 9423 7937
rect 9449 7911 9450 7937
rect 9310 7770 9338 7775
rect 9254 7769 9338 7770
rect 9254 7743 9311 7769
rect 9337 7743 9338 7769
rect 9254 7742 9338 7743
rect 9310 7737 9338 7742
rect 9422 7770 9450 7911
rect 9478 7938 9506 7943
rect 9478 7891 9506 7910
rect 9422 7737 9450 7742
rect 9086 7658 9114 7663
rect 9086 7611 9114 7630
rect 9422 7658 9450 7663
rect 9422 7611 9450 7630
rect 9254 7321 9282 7327
rect 9254 7295 9255 7321
rect 9281 7295 9282 7321
rect 9254 7266 9282 7295
rect 9534 7266 9562 8414
rect 9646 8386 9674 8391
rect 9646 8049 9674 8358
rect 9646 8023 9647 8049
rect 9673 8023 9674 8049
rect 9646 8017 9674 8023
rect 9702 7994 9730 9087
rect 9870 8778 9898 8783
rect 9814 8750 9870 8778
rect 9814 8050 9842 8750
rect 9870 8745 9898 8750
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 10094 8106 10122 9311
rect 10486 9225 10514 9231
rect 10486 9199 10487 9225
rect 10513 9199 10514 9225
rect 10486 9114 10514 9199
rect 10486 9081 10514 9086
rect 10542 9113 10570 10766
rect 10598 10747 10626 10766
rect 10654 10793 10682 10799
rect 10654 10767 10655 10793
rect 10681 10767 10682 10793
rect 10654 10738 10682 10767
rect 10654 10514 10682 10710
rect 10878 10737 10906 11102
rect 10990 10962 11018 11158
rect 11830 11186 11858 11191
rect 11550 11129 11578 11135
rect 11550 11103 11551 11129
rect 11577 11103 11578 11129
rect 11550 10962 11578 11103
rect 11830 11129 11858 11158
rect 11830 11103 11831 11129
rect 11857 11103 11858 11129
rect 11830 11097 11858 11103
rect 10990 10929 11018 10934
rect 11326 10934 11578 10962
rect 11662 11074 11690 11079
rect 10934 10906 10962 10911
rect 10934 10859 10962 10878
rect 11214 10906 11242 10911
rect 10878 10711 10879 10737
rect 10905 10711 10906 10737
rect 10878 10705 10906 10711
rect 10598 10486 10682 10514
rect 10766 10514 10794 10519
rect 10598 9954 10626 10486
rect 10766 10467 10794 10486
rect 10654 10402 10682 10407
rect 10654 10401 10906 10402
rect 10654 10375 10655 10401
rect 10681 10375 10906 10401
rect 10654 10374 10906 10375
rect 10654 10369 10682 10374
rect 10710 9954 10738 9959
rect 10598 9926 10710 9954
rect 10542 9087 10543 9113
rect 10569 9087 10570 9113
rect 10094 8073 10122 8078
rect 9870 8050 9898 8055
rect 9842 8049 9898 8050
rect 9842 8023 9871 8049
rect 9897 8023 9898 8049
rect 9842 8022 9898 8023
rect 9814 8003 9842 8022
rect 9870 8017 9898 8022
rect 10206 8050 10234 8055
rect 10542 8050 10570 9087
rect 10598 9562 10626 9567
rect 10598 8553 10626 9534
rect 10710 9561 10738 9926
rect 10822 9618 10850 9623
rect 10710 9535 10711 9561
rect 10737 9535 10738 9561
rect 10710 9529 10738 9535
rect 10766 9617 10850 9618
rect 10766 9591 10823 9617
rect 10849 9591 10850 9617
rect 10766 9590 10850 9591
rect 10766 9281 10794 9590
rect 10822 9585 10850 9590
rect 10878 9618 10906 10374
rect 10934 10289 10962 10295
rect 10934 10263 10935 10289
rect 10961 10263 10962 10289
rect 10934 10178 10962 10263
rect 11102 10290 11130 10295
rect 11102 10243 11130 10262
rect 10934 10145 10962 10150
rect 11214 10234 11242 10878
rect 10766 9255 10767 9281
rect 10793 9255 10794 9281
rect 10654 9225 10682 9231
rect 10654 9199 10655 9225
rect 10681 9199 10682 9225
rect 10654 9058 10682 9199
rect 10766 9226 10794 9255
rect 10822 9506 10850 9511
rect 10878 9506 10906 9590
rect 11158 9561 11186 9567
rect 11158 9535 11159 9561
rect 11185 9535 11186 9561
rect 11158 9506 11186 9535
rect 10878 9478 11186 9506
rect 10822 9281 10850 9478
rect 10822 9255 10823 9281
rect 10849 9255 10850 9281
rect 10822 9249 10850 9255
rect 10766 9193 10794 9198
rect 10654 9025 10682 9030
rect 10598 8527 10599 8553
rect 10625 8527 10626 8553
rect 10598 8521 10626 8527
rect 10710 8498 10738 8503
rect 10710 8451 10738 8470
rect 10934 8441 10962 9478
rect 11046 9226 11074 9231
rect 10990 9170 11018 9175
rect 10990 9123 11018 9142
rect 10934 8415 10935 8441
rect 10961 8415 10962 8441
rect 10934 8409 10962 8415
rect 11046 9113 11074 9198
rect 11046 9087 11047 9113
rect 11073 9087 11074 9113
rect 11046 8441 11074 9087
rect 11158 8946 11186 8951
rect 11214 8946 11242 10206
rect 11186 8918 11242 8946
rect 11270 10794 11298 10799
rect 11326 10794 11354 10934
rect 11382 10850 11410 10855
rect 11382 10803 11410 10822
rect 11550 10850 11578 10855
rect 11550 10803 11578 10822
rect 11270 10793 11354 10794
rect 11270 10767 11271 10793
rect 11297 10767 11354 10793
rect 11270 10766 11354 10767
rect 11494 10793 11522 10799
rect 11494 10767 11495 10793
rect 11521 10767 11522 10793
rect 11270 10289 11298 10766
rect 11270 10263 11271 10289
rect 11297 10263 11298 10289
rect 11158 8913 11186 8918
rect 11270 8498 11298 10263
rect 11494 10010 11522 10767
rect 11662 10737 11690 11046
rect 11662 10711 11663 10737
rect 11689 10711 11690 10737
rect 11662 10705 11690 10711
rect 11830 10793 11858 10799
rect 11830 10767 11831 10793
rect 11857 10767 11858 10793
rect 11718 10402 11746 10407
rect 11774 10402 11802 10407
rect 11746 10401 11802 10402
rect 11746 10375 11775 10401
rect 11801 10375 11802 10401
rect 11746 10374 11802 10375
rect 11326 9562 11354 9567
rect 11326 9515 11354 9534
rect 11494 9282 11522 9982
rect 11662 10178 11690 10183
rect 11606 9730 11634 9735
rect 11606 9617 11634 9702
rect 11606 9591 11607 9617
rect 11633 9591 11634 9617
rect 11550 9505 11578 9511
rect 11550 9479 11551 9505
rect 11577 9479 11578 9505
rect 11550 9450 11578 9479
rect 11606 9506 11634 9591
rect 11606 9473 11634 9478
rect 11550 9417 11578 9422
rect 11494 9249 11522 9254
rect 11606 9281 11634 9287
rect 11606 9255 11607 9281
rect 11633 9255 11634 9281
rect 11438 9225 11466 9231
rect 11438 9199 11439 9225
rect 11465 9199 11466 9225
rect 11438 9114 11466 9199
rect 11438 9081 11466 9086
rect 11606 9002 11634 9255
rect 11606 8969 11634 8974
rect 11270 8451 11298 8470
rect 11046 8415 11047 8441
rect 11073 8415 11074 8441
rect 11046 8409 11074 8415
rect 11102 8441 11130 8447
rect 11102 8415 11103 8441
rect 11129 8415 11130 8441
rect 10654 8385 10682 8391
rect 10654 8359 10655 8385
rect 10681 8359 10682 8385
rect 10654 8162 10682 8359
rect 10822 8162 10850 8167
rect 10654 8161 10850 8162
rect 10654 8135 10823 8161
rect 10849 8135 10850 8161
rect 10654 8134 10850 8135
rect 10822 8129 10850 8134
rect 10934 8162 10962 8167
rect 10934 8115 10962 8134
rect 11046 8106 11074 8111
rect 11046 8059 11074 8078
rect 10206 8049 10570 8050
rect 10206 8023 10207 8049
rect 10233 8023 10570 8049
rect 10206 8022 10570 8023
rect 10206 8017 10234 8022
rect 9646 7658 9674 7663
rect 9646 7611 9674 7630
rect 9702 7574 9730 7966
rect 10094 7938 10122 7943
rect 10094 7891 10122 7910
rect 10150 7937 10178 7943
rect 10150 7911 10151 7937
rect 10177 7911 10178 7937
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9814 7713 9842 7719
rect 9814 7687 9815 7713
rect 9841 7687 9842 7713
rect 9702 7546 9786 7574
rect 9254 7238 9562 7266
rect 9478 7153 9506 7159
rect 9478 7127 9479 7153
rect 9505 7127 9506 7153
rect 9254 6818 9282 6823
rect 9478 6818 9506 7127
rect 9254 6817 9506 6818
rect 9254 6791 9255 6817
rect 9281 6791 9506 6817
rect 9254 6790 9506 6791
rect 9030 6762 9058 6767
rect 9254 6762 9282 6790
rect 9030 6761 9114 6762
rect 9030 6735 9031 6761
rect 9057 6735 9114 6761
rect 9030 6734 9114 6735
rect 9030 6729 9058 6734
rect 8974 6622 9058 6650
rect 8806 6481 8946 6482
rect 8806 6455 8919 6481
rect 8945 6455 8946 6481
rect 8806 6454 8946 6455
rect 8806 6201 8834 6454
rect 8918 6449 8946 6454
rect 8806 6175 8807 6201
rect 8833 6175 8834 6201
rect 8806 6169 8834 6175
rect 8974 6090 9002 6095
rect 8750 6089 9002 6090
rect 8750 6063 8975 6089
rect 9001 6063 9002 6089
rect 8750 6062 9002 6063
rect 9030 6090 9058 6622
rect 9086 6201 9114 6734
rect 9198 6734 9282 6762
rect 9142 6706 9170 6711
rect 9198 6706 9226 6734
rect 9170 6678 9226 6706
rect 9142 6673 9170 6678
rect 9310 6426 9338 6431
rect 9310 6379 9338 6398
rect 9086 6175 9087 6201
rect 9113 6175 9114 6201
rect 9086 6169 9114 6175
rect 9142 6090 9170 6095
rect 9030 6089 9170 6090
rect 9030 6063 9143 6089
rect 9169 6063 9170 6089
rect 9030 6062 9170 6063
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 8974 4214 9002 6062
rect 9142 6057 9170 6062
rect 8806 4186 9002 4214
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8806 1777 8834 4186
rect 9534 2169 9562 7238
rect 9758 6986 9786 7546
rect 9758 6953 9786 6958
rect 9814 6930 9842 7687
rect 10150 7574 10178 7911
rect 11102 7574 11130 8415
rect 11214 8385 11242 8391
rect 11214 8359 11215 8385
rect 11241 8359 11242 8385
rect 11214 8106 11242 8359
rect 11214 8078 11354 8106
rect 11158 7937 11186 7943
rect 11158 7911 11159 7937
rect 11185 7911 11186 7937
rect 11158 7770 11186 7911
rect 11158 7737 11186 7742
rect 11214 7937 11242 7943
rect 11214 7911 11215 7937
rect 11241 7911 11242 7937
rect 11158 7658 11186 7663
rect 11158 7611 11186 7630
rect 10038 7546 10178 7574
rect 10990 7546 11130 7574
rect 10038 7154 10066 7546
rect 10038 7126 10122 7154
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9870 6986 9898 6991
rect 9870 6939 9898 6958
rect 9982 6986 10010 6991
rect 10094 6986 10122 7126
rect 9982 6985 10122 6986
rect 9982 6959 9983 6985
rect 10009 6959 10122 6985
rect 9982 6958 10122 6959
rect 9982 6953 10010 6958
rect 9814 6897 9842 6902
rect 10206 6930 10234 6935
rect 10206 6883 10234 6902
rect 10990 6930 11018 7546
rect 10990 6897 11018 6902
rect 9758 6874 9786 6879
rect 9758 6827 9786 6846
rect 10262 6874 10290 6879
rect 10262 6827 10290 6846
rect 10374 6873 10402 6879
rect 10934 6874 10962 6879
rect 10374 6847 10375 6873
rect 10401 6847 10402 6873
rect 9814 6817 9842 6823
rect 9814 6791 9815 6817
rect 9841 6791 9842 6817
rect 9814 6426 9842 6791
rect 9814 6393 9842 6398
rect 10374 6537 10402 6847
rect 10374 6511 10375 6537
rect 10401 6511 10402 6537
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 10374 4214 10402 6511
rect 10878 6873 10962 6874
rect 10878 6847 10935 6873
rect 10961 6847 10962 6873
rect 10878 6846 10962 6847
rect 10878 6762 10906 6846
rect 10934 6841 10962 6846
rect 10822 6482 10850 6487
rect 10878 6482 10906 6734
rect 11158 6538 11186 6543
rect 11214 6538 11242 7911
rect 11270 7938 11298 7943
rect 11270 7891 11298 7910
rect 11326 7657 11354 8078
rect 11382 7938 11410 7943
rect 11382 7769 11410 7910
rect 11382 7743 11383 7769
rect 11409 7743 11410 7769
rect 11382 7737 11410 7743
rect 11438 7770 11466 7775
rect 11466 7742 11578 7770
rect 11438 7737 11466 7742
rect 11326 7631 11327 7657
rect 11353 7631 11354 7657
rect 11326 7625 11354 7631
rect 11494 7657 11522 7663
rect 11494 7631 11495 7657
rect 11521 7631 11522 7657
rect 11438 7601 11466 7607
rect 11438 7575 11439 7601
rect 11465 7575 11466 7601
rect 11270 6930 11298 6935
rect 11438 6930 11466 7575
rect 11494 7378 11522 7631
rect 11494 7345 11522 7350
rect 11550 7321 11578 7742
rect 11662 7658 11690 10150
rect 11718 10065 11746 10374
rect 11774 10369 11802 10374
rect 11718 10039 11719 10065
rect 11745 10039 11746 10065
rect 11718 10033 11746 10039
rect 11774 10122 11802 10127
rect 11774 9617 11802 10094
rect 11830 9674 11858 10767
rect 11886 10737 11914 11774
rect 11998 11185 12026 11191
rect 11998 11159 11999 11185
rect 12025 11159 12026 11185
rect 11998 10906 12026 11159
rect 12054 11130 12082 13230
rect 12670 13201 12698 13426
rect 13062 13425 13090 13431
rect 13062 13399 13063 13425
rect 13089 13399 13090 13425
rect 13062 13314 13090 13399
rect 12894 13286 13090 13314
rect 12670 13175 12671 13201
rect 12697 13175 12698 13201
rect 12558 13146 12586 13151
rect 12558 13099 12586 13118
rect 12670 12810 12698 13175
rect 12726 13202 12754 13207
rect 12726 13155 12754 13174
rect 12894 12810 12922 13286
rect 13174 13258 13202 13510
rect 13230 13482 13258 13487
rect 13230 13435 13258 13454
rect 14294 13482 14322 18999
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 14294 13449 14322 13454
rect 13062 13257 13202 13258
rect 13062 13231 13175 13257
rect 13201 13231 13202 13257
rect 13062 13230 13202 13231
rect 13006 12810 13034 12815
rect 12670 12809 13034 12810
rect 12670 12783 13007 12809
rect 13033 12783 13034 12809
rect 12670 12782 13034 12783
rect 13006 12777 13034 12782
rect 12950 12362 12978 12367
rect 13062 12362 13090 13230
rect 13174 13225 13202 13230
rect 13230 13202 13258 13207
rect 13230 12753 13258 13174
rect 14350 13146 14378 13151
rect 13230 12727 13231 12753
rect 13257 12727 13258 12753
rect 13230 12721 13258 12727
rect 13398 12754 13426 12759
rect 13398 12753 13594 12754
rect 13398 12727 13399 12753
rect 13425 12727 13594 12753
rect 13398 12726 13594 12727
rect 13398 12721 13426 12726
rect 13286 12698 13314 12703
rect 13286 12651 13314 12670
rect 13566 12697 13594 12726
rect 13566 12671 13567 12697
rect 13593 12671 13594 12697
rect 13566 12665 13594 12671
rect 13622 12697 13650 12703
rect 13622 12671 13623 12697
rect 13649 12671 13650 12697
rect 13454 12642 13482 12647
rect 13342 12641 13482 12642
rect 13342 12615 13455 12641
rect 13481 12615 13482 12641
rect 13342 12614 13482 12615
rect 13286 12418 13314 12423
rect 13342 12418 13370 12614
rect 13454 12609 13482 12614
rect 13622 12586 13650 12671
rect 13510 12558 13650 12586
rect 14350 12698 14378 13118
rect 18830 13146 18858 13151
rect 18830 13099 18858 13118
rect 20006 13033 20034 13039
rect 20006 13007 20007 13033
rect 20033 13007 20034 13033
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 20006 12810 20034 13007
rect 20006 12777 20034 12782
rect 13510 12530 13538 12558
rect 13286 12417 13370 12418
rect 13286 12391 13287 12417
rect 13313 12391 13370 12417
rect 13286 12390 13370 12391
rect 13398 12502 13538 12530
rect 13286 12385 13314 12390
rect 12950 12361 13090 12362
rect 12950 12335 12951 12361
rect 12977 12335 13090 12361
rect 12950 12334 13090 12335
rect 12390 11802 12418 11807
rect 12222 11522 12250 11527
rect 12222 11297 12250 11494
rect 12222 11271 12223 11297
rect 12249 11271 12250 11297
rect 12222 11265 12250 11271
rect 12334 11521 12362 11527
rect 12334 11495 12335 11521
rect 12361 11495 12362 11521
rect 12334 11466 12362 11495
rect 12166 11130 12194 11135
rect 12054 11129 12138 11130
rect 12054 11103 12055 11129
rect 12081 11103 12138 11129
rect 12054 11102 12138 11103
rect 12054 11097 12082 11102
rect 11998 10873 12026 10878
rect 12054 10849 12082 10855
rect 12054 10823 12055 10849
rect 12081 10823 12082 10849
rect 11942 10794 11970 10799
rect 11942 10747 11970 10766
rect 11886 10711 11887 10737
rect 11913 10711 11914 10737
rect 11886 10705 11914 10711
rect 12054 10122 12082 10823
rect 12054 10089 12082 10094
rect 11942 9674 11970 9679
rect 11830 9646 11942 9674
rect 11774 9591 11775 9617
rect 11801 9591 11802 9617
rect 11774 9585 11802 9591
rect 11942 9617 11970 9646
rect 11942 9591 11943 9617
rect 11969 9591 11970 9617
rect 11886 9561 11914 9567
rect 11886 9535 11887 9561
rect 11913 9535 11914 9561
rect 11774 9281 11802 9287
rect 11774 9255 11775 9281
rect 11801 9255 11802 9281
rect 11774 9226 11802 9255
rect 11774 9193 11802 9198
rect 11886 9114 11914 9535
rect 11942 9337 11970 9591
rect 11942 9311 11943 9337
rect 11969 9311 11970 9337
rect 11942 9305 11970 9311
rect 11886 9081 11914 9086
rect 12110 8386 12138 11102
rect 12166 11083 12194 11102
rect 12278 11074 12306 11079
rect 12278 11027 12306 11046
rect 12334 10850 12362 11438
rect 12390 11185 12418 11774
rect 12670 11578 12698 11583
rect 12950 11578 12978 12334
rect 12698 11550 12950 11578
rect 12670 11531 12698 11550
rect 12390 11159 12391 11185
rect 12417 11159 12418 11185
rect 12390 11153 12418 11159
rect 12502 11129 12530 11135
rect 12502 11103 12503 11129
rect 12529 11103 12530 11129
rect 12502 11074 12530 11103
rect 12502 11018 12530 11046
rect 12334 10817 12362 10822
rect 12390 10990 12530 11018
rect 12334 10122 12362 10127
rect 12334 9617 12362 10094
rect 12334 9591 12335 9617
rect 12361 9591 12362 9617
rect 12334 9585 12362 9591
rect 12166 9505 12194 9511
rect 12166 9479 12167 9505
rect 12193 9479 12194 9505
rect 12166 8834 12194 9479
rect 12390 9450 12418 10990
rect 12782 10906 12810 10911
rect 12614 10849 12642 10855
rect 12614 10823 12615 10849
rect 12641 10823 12642 10849
rect 12614 10738 12642 10823
rect 12614 10705 12642 10710
rect 12726 10793 12754 10799
rect 12726 10767 12727 10793
rect 12753 10767 12754 10793
rect 12670 10010 12698 10015
rect 12446 10009 12698 10010
rect 12446 9983 12671 10009
rect 12697 9983 12698 10009
rect 12446 9982 12698 9983
rect 12446 9673 12474 9982
rect 12670 9977 12698 9982
rect 12726 9786 12754 10767
rect 12782 10737 12810 10878
rect 12782 10711 12783 10737
rect 12809 10711 12810 10737
rect 12782 10705 12810 10711
rect 12838 10850 12866 10855
rect 12838 10234 12866 10822
rect 12894 10458 12922 11550
rect 12950 11531 12978 11550
rect 13286 11522 13314 11527
rect 13006 11521 13314 11522
rect 13006 11495 13287 11521
rect 13313 11495 13314 11521
rect 13006 11494 13314 11495
rect 13006 11241 13034 11494
rect 13286 11489 13314 11494
rect 13398 11354 13426 12502
rect 14350 12305 14378 12670
rect 14350 12279 14351 12305
rect 14377 12279 14378 12305
rect 14350 12273 14378 12279
rect 14574 12305 14602 12311
rect 14574 12279 14575 12305
rect 14601 12279 14602 12305
rect 13006 11215 13007 11241
rect 13033 11215 13034 11241
rect 13006 11209 13034 11215
rect 13230 11326 13426 11354
rect 13622 11634 13650 11639
rect 13062 11186 13090 11191
rect 13062 11139 13090 11158
rect 12950 11074 12978 11079
rect 12950 11027 12978 11046
rect 13230 10906 13258 11326
rect 13286 11270 13426 11298
rect 13286 11185 13314 11270
rect 13398 11242 13426 11270
rect 13454 11242 13482 11247
rect 13398 11241 13482 11242
rect 13398 11215 13455 11241
rect 13481 11215 13482 11241
rect 13398 11214 13482 11215
rect 13454 11209 13482 11214
rect 13286 11159 13287 11185
rect 13313 11159 13314 11185
rect 13286 11153 13314 11159
rect 13342 11185 13370 11191
rect 13342 11159 13343 11185
rect 13369 11159 13370 11185
rect 13342 11130 13370 11159
rect 13342 11097 13370 11102
rect 13622 11129 13650 11606
rect 14350 11634 14378 11639
rect 14350 11521 14378 11606
rect 14574 11578 14602 12279
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 18830 11969 18858 11975
rect 18830 11943 18831 11969
rect 18857 11943 18858 11969
rect 18830 11634 18858 11943
rect 20006 11802 20034 11999
rect 20006 11769 20034 11774
rect 18830 11601 18858 11606
rect 20118 11633 20146 11639
rect 20118 11607 20119 11633
rect 20145 11607 20146 11633
rect 14574 11531 14602 11550
rect 14350 11495 14351 11521
rect 14377 11495 14378 11521
rect 14350 11489 14378 11495
rect 18830 11466 18858 11471
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 18830 11185 18858 11438
rect 20118 11466 20146 11607
rect 20118 11433 20146 11438
rect 18830 11159 18831 11185
rect 18857 11159 18858 11185
rect 18830 11153 18858 11159
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 13622 11103 13623 11129
rect 13649 11103 13650 11129
rect 13622 11097 13650 11103
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 13510 11073 13538 11079
rect 13510 11047 13511 11073
rect 13537 11047 13538 11073
rect 13286 10906 13314 10911
rect 13258 10905 13314 10906
rect 13258 10879 13287 10905
rect 13313 10879 13314 10905
rect 13258 10878 13314 10879
rect 13230 10859 13258 10878
rect 13286 10873 13314 10878
rect 13510 10906 13538 11047
rect 13510 10873 13538 10878
rect 14182 10906 14210 10911
rect 14210 10878 14378 10906
rect 13678 10849 13706 10855
rect 13678 10823 13679 10849
rect 13705 10823 13706 10849
rect 13174 10793 13202 10799
rect 13174 10767 13175 10793
rect 13201 10767 13202 10793
rect 12894 10457 12978 10458
rect 12894 10431 12895 10457
rect 12921 10431 12978 10457
rect 12894 10430 12978 10431
rect 12894 10425 12922 10430
rect 12502 9758 12754 9786
rect 12782 10206 12866 10234
rect 12894 10234 12922 10239
rect 12502 9730 12530 9758
rect 12502 9683 12530 9702
rect 12446 9647 12447 9673
rect 12473 9647 12474 9673
rect 12446 9641 12474 9647
rect 12446 9450 12474 9455
rect 12390 9422 12446 9450
rect 12446 9417 12474 9422
rect 12390 9226 12418 9231
rect 12166 8801 12194 8806
rect 12334 9198 12390 9226
rect 12222 8778 12250 8783
rect 12222 8731 12250 8750
rect 12334 8778 12362 9198
rect 12390 9193 12418 9198
rect 12782 9226 12810 10206
rect 12838 10122 12866 10127
rect 12838 10075 12866 10094
rect 12894 10065 12922 10206
rect 12894 10039 12895 10065
rect 12921 10039 12922 10065
rect 12894 9898 12922 10039
rect 12950 10066 12978 10430
rect 13174 10122 13202 10767
rect 13398 10794 13426 10799
rect 13398 10747 13426 10766
rect 13510 10793 13538 10799
rect 13510 10767 13511 10793
rect 13537 10767 13538 10793
rect 13342 10737 13370 10743
rect 13342 10711 13343 10737
rect 13369 10711 13370 10737
rect 13342 10178 13370 10711
rect 13342 10150 13426 10178
rect 13174 10089 13202 10094
rect 12950 10033 12978 10038
rect 13342 10066 13370 10071
rect 13006 10010 13034 10015
rect 13034 9982 13146 10010
rect 13006 9963 13034 9982
rect 12894 9870 13090 9898
rect 13062 9561 13090 9870
rect 13062 9535 13063 9561
rect 13089 9535 13090 9561
rect 13062 9529 13090 9535
rect 13118 9561 13146 9982
rect 13342 10009 13370 10038
rect 13342 9983 13343 10009
rect 13369 9983 13370 10009
rect 13118 9535 13119 9561
rect 13145 9535 13146 9561
rect 13118 9529 13146 9535
rect 13286 9617 13314 9623
rect 13286 9591 13287 9617
rect 13313 9591 13314 9617
rect 13286 9562 13314 9591
rect 13286 9529 13314 9534
rect 12950 9506 12978 9511
rect 12782 9193 12810 9198
rect 12894 9505 12978 9506
rect 12894 9479 12951 9505
rect 12977 9479 12978 9505
rect 12894 9478 12978 9479
rect 12838 9002 12866 9007
rect 12894 9002 12922 9478
rect 12950 9473 12978 9478
rect 13006 9505 13034 9511
rect 13006 9479 13007 9505
rect 13033 9479 13034 9505
rect 13006 9002 13034 9479
rect 13174 9450 13202 9455
rect 13118 9282 13146 9287
rect 13118 9226 13146 9254
rect 12866 8974 12922 9002
rect 12950 8974 13034 9002
rect 13062 9225 13146 9226
rect 13062 9199 13119 9225
rect 13145 9199 13146 9225
rect 13062 9198 13146 9199
rect 12838 8969 12866 8974
rect 12390 8890 12418 8895
rect 12390 8843 12418 8862
rect 12782 8890 12810 8895
rect 12782 8833 12810 8862
rect 12782 8807 12783 8833
rect 12809 8807 12810 8833
rect 12782 8801 12810 8807
rect 12894 8834 12922 8839
rect 12334 8731 12362 8750
rect 12894 8777 12922 8806
rect 12894 8751 12895 8777
rect 12921 8751 12922 8777
rect 12782 8442 12810 8447
rect 12110 8353 12138 8358
rect 12726 8414 12782 8442
rect 11662 7625 11690 7630
rect 12726 7657 12754 8414
rect 12782 8409 12810 8414
rect 12894 8050 12922 8751
rect 12950 8777 12978 8974
rect 12950 8751 12951 8777
rect 12977 8751 12978 8777
rect 12950 8745 12978 8751
rect 12950 8442 12978 8447
rect 13062 8442 13090 9198
rect 13118 9193 13146 9198
rect 13174 9114 13202 9422
rect 13342 9282 13370 9983
rect 13398 10010 13426 10150
rect 13510 10122 13538 10767
rect 13678 10458 13706 10823
rect 13790 10794 13818 10799
rect 14014 10794 14042 10799
rect 13790 10793 14042 10794
rect 13790 10767 13791 10793
rect 13817 10767 14015 10793
rect 14041 10767 14042 10793
rect 13790 10766 14042 10767
rect 13790 10570 13818 10766
rect 14014 10761 14042 10766
rect 13790 10537 13818 10542
rect 13678 10425 13706 10430
rect 14182 10094 14210 10878
rect 14350 10849 14378 10878
rect 14350 10823 14351 10849
rect 14377 10823 14378 10849
rect 14350 10817 14378 10823
rect 14406 10850 14434 10855
rect 14406 10803 14434 10822
rect 14798 10850 14826 10855
rect 14518 10794 14546 10799
rect 14518 10747 14546 10766
rect 13510 10066 13650 10094
rect 13398 9977 13426 9982
rect 13342 9249 13370 9254
rect 13566 9505 13594 9511
rect 13566 9479 13567 9505
rect 13593 9479 13594 9505
rect 13566 9282 13594 9479
rect 13566 9249 13594 9254
rect 13118 9086 13202 9114
rect 13510 9169 13538 9175
rect 13510 9143 13511 9169
rect 13537 9143 13538 9169
rect 13118 8833 13146 9086
rect 13454 8946 13482 8951
rect 13174 8890 13202 8895
rect 13398 8890 13426 8895
rect 13174 8843 13202 8862
rect 13286 8889 13426 8890
rect 13286 8863 13399 8889
rect 13425 8863 13426 8889
rect 13286 8862 13426 8863
rect 13118 8807 13119 8833
rect 13145 8807 13146 8833
rect 13118 8801 13146 8807
rect 13286 8497 13314 8862
rect 13398 8857 13426 8862
rect 13454 8833 13482 8918
rect 13510 8890 13538 9143
rect 13510 8857 13538 8862
rect 13454 8807 13455 8833
rect 13481 8807 13482 8833
rect 13454 8801 13482 8807
rect 13622 8833 13650 10066
rect 14070 10066 14210 10094
rect 13734 10010 13762 10015
rect 13734 9963 13762 9982
rect 13622 8807 13623 8833
rect 13649 8807 13650 8833
rect 13342 8778 13370 8783
rect 13342 8722 13370 8750
rect 13398 8722 13426 8727
rect 13342 8721 13426 8722
rect 13342 8695 13399 8721
rect 13425 8695 13426 8721
rect 13342 8694 13426 8695
rect 13398 8689 13426 8694
rect 13566 8721 13594 8727
rect 13566 8695 13567 8721
rect 13593 8695 13594 8721
rect 13286 8471 13287 8497
rect 13313 8471 13314 8497
rect 13286 8465 13314 8471
rect 12950 8441 13062 8442
rect 12950 8415 12951 8441
rect 12977 8415 13062 8441
rect 12950 8414 13062 8415
rect 12950 8409 12978 8414
rect 13062 8395 13090 8414
rect 13174 8386 13202 8391
rect 13006 8050 13034 8055
rect 12894 8049 13034 8050
rect 12894 8023 13007 8049
rect 13033 8023 13034 8049
rect 12894 8022 13034 8023
rect 13006 8017 13034 8022
rect 13174 8049 13202 8358
rect 13174 8023 13175 8049
rect 13201 8023 13202 8049
rect 13174 8017 13202 8023
rect 13566 8050 13594 8695
rect 13622 8386 13650 8807
rect 13622 8353 13650 8358
rect 13734 8386 13762 8391
rect 13622 8050 13650 8055
rect 13566 8049 13650 8050
rect 13566 8023 13623 8049
rect 13649 8023 13650 8049
rect 13566 8022 13650 8023
rect 13622 8017 13650 8022
rect 13286 7994 13314 7999
rect 13286 7947 13314 7966
rect 13734 7993 13762 8358
rect 13790 8050 13818 8055
rect 14070 8050 14098 10066
rect 14798 9953 14826 10822
rect 18830 10794 18858 10799
rect 18830 10747 18858 10766
rect 20006 10681 20034 10687
rect 20006 10655 20007 10681
rect 20033 10655 20034 10681
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 20006 10458 20034 10655
rect 20006 10425 20034 10430
rect 14798 9927 14799 9953
rect 14825 9927 14826 9953
rect 14798 9921 14826 9927
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 14574 9562 14602 9567
rect 14574 9170 14602 9534
rect 18830 9226 18858 9231
rect 18830 9179 18858 9198
rect 14574 9123 14602 9142
rect 14798 9169 14826 9175
rect 14798 9143 14799 9169
rect 14825 9143 14826 9169
rect 14406 8442 14434 8447
rect 14350 8386 14378 8391
rect 14350 8339 14378 8358
rect 14406 8386 14434 8414
rect 14574 8386 14602 8391
rect 14798 8386 14826 9143
rect 20006 9114 20034 9119
rect 20006 9067 20034 9086
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 14406 8385 14826 8386
rect 14406 8359 14575 8385
rect 14601 8359 14826 8385
rect 14406 8358 14826 8359
rect 18830 8833 18858 8839
rect 18830 8807 18831 8833
rect 18857 8807 18858 8833
rect 18830 8386 18858 8807
rect 20006 8442 20034 8863
rect 20006 8409 20034 8414
rect 13790 8049 14098 8050
rect 13790 8023 13791 8049
rect 13817 8023 14071 8049
rect 14097 8023 14098 8049
rect 13790 8022 14098 8023
rect 13790 8017 13818 8022
rect 14070 8017 14098 8022
rect 13734 7967 13735 7993
rect 13761 7967 13762 7993
rect 13734 7961 13762 7967
rect 13174 7937 13202 7943
rect 13174 7911 13175 7937
rect 13201 7911 13202 7937
rect 13118 7714 13146 7719
rect 13174 7714 13202 7911
rect 13902 7938 13930 7943
rect 13902 7891 13930 7910
rect 14014 7937 14042 7943
rect 14014 7911 14015 7937
rect 14041 7911 14042 7937
rect 13118 7713 13202 7714
rect 13118 7687 13119 7713
rect 13145 7687 13202 7713
rect 13118 7686 13202 7687
rect 13118 7681 13146 7686
rect 12726 7631 12727 7657
rect 12753 7631 12754 7657
rect 11550 7295 11551 7321
rect 11577 7295 11578 7321
rect 11550 7289 11578 7295
rect 11886 7378 11914 7383
rect 11886 7321 11914 7350
rect 11886 7295 11887 7321
rect 11913 7295 11914 7321
rect 11886 7289 11914 7295
rect 11662 7265 11690 7271
rect 11662 7239 11663 7265
rect 11689 7239 11690 7265
rect 11270 6929 11466 6930
rect 11270 6903 11271 6929
rect 11297 6903 11466 6929
rect 11270 6902 11466 6903
rect 11494 7210 11522 7215
rect 11494 6930 11522 7182
rect 11270 6897 11298 6902
rect 11494 6897 11522 6902
rect 11158 6537 11242 6538
rect 11158 6511 11159 6537
rect 11185 6511 11242 6537
rect 11158 6510 11242 6511
rect 11662 6538 11690 7239
rect 11998 7265 12026 7271
rect 11998 7239 11999 7265
rect 12025 7239 12026 7265
rect 11830 7210 11858 7215
rect 11830 7163 11858 7182
rect 11998 7154 12026 7239
rect 11998 7121 12026 7126
rect 12334 7154 12362 7159
rect 12334 6818 12362 7126
rect 12670 6818 12698 6823
rect 12726 6818 12754 7631
rect 14014 7602 14042 7911
rect 14406 7769 14434 8358
rect 14574 8353 14602 8358
rect 18830 8353 18858 8358
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 20006 8105 20034 8111
rect 20006 8079 20007 8105
rect 20033 8079 20034 8105
rect 14406 7743 14407 7769
rect 14433 7743 14434 7769
rect 14406 7737 14434 7743
rect 18830 8049 18858 8055
rect 18830 8023 18831 8049
rect 18857 8023 18858 8049
rect 14182 7602 14210 7607
rect 14014 7574 14182 7602
rect 14182 7555 14210 7574
rect 18830 7602 18858 8023
rect 20006 7770 20034 8079
rect 20006 7737 20034 7742
rect 18830 7569 18858 7574
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 12334 6817 12474 6818
rect 12334 6791 12335 6817
rect 12361 6791 12474 6817
rect 12334 6790 12474 6791
rect 12334 6785 12362 6790
rect 11158 6505 11186 6510
rect 11662 6505 11690 6510
rect 12222 6538 12250 6543
rect 12250 6510 12306 6538
rect 12222 6491 12250 6510
rect 10822 6481 10906 6482
rect 10822 6455 10823 6481
rect 10849 6455 10906 6481
rect 10822 6454 10906 6455
rect 10822 6449 10850 6454
rect 10374 4186 10570 4214
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9534 2143 9535 2169
rect 9561 2143 9562 2169
rect 9534 2137 9562 2143
rect 9422 2058 9450 2063
rect 9310 1834 9338 1839
rect 8806 1751 8807 1777
rect 8833 1751 8834 1777
rect 8806 1745 8834 1751
rect 9086 1833 9338 1834
rect 9086 1807 9311 1833
rect 9337 1807 9338 1833
rect 9086 1806 9338 1807
rect 7518 1666 7546 1671
rect 7406 1665 7546 1666
rect 7406 1639 7519 1665
rect 7545 1639 7546 1665
rect 7406 1638 7546 1639
rect 7406 400 7434 1638
rect 7518 1633 7546 1638
rect 9086 400 9114 1806
rect 9310 1801 9338 1806
rect 9422 400 9450 2030
rect 10038 2058 10066 2063
rect 10038 2011 10066 2030
rect 10430 1834 10458 1839
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10430 400 10458 1806
rect 10542 1777 10570 4186
rect 12110 2058 12138 2063
rect 11046 1834 11074 1839
rect 11046 1787 11074 1806
rect 11774 1834 11802 1839
rect 10542 1751 10543 1777
rect 10569 1751 10570 1777
rect 10542 1745 10570 1751
rect 11774 400 11802 1806
rect 12110 400 12138 2030
rect 12278 1777 12306 6510
rect 12446 6426 12474 6790
rect 12670 6817 12754 6818
rect 12670 6791 12671 6817
rect 12697 6791 12754 6817
rect 12670 6790 12754 6791
rect 12502 6762 12530 6767
rect 12670 6762 12698 6790
rect 12530 6734 12698 6762
rect 12502 6537 12530 6734
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 12502 6511 12503 6537
rect 12529 6511 12530 6537
rect 12502 6505 12530 6511
rect 12446 6398 12642 6426
rect 12614 2169 12642 6398
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 12614 2143 12615 2169
rect 12641 2143 12642 2169
rect 12614 2137 12642 2143
rect 13118 2058 13146 2063
rect 13118 2011 13146 2030
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1745 12306 1751
rect 7392 0 7448 400
rect 9072 0 9128 400
rect 9408 0 9464 400
rect 10416 0 10472 400
rect 11760 0 11816 400
rect 12096 0 12152 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 7742 19110 7770 19138
rect 8974 19137 9002 19138
rect 8974 19111 8975 19137
rect 8975 19111 9001 19137
rect 9001 19111 9002 19137
rect 8974 19110 9002 19111
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 7854 13230 7882 13258
rect 2086 13118 2114 13146
rect 966 12446 994 12474
rect 966 12249 994 12250
rect 966 12223 967 12249
rect 967 12223 993 12249
rect 993 12223 994 12249
rect 966 12222 994 12223
rect 966 11465 994 11466
rect 966 11439 967 11465
rect 967 11439 993 11465
rect 993 11439 994 11465
rect 966 11438 994 11439
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 2142 12753 2170 12754
rect 2142 12727 2143 12753
rect 2143 12727 2169 12753
rect 2169 12727 2170 12753
rect 2142 12726 2170 12727
rect 5054 12726 5082 12754
rect 2142 12361 2170 12362
rect 2142 12335 2143 12361
rect 2143 12335 2169 12361
rect 2169 12335 2170 12361
rect 2142 12334 2170 12335
rect 6174 12726 6202 12754
rect 6230 12697 6258 12698
rect 6230 12671 6231 12697
rect 6231 12671 6257 12697
rect 6257 12671 6258 12697
rect 6230 12670 6258 12671
rect 6454 12670 6482 12698
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 8078 13257 8106 13258
rect 8078 13231 8079 13257
rect 8079 13231 8105 13257
rect 8105 13231 8106 13257
rect 8078 13230 8106 13231
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 10766 19110 10794 19138
rect 11214 19137 11242 19138
rect 11214 19111 11215 19137
rect 11215 19111 11241 19137
rect 11241 19111 11242 19137
rect 11214 19110 11242 19111
rect 12110 19110 12138 19138
rect 10430 18718 10458 18746
rect 10094 18326 10122 18354
rect 10150 18214 10178 18242
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 8470 13230 8498 13258
rect 8134 13145 8162 13146
rect 8134 13119 8135 13145
rect 8135 13119 8161 13145
rect 8161 13119 8162 13145
rect 8134 13118 8162 13119
rect 8638 13118 8666 13146
rect 7406 13006 7434 13034
rect 8078 13033 8106 13034
rect 8078 13007 8079 13033
rect 8079 13007 8105 13033
rect 8105 13007 8106 13033
rect 8078 13006 8106 13007
rect 8134 12726 8162 12754
rect 6958 12334 6986 12362
rect 6342 11857 6370 11858
rect 6342 11831 6343 11857
rect 6343 11831 6369 11857
rect 6369 11831 6370 11857
rect 6342 11830 6370 11831
rect 4830 11606 4858 11634
rect 2142 11577 2170 11578
rect 2142 11551 2143 11577
rect 2143 11551 2169 11577
rect 2169 11551 2170 11577
rect 2142 11550 2170 11551
rect 5782 11438 5810 11466
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 2086 10710 2114 10738
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 6006 11073 6034 11074
rect 6006 11047 6007 11073
rect 6007 11047 6033 11073
rect 6033 11047 6034 11073
rect 6006 11046 6034 11047
rect 6566 11633 6594 11634
rect 6566 11607 6567 11633
rect 6567 11607 6593 11633
rect 6593 11607 6594 11633
rect 6566 11606 6594 11607
rect 7070 11830 7098 11858
rect 6566 11465 6594 11466
rect 6566 11439 6567 11465
rect 6567 11439 6593 11465
rect 6593 11439 6594 11465
rect 6566 11438 6594 11439
rect 6454 11102 6482 11130
rect 6902 11129 6930 11130
rect 6902 11103 6903 11129
rect 6903 11103 6929 11129
rect 6929 11103 6930 11129
rect 6902 11102 6930 11103
rect 6342 11046 6370 11074
rect 6342 10934 6370 10962
rect 6790 11046 6818 11074
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 5894 9926 5922 9954
rect 5726 9225 5754 9226
rect 5726 9199 5727 9225
rect 5727 9199 5753 9225
rect 5753 9199 5754 9225
rect 5726 9198 5754 9199
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 2142 8833 2170 8834
rect 2142 8807 2143 8833
rect 2143 8807 2169 8833
rect 2169 8807 2170 8833
rect 2142 8806 2170 8807
rect 966 8414 994 8442
rect 6118 9169 6146 9170
rect 6118 9143 6119 9169
rect 6119 9143 6145 9169
rect 6145 9143 6146 9169
rect 6118 9142 6146 9143
rect 6342 8806 6370 8834
rect 6734 8833 6762 8834
rect 6734 8807 6735 8833
rect 6735 8807 6761 8833
rect 6761 8807 6762 8833
rect 6734 8806 6762 8807
rect 6846 10990 6874 11018
rect 8358 12614 8386 12642
rect 7910 12334 7938 12362
rect 8022 12166 8050 12194
rect 9534 13118 9562 13146
rect 8470 12641 8498 12642
rect 8470 12615 8471 12641
rect 8471 12615 8497 12641
rect 8497 12615 8498 12641
rect 8470 12614 8498 12615
rect 8750 12305 8778 12306
rect 8750 12279 8751 12305
rect 8751 12279 8777 12305
rect 8777 12279 8778 12305
rect 8750 12278 8778 12279
rect 8358 11913 8386 11914
rect 8358 11887 8359 11913
rect 8359 11887 8385 11913
rect 8385 11887 8386 11913
rect 8358 11886 8386 11887
rect 7294 11857 7322 11858
rect 7294 11831 7295 11857
rect 7295 11831 7321 11857
rect 7321 11831 7322 11857
rect 7294 11830 7322 11831
rect 7462 11857 7490 11858
rect 7462 11831 7463 11857
rect 7463 11831 7489 11857
rect 7489 11831 7490 11857
rect 7462 11830 7490 11831
rect 8078 11185 8106 11186
rect 8078 11159 8079 11185
rect 8079 11159 8105 11185
rect 8105 11159 8106 11185
rect 8078 11158 8106 11159
rect 7182 10990 7210 11018
rect 7910 11073 7938 11074
rect 7910 11047 7911 11073
rect 7911 11047 7937 11073
rect 7937 11047 7938 11073
rect 7910 11046 7938 11047
rect 8302 11830 8330 11858
rect 8302 11550 8330 11578
rect 8246 11158 8274 11186
rect 8302 11326 8330 11354
rect 6958 10934 6986 10962
rect 7742 10766 7770 10794
rect 6902 9702 6930 9730
rect 7126 9198 7154 9226
rect 7406 9617 7434 9618
rect 7406 9591 7407 9617
rect 7407 9591 7433 9617
rect 7433 9591 7434 9617
rect 7406 9590 7434 9591
rect 6902 9142 6930 9170
rect 6454 8777 6482 8778
rect 6454 8751 6455 8777
rect 6455 8751 6481 8777
rect 6481 8751 6482 8777
rect 6454 8750 6482 8751
rect 7742 9617 7770 9618
rect 7742 9591 7743 9617
rect 7743 9591 7769 9617
rect 7769 9591 7770 9617
rect 7742 9590 7770 9591
rect 7574 9561 7602 9562
rect 7574 9535 7575 9561
rect 7575 9535 7601 9561
rect 7601 9535 7602 9561
rect 7574 9534 7602 9535
rect 7462 9198 7490 9226
rect 7014 8638 7042 8666
rect 7070 8694 7098 8722
rect 5726 8441 5754 8442
rect 5726 8415 5727 8441
rect 5727 8415 5753 8441
rect 5753 8415 5754 8441
rect 5726 8414 5754 8415
rect 6174 8358 6202 8386
rect 7406 8806 7434 8834
rect 7350 8777 7378 8778
rect 7350 8751 7351 8777
rect 7351 8751 7377 8777
rect 7377 8751 7378 8777
rect 7350 8750 7378 8751
rect 7238 8638 7266 8666
rect 7406 8721 7434 8722
rect 7406 8695 7407 8721
rect 7407 8695 7433 8721
rect 7433 8695 7434 8721
rect 7406 8694 7434 8695
rect 7518 9142 7546 9170
rect 7742 9198 7770 9226
rect 7630 8918 7658 8946
rect 7294 8414 7322 8442
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 6566 7742 6594 7770
rect 7630 7601 7658 7602
rect 7630 7575 7631 7601
rect 7631 7575 7657 7601
rect 7657 7575 7658 7601
rect 7630 7574 7658 7575
rect 7966 10934 7994 10962
rect 8246 10766 8274 10794
rect 7854 9673 7882 9674
rect 7854 9647 7855 9673
rect 7855 9647 7881 9673
rect 7881 9647 7882 9673
rect 7854 9646 7882 9647
rect 8078 10542 8106 10570
rect 8694 12166 8722 12194
rect 8526 11969 8554 11970
rect 8526 11943 8527 11969
rect 8527 11943 8553 11969
rect 8553 11943 8554 11969
rect 8526 11942 8554 11943
rect 8638 11830 8666 11858
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 10654 18241 10682 18242
rect 10654 18215 10655 18241
rect 10655 18215 10681 18241
rect 10681 18215 10682 18241
rect 10654 18214 10682 18215
rect 10318 13145 10346 13146
rect 10318 13119 10319 13145
rect 10319 13119 10345 13145
rect 10345 13119 10346 13145
rect 10318 13118 10346 13119
rect 10038 13006 10066 13034
rect 9534 12753 9562 12754
rect 9534 12727 9535 12753
rect 9535 12727 9561 12753
rect 9561 12727 9562 12753
rect 9534 12726 9562 12727
rect 9478 12697 9506 12698
rect 9478 12671 9479 12697
rect 9479 12671 9505 12697
rect 9505 12671 9506 12697
rect 9478 12670 9506 12671
rect 10374 13033 10402 13034
rect 10374 13007 10375 13033
rect 10375 13007 10401 13033
rect 10401 13007 10402 13033
rect 10374 13006 10402 13007
rect 10150 12670 10178 12698
rect 9198 12305 9226 12306
rect 9198 12279 9199 12305
rect 9199 12279 9225 12305
rect 9225 12279 9226 12305
rect 9198 12278 9226 12279
rect 9086 12054 9114 12082
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9422 12278 9450 12306
rect 9422 12081 9450 12082
rect 9422 12055 9423 12081
rect 9423 12055 9449 12081
rect 9449 12055 9450 12081
rect 9422 12054 9450 12055
rect 9646 11969 9674 11970
rect 9646 11943 9647 11969
rect 9647 11943 9673 11969
rect 9673 11943 9674 11969
rect 9646 11942 9674 11943
rect 9478 11913 9506 11914
rect 9478 11887 9479 11913
rect 9479 11887 9505 11913
rect 9505 11887 9506 11913
rect 9478 11886 9506 11887
rect 8694 11185 8722 11186
rect 8694 11159 8695 11185
rect 8695 11159 8721 11185
rect 8721 11159 8722 11185
rect 8694 11158 8722 11159
rect 8358 10934 8386 10962
rect 8694 10934 8722 10962
rect 8414 10878 8442 10906
rect 7966 9198 7994 9226
rect 8302 9422 8330 9450
rect 8414 9086 8442 9114
rect 7854 8358 7882 8386
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 8694 10793 8722 10794
rect 8694 10767 8695 10793
rect 8695 10767 8721 10793
rect 8721 10767 8722 10793
rect 8694 10766 8722 10767
rect 9478 11214 9506 11242
rect 9478 10934 9506 10962
rect 9590 11830 9618 11858
rect 8806 10542 8834 10570
rect 9142 10542 9170 10570
rect 8862 10262 8890 10290
rect 8694 9534 8722 9562
rect 8750 9702 8778 9730
rect 9590 10486 9618 10514
rect 9366 10262 9394 10290
rect 9534 9617 9562 9618
rect 9534 9591 9535 9617
rect 9535 9591 9561 9617
rect 9561 9591 9562 9617
rect 9534 9590 9562 9591
rect 9198 9561 9226 9562
rect 9198 9535 9199 9561
rect 9199 9535 9225 9561
rect 9225 9535 9226 9561
rect 9198 9534 9226 9535
rect 9310 9534 9338 9562
rect 8470 9030 8498 9058
rect 8694 9142 8722 9170
rect 8526 8777 8554 8778
rect 8526 8751 8527 8777
rect 8527 8751 8553 8777
rect 8553 8751 8554 8777
rect 8526 8750 8554 8751
rect 9142 9225 9170 9226
rect 9142 9199 9143 9225
rect 9143 9199 9169 9225
rect 9169 9199 9170 9225
rect 9142 9198 9170 9199
rect 9254 9422 9282 9450
rect 9590 9561 9618 9562
rect 9590 9535 9591 9561
rect 9591 9535 9617 9561
rect 9617 9535 9618 9561
rect 9590 9534 9618 9535
rect 9478 9198 9506 9226
rect 9590 9225 9618 9226
rect 9590 9199 9591 9225
rect 9591 9199 9617 9225
rect 9617 9199 9618 9225
rect 9590 9198 9618 9199
rect 8918 8833 8946 8834
rect 8918 8807 8919 8833
rect 8919 8807 8945 8833
rect 8945 8807 8946 8833
rect 8918 8806 8946 8807
rect 8862 8750 8890 8778
rect 9254 8806 9282 8834
rect 9702 11718 9730 11746
rect 9814 11830 9842 11858
rect 10654 12278 10682 12306
rect 11046 18745 11074 18746
rect 11046 18719 11047 18745
rect 11047 18719 11073 18745
rect 11073 18719 11074 18745
rect 11046 18718 11074 18719
rect 11158 18353 11186 18354
rect 11158 18327 11159 18353
rect 11159 18327 11185 18353
rect 11185 18327 11186 18353
rect 11158 18326 11186 18327
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 12446 18718 12474 18746
rect 11494 13790 11522 13818
rect 10934 13537 10962 13538
rect 10934 13511 10935 13537
rect 10935 13511 10961 13537
rect 10961 13511 10962 13537
rect 10934 13510 10962 13511
rect 11942 13817 11970 13818
rect 11942 13791 11943 13817
rect 11943 13791 11969 13817
rect 11969 13791 11970 13817
rect 11942 13790 11970 13791
rect 11494 13510 11522 13538
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 9870 11662 9898 11690
rect 9926 11158 9954 11186
rect 10934 11577 10962 11578
rect 10934 11551 10935 11577
rect 10935 11551 10961 11577
rect 10961 11551 10962 11577
rect 10934 11550 10962 11551
rect 10094 11270 10122 11298
rect 9758 10737 9786 10738
rect 9758 10711 9759 10737
rect 9759 10711 9785 10737
rect 9785 10711 9786 10737
rect 9758 10710 9786 10711
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 10038 10401 10066 10402
rect 10038 10375 10039 10401
rect 10039 10375 10065 10401
rect 10065 10375 10066 10401
rect 10038 10374 10066 10375
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9982 10094 10010 10122
rect 9870 9702 9898 9730
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 10934 11326 10962 11354
rect 10262 11046 10290 11074
rect 10374 11102 10402 11130
rect 10206 10262 10234 10290
rect 10486 10094 10514 10122
rect 10654 11073 10682 11074
rect 10654 11047 10655 11073
rect 10655 11047 10681 11073
rect 10681 11047 10682 11073
rect 10654 11046 10682 11047
rect 12558 13537 12586 13538
rect 12558 13511 12559 13537
rect 12559 13511 12585 13537
rect 12585 13511 12586 13537
rect 12558 13510 12586 13511
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 13118 19110 13146 19138
rect 14686 19137 14714 19138
rect 14686 19111 14687 19137
rect 14687 19111 14713 19137
rect 14713 19111 14714 19137
rect 14686 19110 14714 19111
rect 13118 18745 13146 18746
rect 13118 18719 13119 18745
rect 13119 18719 13145 18745
rect 13145 18719 13146 18745
rect 13118 18718 13146 18719
rect 12894 18326 12922 18354
rect 13398 18353 13426 18354
rect 13398 18327 13399 18353
rect 13399 18327 13425 18353
rect 13425 18327 13426 18353
rect 13398 18326 13426 18327
rect 13174 13510 13202 13538
rect 11886 13174 11914 13202
rect 11998 13145 12026 13146
rect 11998 13119 11999 13145
rect 11999 13119 12025 13145
rect 12025 13119 12026 13145
rect 11998 13118 12026 13119
rect 11438 11774 11466 11802
rect 11886 11774 11914 11802
rect 11270 11521 11298 11522
rect 11270 11495 11271 11521
rect 11271 11495 11297 11521
rect 11297 11495 11298 11521
rect 11270 11494 11298 11495
rect 10822 10990 10850 11018
rect 10878 11102 10906 11130
rect 10598 10766 10626 10794
rect 10318 9505 10346 9506
rect 10318 9479 10319 9505
rect 10319 9479 10345 9505
rect 10345 9479 10346 9505
rect 10318 9478 10346 9479
rect 9926 9225 9954 9226
rect 9926 9199 9927 9225
rect 9927 9199 9953 9225
rect 9953 9199 9954 9225
rect 9926 9198 9954 9199
rect 9814 9142 9842 9170
rect 9646 8974 9674 9002
rect 9590 8806 9618 8834
rect 9310 8750 9338 8778
rect 9366 8638 9394 8666
rect 7910 7574 7938 7602
rect 8190 7910 8218 7938
rect 8862 7937 8890 7938
rect 8862 7911 8863 7937
rect 8863 7911 8889 7937
rect 8889 7911 8890 7937
rect 8862 7910 8890 7911
rect 9030 8049 9058 8050
rect 9030 8023 9031 8049
rect 9031 8023 9057 8049
rect 9057 8023 9058 8049
rect 9030 8022 9058 8023
rect 8974 7910 9002 7938
rect 8750 7657 8778 7658
rect 8750 7631 8751 7657
rect 8751 7631 8777 7657
rect 8777 7631 8778 7657
rect 8750 7630 8778 7631
rect 8694 7601 8722 7602
rect 8694 7575 8695 7601
rect 8695 7575 8721 7601
rect 8721 7575 8722 7601
rect 8694 7574 8722 7575
rect 7686 6734 7714 6762
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 7350 6678 7378 6706
rect 8918 6985 8946 6986
rect 8918 6959 8919 6985
rect 8919 6959 8945 6985
rect 8945 6959 8946 6985
rect 8918 6958 8946 6959
rect 8862 6761 8890 6762
rect 8862 6735 8863 6761
rect 8863 6735 8889 6761
rect 8889 6735 8890 6761
rect 8862 6734 8890 6735
rect 7854 6678 7882 6706
rect 8918 6678 8946 6706
rect 9310 8385 9338 8386
rect 9310 8359 9311 8385
rect 9311 8359 9337 8385
rect 9337 8359 9338 8385
rect 9310 8358 9338 8359
rect 9646 8638 9674 8666
rect 9366 8134 9394 8162
rect 9478 7937 9506 7938
rect 9478 7911 9479 7937
rect 9479 7911 9505 7937
rect 9505 7911 9506 7937
rect 9478 7910 9506 7911
rect 9422 7742 9450 7770
rect 9086 7657 9114 7658
rect 9086 7631 9087 7657
rect 9087 7631 9113 7657
rect 9113 7631 9114 7657
rect 9086 7630 9114 7631
rect 9422 7657 9450 7658
rect 9422 7631 9423 7657
rect 9423 7631 9449 7657
rect 9449 7631 9450 7657
rect 9422 7630 9450 7631
rect 9646 8358 9674 8386
rect 9870 8750 9898 8778
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 10486 9086 10514 9114
rect 10654 10710 10682 10738
rect 11830 11158 11858 11186
rect 10990 10934 11018 10962
rect 11662 11046 11690 11074
rect 10934 10905 10962 10906
rect 10934 10879 10935 10905
rect 10935 10879 10961 10905
rect 10961 10879 10962 10905
rect 10934 10878 10962 10879
rect 11214 10878 11242 10906
rect 10766 10513 10794 10514
rect 10766 10487 10767 10513
rect 10767 10487 10793 10513
rect 10793 10487 10794 10513
rect 10766 10486 10794 10487
rect 10710 9926 10738 9954
rect 10094 8078 10122 8106
rect 9814 8022 9842 8050
rect 10598 9534 10626 9562
rect 11102 10289 11130 10290
rect 11102 10263 11103 10289
rect 11103 10263 11129 10289
rect 11129 10263 11130 10289
rect 11102 10262 11130 10263
rect 10934 10150 10962 10178
rect 11214 10206 11242 10234
rect 10878 9590 10906 9618
rect 10822 9478 10850 9506
rect 10766 9198 10794 9226
rect 10654 9030 10682 9058
rect 10710 8497 10738 8498
rect 10710 8471 10711 8497
rect 10711 8471 10737 8497
rect 10737 8471 10738 8497
rect 10710 8470 10738 8471
rect 11046 9198 11074 9226
rect 10990 9169 11018 9170
rect 10990 9143 10991 9169
rect 10991 9143 11017 9169
rect 11017 9143 11018 9169
rect 10990 9142 11018 9143
rect 11158 8918 11186 8946
rect 11382 10849 11410 10850
rect 11382 10823 11383 10849
rect 11383 10823 11409 10849
rect 11409 10823 11410 10849
rect 11382 10822 11410 10823
rect 11550 10849 11578 10850
rect 11550 10823 11551 10849
rect 11551 10823 11577 10849
rect 11577 10823 11578 10849
rect 11550 10822 11578 10823
rect 11718 10374 11746 10402
rect 11494 9982 11522 10010
rect 11326 9561 11354 9562
rect 11326 9535 11327 9561
rect 11327 9535 11353 9561
rect 11353 9535 11354 9561
rect 11326 9534 11354 9535
rect 11662 10150 11690 10178
rect 11606 9702 11634 9730
rect 11606 9478 11634 9506
rect 11550 9422 11578 9450
rect 11494 9254 11522 9282
rect 11438 9086 11466 9114
rect 11606 8974 11634 9002
rect 11270 8497 11298 8498
rect 11270 8471 11271 8497
rect 11271 8471 11297 8497
rect 11297 8471 11298 8497
rect 11270 8470 11298 8471
rect 10934 8161 10962 8162
rect 10934 8135 10935 8161
rect 10935 8135 10961 8161
rect 10961 8135 10962 8161
rect 10934 8134 10962 8135
rect 11046 8105 11074 8106
rect 11046 8079 11047 8105
rect 11047 8079 11073 8105
rect 11073 8079 11074 8105
rect 11046 8078 11074 8079
rect 9702 7966 9730 7994
rect 9646 7657 9674 7658
rect 9646 7631 9647 7657
rect 9647 7631 9673 7657
rect 9673 7631 9674 7657
rect 9646 7630 9674 7631
rect 10094 7937 10122 7938
rect 10094 7911 10095 7937
rect 10095 7911 10121 7937
rect 10121 7911 10122 7937
rect 10094 7910 10122 7911
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 9142 6678 9170 6706
rect 9310 6425 9338 6426
rect 9310 6399 9311 6425
rect 9311 6399 9337 6425
rect 9337 6399 9338 6425
rect 9310 6398 9338 6399
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9758 6958 9786 6986
rect 11158 7742 11186 7770
rect 11158 7657 11186 7658
rect 11158 7631 11159 7657
rect 11159 7631 11185 7657
rect 11185 7631 11186 7657
rect 11158 7630 11186 7631
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 9870 6985 9898 6986
rect 9870 6959 9871 6985
rect 9871 6959 9897 6985
rect 9897 6959 9898 6985
rect 9870 6958 9898 6959
rect 9814 6902 9842 6930
rect 10206 6929 10234 6930
rect 10206 6903 10207 6929
rect 10207 6903 10233 6929
rect 10233 6903 10234 6929
rect 10206 6902 10234 6903
rect 10990 6902 11018 6930
rect 9758 6873 9786 6874
rect 9758 6847 9759 6873
rect 9759 6847 9785 6873
rect 9785 6847 9786 6873
rect 9758 6846 9786 6847
rect 10262 6873 10290 6874
rect 10262 6847 10263 6873
rect 10263 6847 10289 6873
rect 10289 6847 10290 6873
rect 10262 6846 10290 6847
rect 9814 6398 9842 6426
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 10878 6734 10906 6762
rect 11270 7937 11298 7938
rect 11270 7911 11271 7937
rect 11271 7911 11297 7937
rect 11297 7911 11298 7937
rect 11270 7910 11298 7911
rect 11382 7910 11410 7938
rect 11438 7742 11466 7770
rect 11494 7350 11522 7378
rect 11774 10094 11802 10122
rect 12558 13145 12586 13146
rect 12558 13119 12559 13145
rect 12559 13119 12585 13145
rect 12585 13119 12586 13145
rect 12558 13118 12586 13119
rect 12726 13201 12754 13202
rect 12726 13175 12727 13201
rect 12727 13175 12753 13201
rect 12753 13175 12754 13201
rect 12726 13174 12754 13175
rect 13230 13481 13258 13482
rect 13230 13455 13231 13481
rect 13231 13455 13257 13481
rect 13257 13455 13258 13481
rect 13230 13454 13258 13455
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 14294 13454 14322 13482
rect 13230 13174 13258 13202
rect 14350 13118 14378 13146
rect 13286 12697 13314 12698
rect 13286 12671 13287 12697
rect 13287 12671 13313 12697
rect 13313 12671 13314 12697
rect 13286 12670 13314 12671
rect 18830 13145 18858 13146
rect 18830 13119 18831 13145
rect 18831 13119 18857 13145
rect 18857 13119 18858 13145
rect 18830 13118 18858 13119
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 20006 12782 20034 12810
rect 14350 12670 14378 12698
rect 12390 11774 12418 11802
rect 12222 11494 12250 11522
rect 12334 11438 12362 11466
rect 11998 10878 12026 10906
rect 11942 10793 11970 10794
rect 11942 10767 11943 10793
rect 11943 10767 11969 10793
rect 11969 10767 11970 10793
rect 11942 10766 11970 10767
rect 12054 10094 12082 10122
rect 11942 9646 11970 9674
rect 11774 9198 11802 9226
rect 11886 9086 11914 9114
rect 12166 11129 12194 11130
rect 12166 11103 12167 11129
rect 12167 11103 12193 11129
rect 12193 11103 12194 11129
rect 12166 11102 12194 11103
rect 12278 11073 12306 11074
rect 12278 11047 12279 11073
rect 12279 11047 12305 11073
rect 12305 11047 12306 11073
rect 12278 11046 12306 11047
rect 12670 11577 12698 11578
rect 12670 11551 12671 11577
rect 12671 11551 12697 11577
rect 12697 11551 12698 11577
rect 12670 11550 12698 11551
rect 12950 11577 12978 11578
rect 12950 11551 12951 11577
rect 12951 11551 12977 11577
rect 12977 11551 12978 11577
rect 12950 11550 12978 11551
rect 12502 11046 12530 11074
rect 12334 10822 12362 10850
rect 12334 10094 12362 10122
rect 12782 10878 12810 10906
rect 12614 10710 12642 10738
rect 12838 10849 12866 10850
rect 12838 10823 12839 10849
rect 12839 10823 12865 10849
rect 12865 10823 12866 10849
rect 12838 10822 12866 10823
rect 13622 11606 13650 11634
rect 13062 11185 13090 11186
rect 13062 11159 13063 11185
rect 13063 11159 13089 11185
rect 13089 11159 13090 11185
rect 13062 11158 13090 11159
rect 12950 11073 12978 11074
rect 12950 11047 12951 11073
rect 12951 11047 12977 11073
rect 12977 11047 12978 11073
rect 12950 11046 12978 11047
rect 13342 11102 13370 11130
rect 14350 11606 14378 11634
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 20006 11774 20034 11802
rect 18830 11606 18858 11634
rect 14574 11577 14602 11578
rect 14574 11551 14575 11577
rect 14575 11551 14601 11577
rect 14601 11551 14602 11577
rect 14574 11550 14602 11551
rect 18830 11438 18858 11466
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 20118 11438 20146 11466
rect 20006 11102 20034 11130
rect 13230 10878 13258 10906
rect 13510 10878 13538 10906
rect 14182 10905 14210 10906
rect 14182 10879 14183 10905
rect 14183 10879 14209 10905
rect 14209 10879 14210 10905
rect 14182 10878 14210 10879
rect 12894 10206 12922 10234
rect 12502 9729 12530 9730
rect 12502 9703 12503 9729
rect 12503 9703 12529 9729
rect 12529 9703 12530 9729
rect 12502 9702 12530 9703
rect 12446 9422 12474 9450
rect 12166 8806 12194 8834
rect 12390 9198 12418 9226
rect 12222 8777 12250 8778
rect 12222 8751 12223 8777
rect 12223 8751 12249 8777
rect 12249 8751 12250 8777
rect 12222 8750 12250 8751
rect 12838 10121 12866 10122
rect 12838 10095 12839 10121
rect 12839 10095 12865 10121
rect 12865 10095 12866 10121
rect 12838 10094 12866 10095
rect 13398 10793 13426 10794
rect 13398 10767 13399 10793
rect 13399 10767 13425 10793
rect 13425 10767 13426 10793
rect 13398 10766 13426 10767
rect 13174 10094 13202 10122
rect 12950 10038 12978 10066
rect 13342 10038 13370 10066
rect 13006 10009 13034 10010
rect 13006 9983 13007 10009
rect 13007 9983 13033 10009
rect 13033 9983 13034 10009
rect 13006 9982 13034 9983
rect 13286 9534 13314 9562
rect 12782 9198 12810 9226
rect 13174 9422 13202 9450
rect 13118 9254 13146 9282
rect 12838 8974 12866 9002
rect 12390 8889 12418 8890
rect 12390 8863 12391 8889
rect 12391 8863 12417 8889
rect 12417 8863 12418 8889
rect 12390 8862 12418 8863
rect 12782 8862 12810 8890
rect 12894 8806 12922 8834
rect 12334 8777 12362 8778
rect 12334 8751 12335 8777
rect 12335 8751 12361 8777
rect 12361 8751 12362 8777
rect 12334 8750 12362 8751
rect 12110 8358 12138 8386
rect 12782 8414 12810 8442
rect 11662 7630 11690 7658
rect 13790 10542 13818 10570
rect 13678 10430 13706 10458
rect 13510 10094 13538 10122
rect 14406 10849 14434 10850
rect 14406 10823 14407 10849
rect 14407 10823 14433 10849
rect 14433 10823 14434 10849
rect 14406 10822 14434 10823
rect 14798 10822 14826 10850
rect 14518 10793 14546 10794
rect 14518 10767 14519 10793
rect 14519 10767 14545 10793
rect 14545 10767 14546 10793
rect 14518 10766 14546 10767
rect 13398 9982 13426 10010
rect 13342 9254 13370 9282
rect 13566 9254 13594 9282
rect 13454 8918 13482 8946
rect 13174 8889 13202 8890
rect 13174 8863 13175 8889
rect 13175 8863 13201 8889
rect 13201 8863 13202 8889
rect 13174 8862 13202 8863
rect 13510 8862 13538 8890
rect 13734 10009 13762 10010
rect 13734 9983 13735 10009
rect 13735 9983 13761 10009
rect 13761 9983 13762 10009
rect 13734 9982 13762 9983
rect 13342 8750 13370 8778
rect 13062 8414 13090 8442
rect 13174 8358 13202 8386
rect 13622 8358 13650 8386
rect 13734 8358 13762 8386
rect 13286 7993 13314 7994
rect 13286 7967 13287 7993
rect 13287 7967 13313 7993
rect 13313 7967 13314 7993
rect 13286 7966 13314 7967
rect 18830 10793 18858 10794
rect 18830 10767 18831 10793
rect 18831 10767 18857 10793
rect 18857 10767 18858 10793
rect 18830 10766 18858 10767
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 20006 10430 20034 10458
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 14574 9534 14602 9562
rect 18830 9225 18858 9226
rect 18830 9199 18831 9225
rect 18831 9199 18857 9225
rect 18857 9199 18858 9225
rect 18830 9198 18858 9199
rect 14574 9169 14602 9170
rect 14574 9143 14575 9169
rect 14575 9143 14601 9169
rect 14601 9143 14602 9169
rect 14574 9142 14602 9143
rect 14406 8414 14434 8442
rect 14350 8385 14378 8386
rect 14350 8359 14351 8385
rect 14351 8359 14377 8385
rect 14377 8359 14378 8385
rect 14350 8358 14378 8359
rect 20006 9113 20034 9114
rect 20006 9087 20007 9113
rect 20007 9087 20033 9113
rect 20033 9087 20034 9113
rect 20006 9086 20034 9087
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 20006 8414 20034 8442
rect 18830 8358 18858 8386
rect 13902 7937 13930 7938
rect 13902 7911 13903 7937
rect 13903 7911 13929 7937
rect 13929 7911 13930 7937
rect 13902 7910 13930 7911
rect 11886 7350 11914 7378
rect 11494 7209 11522 7210
rect 11494 7183 11495 7209
rect 11495 7183 11521 7209
rect 11521 7183 11522 7209
rect 11494 7182 11522 7183
rect 11494 6902 11522 6930
rect 11830 7209 11858 7210
rect 11830 7183 11831 7209
rect 11831 7183 11857 7209
rect 11857 7183 11858 7209
rect 11830 7182 11858 7183
rect 11998 7126 12026 7154
rect 12334 7126 12362 7154
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 14182 7601 14210 7602
rect 14182 7575 14183 7601
rect 14183 7575 14209 7601
rect 14209 7575 14210 7601
rect 14182 7574 14210 7575
rect 20006 7742 20034 7770
rect 18830 7574 18858 7602
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 11662 6510 11690 6538
rect 12222 6537 12250 6538
rect 12222 6511 12223 6537
rect 12223 6511 12249 6537
rect 12249 6511 12250 6537
rect 12222 6510 12250 6511
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9422 2030 9450 2058
rect 10038 2057 10066 2058
rect 10038 2031 10039 2057
rect 10039 2031 10065 2057
rect 10065 2031 10066 2057
rect 10038 2030 10066 2031
rect 10430 1806 10458 1834
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 12110 2030 12138 2058
rect 11046 1833 11074 1834
rect 11046 1807 11047 1833
rect 11047 1807 11073 1833
rect 11073 1807 11074 1833
rect 11046 1806 11074 1807
rect 11774 1806 11802 1834
rect 12502 6734 12530 6762
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 13118 2057 13146 2058
rect 13118 2031 13119 2057
rect 13119 2031 13145 2057
rect 13145 2031 13146 2057
rect 13118 2030 13146 2031
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 7737 19110 7742 19138
rect 7770 19110 8974 19138
rect 9002 19110 9007 19138
rect 10761 19110 10766 19138
rect 10794 19110 11214 19138
rect 11242 19110 11247 19138
rect 12105 19110 12110 19138
rect 12138 19110 12782 19138
rect 12810 19110 12815 19138
rect 13113 19110 13118 19138
rect 13146 19110 14686 19138
rect 14714 19110 14719 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 10425 18718 10430 18746
rect 10458 18718 11046 18746
rect 11074 18718 11079 18746
rect 12441 18718 12446 18746
rect 12474 18718 13118 18746
rect 13146 18718 13151 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 10089 18326 10094 18354
rect 10122 18326 11158 18354
rect 11186 18326 11191 18354
rect 12889 18326 12894 18354
rect 12922 18326 13398 18354
rect 13426 18326 13431 18354
rect 10145 18214 10150 18242
rect 10178 18214 10654 18242
rect 10682 18214 10687 18242
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 11489 13790 11494 13818
rect 11522 13790 11942 13818
rect 11970 13790 11975 13818
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 10929 13510 10934 13538
rect 10962 13510 11494 13538
rect 11522 13510 12558 13538
rect 12586 13510 13174 13538
rect 13202 13510 13207 13538
rect 13225 13454 13230 13482
rect 13258 13454 14294 13482
rect 14322 13454 14327 13482
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 7849 13230 7854 13258
rect 7882 13230 8078 13258
rect 8106 13230 8470 13258
rect 8498 13230 8503 13258
rect 8638 13174 11886 13202
rect 11914 13174 12726 13202
rect 12754 13174 13230 13202
rect 13258 13174 13263 13202
rect 0 13146 400 13160
rect 8638 13146 8666 13174
rect 0 13118 2086 13146
rect 2114 13118 2119 13146
rect 8129 13118 8134 13146
rect 8162 13118 8638 13146
rect 8666 13118 8671 13146
rect 9529 13118 9534 13146
rect 9562 13118 10318 13146
rect 10346 13118 10351 13146
rect 11993 13118 11998 13146
rect 12026 13118 12558 13146
rect 12586 13118 12591 13146
rect 14345 13118 14350 13146
rect 14378 13118 18830 13146
rect 18858 13118 18863 13146
rect 0 13104 400 13118
rect 7401 13006 7406 13034
rect 7434 13006 8078 13034
rect 8106 13006 8111 13034
rect 10033 13006 10038 13034
rect 10066 13006 10374 13034
rect 10402 13006 10407 13034
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 20600 12810 21000 12824
rect 20001 12782 20006 12810
rect 20034 12782 21000 12810
rect 20600 12768 21000 12782
rect 2137 12726 2142 12754
rect 2170 12726 5054 12754
rect 5082 12726 6174 12754
rect 6202 12726 6207 12754
rect 7546 12726 8134 12754
rect 8162 12726 9534 12754
rect 9562 12726 9567 12754
rect 7546 12698 7574 12726
rect 6225 12670 6230 12698
rect 6258 12670 6454 12698
rect 6482 12670 7574 12698
rect 9473 12670 9478 12698
rect 9506 12670 10150 12698
rect 10178 12670 10183 12698
rect 13281 12670 13286 12698
rect 13314 12670 14350 12698
rect 14378 12670 14383 12698
rect 8353 12614 8358 12642
rect 8386 12614 8470 12642
rect 8498 12614 8503 12642
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 0 12474 400 12488
rect 0 12446 966 12474
rect 994 12446 999 12474
rect 0 12432 400 12446
rect 2137 12334 2142 12362
rect 2170 12334 6958 12362
rect 6986 12334 7910 12362
rect 7938 12334 7943 12362
rect 8745 12278 8750 12306
rect 8778 12278 9198 12306
rect 9226 12278 9422 12306
rect 9450 12278 10654 12306
rect 10682 12278 10687 12306
rect 961 12222 966 12250
rect 994 12222 999 12250
rect 0 12138 400 12152
rect 966 12138 994 12222
rect 8017 12166 8022 12194
rect 8050 12166 8694 12194
rect 8722 12166 8727 12194
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 0 12110 994 12138
rect 0 12096 400 12110
rect 9081 12054 9086 12082
rect 9114 12054 9422 12082
rect 9450 12054 9455 12082
rect 8521 11942 8526 11970
rect 8554 11942 9646 11970
rect 9674 11942 9679 11970
rect 8353 11886 8358 11914
rect 8386 11886 9478 11914
rect 9506 11886 9511 11914
rect 6337 11830 6342 11858
rect 6370 11830 7070 11858
rect 7098 11830 7294 11858
rect 7322 11830 7327 11858
rect 7457 11830 7462 11858
rect 7490 11830 8302 11858
rect 8330 11830 8638 11858
rect 8666 11830 8671 11858
rect 9585 11830 9590 11858
rect 9618 11830 9814 11858
rect 9842 11830 9847 11858
rect 20600 11802 21000 11816
rect 11433 11774 11438 11802
rect 11466 11774 11886 11802
rect 11914 11774 12390 11802
rect 12418 11774 12423 11802
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 20600 11760 21000 11774
rect 9697 11718 9702 11746
rect 9730 11718 9735 11746
rect 9702 11690 9730 11718
rect 9702 11662 9870 11690
rect 9898 11662 9903 11690
rect 4186 11606 4830 11634
rect 4858 11606 6566 11634
rect 6594 11606 6599 11634
rect 13617 11606 13622 11634
rect 13650 11606 14350 11634
rect 14378 11606 18830 11634
rect 18858 11606 18863 11634
rect 4186 11578 4214 11606
rect 2137 11550 2142 11578
rect 2170 11550 4214 11578
rect 8297 11550 8302 11578
rect 8330 11550 8335 11578
rect 10929 11550 10934 11578
rect 10962 11550 12670 11578
rect 12698 11550 12703 11578
rect 12945 11550 12950 11578
rect 12978 11550 14574 11578
rect 14602 11550 14607 11578
rect 0 11466 400 11480
rect 0 11438 966 11466
rect 994 11438 999 11466
rect 5777 11438 5782 11466
rect 5810 11438 6566 11466
rect 6594 11438 6599 11466
rect 0 11424 400 11438
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 8302 11354 8330 11550
rect 11265 11494 11270 11522
rect 11298 11494 12222 11522
rect 12250 11494 12255 11522
rect 20600 11466 21000 11480
rect 12329 11438 12334 11466
rect 12362 11438 18830 11466
rect 18858 11438 18863 11466
rect 20113 11438 20118 11466
rect 20146 11438 21000 11466
rect 20600 11424 21000 11438
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 8297 11326 8302 11354
rect 8330 11326 10934 11354
rect 10962 11326 10967 11354
rect 10089 11270 10094 11298
rect 10122 11270 13370 11298
rect 9473 11214 9478 11242
rect 9506 11214 11858 11242
rect 11830 11186 11858 11214
rect 8073 11158 8078 11186
rect 8106 11158 8246 11186
rect 8274 11158 8694 11186
rect 8722 11158 8727 11186
rect 9921 11158 9926 11186
rect 9954 11158 9959 11186
rect 11825 11158 11830 11186
rect 11858 11158 13062 11186
rect 13090 11158 13095 11186
rect 9926 11130 9954 11158
rect 13342 11130 13370 11270
rect 20600 11130 21000 11144
rect 6449 11102 6454 11130
rect 6482 11102 6902 11130
rect 6930 11102 10374 11130
rect 10402 11102 10407 11130
rect 10873 11102 10878 11130
rect 10906 11102 12166 11130
rect 12194 11102 12199 11130
rect 13337 11102 13342 11130
rect 13370 11102 13375 11130
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 20600 11088 21000 11102
rect 6001 11046 6006 11074
rect 6034 11046 6342 11074
rect 6370 11046 6790 11074
rect 6818 11046 6823 11074
rect 7905 11046 7910 11074
rect 7938 11046 10178 11074
rect 10257 11046 10262 11074
rect 10290 11046 10654 11074
rect 10682 11046 10687 11074
rect 11657 11046 11662 11074
rect 11690 11046 12278 11074
rect 12306 11046 12311 11074
rect 12497 11046 12502 11074
rect 12530 11046 12950 11074
rect 12978 11046 12983 11074
rect 10150 11018 10178 11046
rect 6841 10990 6846 11018
rect 6874 10990 7182 11018
rect 7210 10990 8498 11018
rect 10150 10990 10822 11018
rect 10850 10990 10855 11018
rect 6337 10934 6342 10962
rect 6370 10934 6958 10962
rect 6986 10934 7966 10962
rect 7994 10934 8358 10962
rect 8386 10934 8391 10962
rect 8470 10906 8498 10990
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 8689 10934 8694 10962
rect 8722 10934 9478 10962
rect 9506 10934 9511 10962
rect 10985 10934 10990 10962
rect 11018 10934 11410 10962
rect 8409 10878 8414 10906
rect 8442 10878 8498 10906
rect 10929 10878 10934 10906
rect 10962 10878 11214 10906
rect 11242 10878 11247 10906
rect 11382 10850 11410 10934
rect 11993 10878 11998 10906
rect 12026 10878 12474 10906
rect 12777 10878 12782 10906
rect 12810 10878 13230 10906
rect 13258 10878 13263 10906
rect 13505 10878 13510 10906
rect 13538 10878 14182 10906
rect 14210 10878 14215 10906
rect 12446 10850 12474 10878
rect 11377 10822 11382 10850
rect 11410 10822 11415 10850
rect 11545 10822 11550 10850
rect 11578 10822 12334 10850
rect 12362 10822 12367 10850
rect 12446 10822 12838 10850
rect 12866 10822 12871 10850
rect 14401 10822 14406 10850
rect 14434 10822 14798 10850
rect 14826 10822 15974 10850
rect 15946 10794 15974 10822
rect 7737 10766 7742 10794
rect 7770 10766 8246 10794
rect 8274 10766 8694 10794
rect 8722 10766 8727 10794
rect 10593 10766 10598 10794
rect 10626 10766 11942 10794
rect 11970 10766 11975 10794
rect 13393 10766 13398 10794
rect 13426 10766 14518 10794
rect 14546 10766 14551 10794
rect 15946 10766 18830 10794
rect 18858 10766 18863 10794
rect 2081 10710 2086 10738
rect 2114 10710 9758 10738
rect 9786 10710 9791 10738
rect 10649 10710 10654 10738
rect 10682 10710 12614 10738
rect 12642 10710 12647 10738
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 8073 10542 8078 10570
rect 8106 10542 8806 10570
rect 8834 10542 9142 10570
rect 9170 10542 13790 10570
rect 13818 10542 13823 10570
rect 9585 10486 9590 10514
rect 9618 10486 10766 10514
rect 10794 10486 10799 10514
rect 20600 10458 21000 10472
rect 13426 10430 13678 10458
rect 13706 10430 13711 10458
rect 20001 10430 20006 10458
rect 20034 10430 21000 10458
rect 10033 10374 10038 10402
rect 10066 10374 11718 10402
rect 11746 10374 11751 10402
rect 8857 10262 8862 10290
rect 8890 10262 9366 10290
rect 9394 10262 10206 10290
rect 10234 10262 11102 10290
rect 11130 10262 11135 10290
rect 13426 10234 13454 10430
rect 20600 10416 21000 10430
rect 11209 10206 11214 10234
rect 11242 10206 12894 10234
rect 12922 10206 13454 10234
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 10929 10150 10934 10178
rect 10962 10150 11662 10178
rect 11690 10150 13454 10178
rect 13426 10122 13454 10150
rect 9977 10094 9982 10122
rect 10010 10094 10486 10122
rect 10514 10094 11774 10122
rect 11802 10094 12054 10122
rect 12082 10094 12334 10122
rect 12362 10094 12367 10122
rect 12833 10094 12838 10122
rect 12866 10094 13174 10122
rect 13202 10094 13207 10122
rect 13426 10094 13510 10122
rect 13538 10094 13543 10122
rect 12945 10038 12950 10066
rect 12978 10038 13342 10066
rect 13370 10038 13375 10066
rect 11489 9982 11494 10010
rect 11522 9982 13006 10010
rect 13034 9982 13039 10010
rect 13393 9982 13398 10010
rect 13426 9982 13734 10010
rect 13762 9982 13767 10010
rect 5889 9926 5894 9954
rect 5922 9926 10710 9954
rect 10738 9926 10743 9954
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 6897 9702 6902 9730
rect 6930 9702 8750 9730
rect 8778 9702 9870 9730
rect 9898 9702 9903 9730
rect 11601 9702 11606 9730
rect 11634 9702 12502 9730
rect 12530 9702 12535 9730
rect 7849 9646 7854 9674
rect 7882 9646 11942 9674
rect 11970 9646 11975 9674
rect 7401 9590 7406 9618
rect 7434 9590 7742 9618
rect 7770 9590 7775 9618
rect 9529 9590 9534 9618
rect 9562 9590 10878 9618
rect 10906 9590 10911 9618
rect 7569 9534 7574 9562
rect 7602 9534 8694 9562
rect 8722 9534 9198 9562
rect 9226 9534 9231 9562
rect 9305 9534 9310 9562
rect 9338 9534 9590 9562
rect 9618 9534 10598 9562
rect 10626 9534 11326 9562
rect 11354 9534 11359 9562
rect 13281 9534 13286 9562
rect 13314 9534 14574 9562
rect 14602 9534 14607 9562
rect 10313 9478 10318 9506
rect 10346 9478 10822 9506
rect 10850 9478 11606 9506
rect 11634 9478 11639 9506
rect 8297 9422 8302 9450
rect 8330 9422 9254 9450
rect 9282 9422 9287 9450
rect 11545 9422 11550 9450
rect 11578 9422 12446 9450
rect 12474 9422 13174 9450
rect 13202 9422 13207 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 8694 9254 11494 9282
rect 11522 9254 11527 9282
rect 13113 9254 13118 9282
rect 13146 9254 13342 9282
rect 13370 9254 13566 9282
rect 13594 9254 13599 9282
rect 5721 9198 5726 9226
rect 5754 9198 7126 9226
rect 7154 9198 7462 9226
rect 7490 9198 7742 9226
rect 7770 9198 7966 9226
rect 7994 9198 7999 9226
rect 8694 9170 8722 9254
rect 9137 9198 9142 9226
rect 9170 9198 9478 9226
rect 9506 9198 9511 9226
rect 9585 9198 9590 9226
rect 9618 9198 9926 9226
rect 9954 9198 9959 9226
rect 10761 9198 10766 9226
rect 10794 9198 11046 9226
rect 11074 9198 11079 9226
rect 11769 9198 11774 9226
rect 11802 9198 12390 9226
rect 12418 9198 12782 9226
rect 12810 9198 12815 9226
rect 15946 9198 18830 9226
rect 18858 9198 18863 9226
rect 15946 9170 15974 9198
rect 6113 9142 6118 9170
rect 6146 9142 6902 9170
rect 6930 9142 6935 9170
rect 7513 9142 7518 9170
rect 7546 9142 8694 9170
rect 8722 9142 8727 9170
rect 9809 9142 9814 9170
rect 9842 9142 10990 9170
rect 11018 9142 11023 9170
rect 14569 9142 14574 9170
rect 14602 9142 15974 9170
rect 20600 9114 21000 9128
rect 8409 9086 8414 9114
rect 8442 9086 10486 9114
rect 10514 9086 11438 9114
rect 11466 9086 11886 9114
rect 11914 9086 11919 9114
rect 20001 9086 20006 9114
rect 20034 9086 21000 9114
rect 20600 9072 21000 9086
rect 8465 9030 8470 9058
rect 8498 9030 10654 9058
rect 10682 9030 10687 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 9641 8974 9646 9002
rect 9674 8974 11606 9002
rect 11634 8974 12838 9002
rect 12866 8974 13454 9002
rect 7625 8918 7630 8946
rect 7658 8918 11158 8946
rect 11186 8918 11191 8946
rect 13426 8918 13454 8974
rect 13482 8918 13487 8946
rect 12385 8862 12390 8890
rect 12418 8862 12782 8890
rect 12810 8862 12815 8890
rect 13169 8862 13174 8890
rect 13202 8862 13510 8890
rect 13538 8862 13543 8890
rect 2137 8806 2142 8834
rect 2170 8806 4214 8834
rect 6337 8806 6342 8834
rect 6370 8806 6734 8834
rect 6762 8806 7406 8834
rect 7434 8806 7439 8834
rect 8913 8806 8918 8834
rect 8946 8806 9254 8834
rect 9282 8806 9590 8834
rect 9618 8806 9623 8834
rect 12161 8806 12166 8834
rect 12194 8806 12894 8834
rect 12922 8806 12927 8834
rect 4186 8722 4214 8806
rect 6449 8750 6454 8778
rect 6482 8750 7350 8778
rect 7378 8750 7383 8778
rect 8521 8750 8526 8778
rect 8554 8750 8862 8778
rect 8890 8750 8895 8778
rect 9305 8750 9310 8778
rect 9338 8750 9870 8778
rect 9898 8750 12222 8778
rect 12250 8750 12255 8778
rect 12329 8750 12334 8778
rect 12362 8750 13342 8778
rect 13370 8750 13375 8778
rect 4186 8694 7070 8722
rect 7098 8694 7406 8722
rect 7434 8694 7439 8722
rect 7009 8638 7014 8666
rect 7042 8638 7238 8666
rect 7266 8638 9366 8666
rect 9394 8638 9646 8666
rect 9674 8638 9679 8666
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 10705 8470 10710 8498
rect 10738 8470 11270 8498
rect 11298 8470 11303 8498
rect 0 8442 400 8456
rect 20600 8442 21000 8456
rect 0 8414 966 8442
rect 994 8414 999 8442
rect 5721 8414 5726 8442
rect 5754 8414 6202 8442
rect 7289 8414 7294 8442
rect 7322 8414 7574 8442
rect 12777 8414 12782 8442
rect 12810 8414 13062 8442
rect 13090 8414 14406 8442
rect 14434 8414 14439 8442
rect 20001 8414 20006 8442
rect 20034 8414 21000 8442
rect 0 8400 400 8414
rect 6174 8386 6202 8414
rect 7546 8386 7574 8414
rect 20600 8400 21000 8414
rect 6169 8358 6174 8386
rect 6202 8358 6207 8386
rect 7546 8358 7854 8386
rect 7882 8358 9310 8386
rect 9338 8358 9343 8386
rect 9641 8358 9646 8386
rect 9674 8358 12110 8386
rect 12138 8358 12143 8386
rect 13169 8358 13174 8386
rect 13202 8358 13622 8386
rect 13650 8358 13655 8386
rect 13729 8358 13734 8386
rect 13762 8358 14350 8386
rect 14378 8358 18830 8386
rect 18858 8358 18863 8386
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 9361 8134 9366 8162
rect 9394 8134 10934 8162
rect 10962 8134 10967 8162
rect 10089 8078 10094 8106
rect 10122 8078 11046 8106
rect 11074 8078 11079 8106
rect 9025 8022 9030 8050
rect 9058 8022 9814 8050
rect 9842 8022 9847 8050
rect 9697 7966 9702 7994
rect 9730 7966 11298 7994
rect 13281 7966 13286 7994
rect 13314 7966 13454 7994
rect 11270 7938 11298 7966
rect 13426 7938 13454 7966
rect 8185 7910 8190 7938
rect 8218 7910 8862 7938
rect 8890 7910 8895 7938
rect 8969 7910 8974 7938
rect 9002 7910 9478 7938
rect 9506 7910 10094 7938
rect 10122 7910 10127 7938
rect 11265 7910 11270 7938
rect 11298 7910 11382 7938
rect 11410 7910 11415 7938
rect 13426 7910 13902 7938
rect 13930 7910 13935 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 20600 7770 21000 7784
rect 6561 7742 6566 7770
rect 6594 7742 9422 7770
rect 9450 7742 9455 7770
rect 11153 7742 11158 7770
rect 11186 7742 11438 7770
rect 11466 7742 11471 7770
rect 20001 7742 20006 7770
rect 20034 7742 21000 7770
rect 20600 7728 21000 7742
rect 8745 7630 8750 7658
rect 8778 7630 9086 7658
rect 9114 7630 9422 7658
rect 9450 7630 9646 7658
rect 9674 7630 9679 7658
rect 11153 7630 11158 7658
rect 11186 7630 11662 7658
rect 11690 7630 11695 7658
rect 7625 7574 7630 7602
rect 7658 7574 7910 7602
rect 7938 7574 8694 7602
rect 8722 7574 8727 7602
rect 14177 7574 14182 7602
rect 14210 7574 18830 7602
rect 18858 7574 18863 7602
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 11489 7350 11494 7378
rect 11522 7350 11886 7378
rect 11914 7350 11919 7378
rect 11489 7182 11494 7210
rect 11522 7182 11830 7210
rect 11858 7182 11863 7210
rect 11993 7126 11998 7154
rect 12026 7126 12334 7154
rect 12362 7126 12367 7154
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 8913 6958 8918 6986
rect 8946 6958 9758 6986
rect 9786 6958 9870 6986
rect 9898 6958 9903 6986
rect 9809 6902 9814 6930
rect 9842 6902 10206 6930
rect 10234 6902 10990 6930
rect 11018 6902 11494 6930
rect 11522 6902 11527 6930
rect 9753 6846 9758 6874
rect 9786 6846 10262 6874
rect 10290 6846 10295 6874
rect 7681 6734 7686 6762
rect 7714 6734 8862 6762
rect 8890 6734 8895 6762
rect 10873 6734 10878 6762
rect 10906 6734 12502 6762
rect 12530 6734 12535 6762
rect 7345 6678 7350 6706
rect 7378 6678 7854 6706
rect 7882 6678 8918 6706
rect 8946 6678 9142 6706
rect 9170 6678 9175 6706
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 11657 6510 11662 6538
rect 11690 6510 12222 6538
rect 12250 6510 12255 6538
rect 9305 6398 9310 6426
rect 9338 6398 9814 6426
rect 9842 6398 9847 6426
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 9417 2030 9422 2058
rect 9450 2030 10038 2058
rect 10066 2030 10071 2058
rect 12105 2030 12110 2058
rect 12138 2030 13118 2058
rect 13146 2030 13151 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 10425 1806 10430 1834
rect 10458 1806 11046 1834
rect 11074 1806 11079 1834
rect 11769 1806 11774 1834
rect 11802 1806 12782 1834
rect 12810 1806 12815 1834
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9072 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _106_
timestamp 1698175906
transform 1 0 8176 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11368 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_
timestamp 1698175906
transform -1 0 9576 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _110_
timestamp 1698175906
transform 1 0 7336 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _111_
timestamp 1698175906
transform 1 0 9128 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9464 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _113_
timestamp 1698175906
transform 1 0 7840 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8624 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform -1 0 8400 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _116_
timestamp 1698175906
transform -1 0 9632 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9296 0 1 11760
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _118_
timestamp 1698175906
transform 1 0 10920 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _119_
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698175906
transform 1 0 10080 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _121_
timestamp 1698175906
transform -1 0 10920 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _122_
timestamp 1698175906
transform 1 0 8008 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _123_
timestamp 1698175906
transform -1 0 8848 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _124_
timestamp 1698175906
transform 1 0 8176 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform -1 0 7560 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform 1 0 8400 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _127_
timestamp 1698175906
transform -1 0 8232 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _128_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7000 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_
timestamp 1698175906
transform 1 0 9744 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10416 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _131_
timestamp 1698175906
transform -1 0 10640 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _132_
timestamp 1698175906
transform -1 0 6328 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _133_
timestamp 1698175906
transform -1 0 6552 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _134_
timestamp 1698175906
transform 1 0 9128 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _135_
timestamp 1698175906
transform 1 0 9856 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _136_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9072 0 -1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _137_
timestamp 1698175906
transform 1 0 9912 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _138_
timestamp 1698175906
transform -1 0 8176 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _139_
timestamp 1698175906
transform -1 0 11200 0 1 10976
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _140_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10360 0 -1 11760
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _141_
timestamp 1698175906
transform -1 0 10976 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform -1 0 7000 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _143_
timestamp 1698175906
transform -1 0 9240 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _144_
timestamp 1698175906
transform 1 0 8680 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _145_
timestamp 1698175906
transform 1 0 9408 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _146_
timestamp 1698175906
transform 1 0 11032 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _147_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7672 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _148_
timestamp 1698175906
transform -1 0 12040 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _149_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12096 0 1 10976
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _150_
timestamp 1698175906
transform 1 0 9296 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _151_
timestamp 1698175906
transform -1 0 9016 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _152_
timestamp 1698175906
transform 1 0 7280 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _153_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7112 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _154_
timestamp 1698175906
transform -1 0 8176 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _155_
timestamp 1698175906
transform 1 0 8176 0 1 11760
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _156_
timestamp 1698175906
transform -1 0 12824 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _157_
timestamp 1698175906
transform -1 0 12096 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698175906
transform 1 0 13160 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _159_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12936 0 -1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform -1 0 13720 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _161_
timestamp 1698175906
transform 1 0 11760 0 -1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _162_
timestamp 1698175906
transform -1 0 12096 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _163_
timestamp 1698175906
transform -1 0 11592 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _164_
timestamp 1698175906
transform 1 0 10248 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _165_
timestamp 1698175906
transform 1 0 9632 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _166_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11704 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _167_
timestamp 1698175906
transform 1 0 9072 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _168_
timestamp 1698175906
transform 1 0 12152 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _169_
timestamp 1698175906
transform -1 0 13944 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _170_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12880 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _171_
timestamp 1698175906
transform -1 0 11704 0 1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _172_
timestamp 1698175906
transform 1 0 12712 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _173_
timestamp 1698175906
transform 1 0 11200 0 -1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _174_
timestamp 1698175906
transform 1 0 10640 0 -1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _175_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12096 0 1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _176_
timestamp 1698175906
transform -1 0 12600 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _177_
timestamp 1698175906
transform 1 0 12656 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _178_
timestamp 1698175906
transform 1 0 13944 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _179_
timestamp 1698175906
transform 1 0 14280 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _180_
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _181_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13608 0 -1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _182_
timestamp 1698175906
transform -1 0 14168 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _183_
timestamp 1698175906
transform -1 0 13384 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _184_
timestamp 1698175906
transform -1 0 13888 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _185_
timestamp 1698175906
transform -1 0 13776 0 1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _186_
timestamp 1698175906
transform -1 0 6720 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _187_
timestamp 1698175906
transform -1 0 6104 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _188_
timestamp 1698175906
transform 1 0 7224 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _189_
timestamp 1698175906
transform -1 0 6552 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _190_
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _191_
timestamp 1698175906
transform 1 0 12880 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _192_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9856 0 -1 9408
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _193_
timestamp 1698175906
transform -1 0 9240 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _194_
timestamp 1698175906
transform -1 0 9128 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _195_
timestamp 1698175906
transform 1 0 8400 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _196_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9016 0 -1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _197_
timestamp 1698175906
transform 1 0 8736 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _198_
timestamp 1698175906
transform 1 0 9576 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _199_
timestamp 1698175906
transform 1 0 10136 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _200_
timestamp 1698175906
transform -1 0 10304 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _201_
timestamp 1698175906
transform 1 0 9688 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _202_
timestamp 1698175906
transform -1 0 10808 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _203_
timestamp 1698175906
transform 1 0 11424 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _204_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10752 0 1 7840
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _205_
timestamp 1698175906
transform 1 0 11760 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _206_
timestamp 1698175906
transform -1 0 11368 0 -1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _207_
timestamp 1698175906
transform 1 0 11088 0 -1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform 1 0 6328 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform -1 0 6608 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 9296 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 5376 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 6216 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 6104 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 5656 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform -1 0 8512 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _217_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11424 0 1 12544
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 12824 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 10808 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 8848 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 13048 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 10808 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 13272 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 12656 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 12824 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform -1 0 6384 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform 1 0 5656 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 12824 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 7224 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 7728 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 8848 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 10696 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform 1 0 10808 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _236_
timestamp 1698175906
transform 1 0 12992 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _237_
timestamp 1698175906
transform 1 0 12656 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10640 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 8344 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 6720 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 7112 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 7952 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 7840 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 7728 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 13160 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 14560 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 12544 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 8736 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 14784 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 13552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 14392 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 14560 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 6832 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 7392 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 14560 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 9240 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 9464 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform -1 0 8848 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform -1 0 12544 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 9744 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9464 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 11368 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_104 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_120 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7392 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_125 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7672 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_133 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8120 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_135
timestamp 1698175906
transform 1 0 8232 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174
timestamp 1698175906
transform 1 0 10416 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698175906
transform 1 0 11928 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698175906
transform 1 0 12040 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698175906
transform 1 0 9072 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_154
timestamp 1698175906
transform 1 0 9296 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_156
timestamp 1698175906
transform 1 0 9408 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_183
timestamp 1698175906
transform 1 0 10920 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_199
timestamp 1698175906
transform 1 0 11816 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 12264 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 14000 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 15792 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 16240 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_146
timestamp 1698175906
transform 1 0 8848 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_153
timestamp 1698175906
transform 1 0 9240 0 -1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_185
timestamp 1698175906
transform 1 0 11032 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_201
timestamp 1698175906
transform 1 0 11928 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698175906
transform 1 0 12376 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_115
timestamp 1698175906
transform 1 0 7112 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_208
timestamp 1698175906
transform 1 0 12320 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_212
timestamp 1698175906
transform 1 0 12544 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698175906
transform 1 0 14336 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_144
timestamp 1698175906
transform 1 0 8736 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_151
timestamp 1698175906
transform 1 0 9128 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_155
timestamp 1698175906
transform 1 0 9352 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_159
timestamp 1698175906
transform 1 0 9576 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_175
timestamp 1698175906
transform 1 0 10472 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_179
timestamp 1698175906
transform 1 0 10696 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_216
timestamp 1698175906
transform 1 0 12768 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_123
timestamp 1698175906
transform 1 0 7560 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_125
timestamp 1698175906
transform 1 0 7672 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_155
timestamp 1698175906
transform 1 0 9352 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_159
timestamp 1698175906
transform 1 0 9576 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_185
timestamp 1698175906
transform 1 0 11032 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_189
timestamp 1698175906
transform 1 0 11256 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_191
timestamp 1698175906
transform 1 0 11368 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_204
timestamp 1698175906
transform 1 0 12096 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_236
timestamp 1698175906
transform 1 0 13888 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 14336 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_88
timestamp 1698175906
transform 1 0 5600 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_96
timestamp 1698175906
transform 1 0 6048 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_126
timestamp 1698175906
transform 1 0 7728 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_130
timestamp 1698175906
transform 1 0 7952 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698175906
transform 1 0 8400 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_146
timestamp 1698175906
transform 1 0 8848 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_165
timestamp 1698175906
transform 1 0 9912 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_181
timestamp 1698175906
transform 1 0 10808 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_185
timestamp 1698175906
transform 1 0 11032 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_196
timestamp 1698175906
transform 1 0 11648 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_204
timestamp 1698175906
transform 1 0 12096 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698175906
transform 1 0 12320 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_243
timestamp 1698175906
transform 1 0 14280 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_247
timestamp 1698175906
transform 1 0 14504 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 16296 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_139
timestamp 1698175906
transform 1 0 8456 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_143
timestamp 1698175906
transform 1 0 8680 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_162
timestamp 1698175906
transform 1 0 9744 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698175906
transform 1 0 10304 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 10416 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_177
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_179
timestamp 1698175906
transform 1 0 10696 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_192
timestamp 1698175906
transform 1 0 11424 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_208
timestamp 1698175906
transform 1 0 12320 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_216
timestamp 1698175906
transform 1 0 12768 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_218
timestamp 1698175906
transform 1 0 12880 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_227
timestamp 1698175906
transform 1 0 13384 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698175906
transform 1 0 14168 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 18648 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_88
timestamp 1698175906
transform 1 0 5600 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_118
timestamp 1698175906
transform 1 0 7280 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_122
timestamp 1698175906
transform 1 0 7504 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698175906
transform 1 0 8400 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_146
timestamp 1698175906
transform 1 0 8848 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_148
timestamp 1698175906
transform 1 0 8960 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_159
timestamp 1698175906
transform 1 0 9576 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_191
timestamp 1698175906
transform 1 0 11368 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698175906
transform 1 0 12264 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 12376 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_216
timestamp 1698175906
transform 1 0 12768 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_246
timestamp 1698175906
transform 1 0 14448 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_250
timestamp 1698175906
transform 1 0 14672 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_266
timestamp 1698175906
transform 1 0 15568 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_274
timestamp 1698175906
transform 1 0 16016 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698175906
transform 1 0 16240 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 20048 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 20160 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_69
timestamp 1698175906
transform 1 0 4536 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_85
timestamp 1698175906
transform 1 0 5432 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_93
timestamp 1698175906
transform 1 0 5880 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_97
timestamp 1698175906
transform 1 0 6104 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_115
timestamp 1698175906
transform 1 0 7112 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_125
timestamp 1698175906
transform 1 0 7672 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_133
timestamp 1698175906
transform 1 0 8120 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_137
timestamp 1698175906
transform 1 0 8344 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_149
timestamp 1698175906
transform 1 0 9016 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_162
timestamp 1698175906
transform 1 0 9744 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_170
timestamp 1698175906
transform 1 0 10192 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 10416 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_177
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_193
timestamp 1698175906
transform 1 0 11480 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_201
timestamp 1698175906
transform 1 0 11928 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_211
timestamp 1698175906
transform 1 0 12488 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_234
timestamp 1698175906
transform 1 0 13776 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_242
timestamp 1698175906
transform 1 0 14224 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 14336 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_88
timestamp 1698175906
transform 1 0 5600 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_124
timestamp 1698175906
transform 1 0 7616 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_128
timestamp 1698175906
transform 1 0 7840 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698175906
transform 1 0 8288 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_148
timestamp 1698175906
transform 1 0 8960 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_170
timestamp 1698175906
transform 1 0 10192 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_187
timestamp 1698175906
transform 1 0 11144 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_203
timestamp 1698175906
transform 1 0 12040 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698175906
transform 1 0 12264 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 12376 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_220
timestamp 1698175906
transform 1 0 12992 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_250
timestamp 1698175906
transform 1 0 14672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_254
timestamp 1698175906
transform 1 0 14896 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_270
timestamp 1698175906
transform 1 0 15792 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 16240 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 18256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 18704 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_115
timestamp 1698175906
transform 1 0 7112 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_139
timestamp 1698175906
transform 1 0 8456 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698175906
transform 1 0 10416 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_177
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_213
timestamp 1698175906
transform 1 0 12600 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_217
timestamp 1698175906
transform 1 0 12824 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_228
timestamp 1698175906
transform 1 0 13440 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_232
timestamp 1698175906
transform 1 0 13664 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_240
timestamp 1698175906
transform 1 0 14112 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 14336 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_80
timestamp 1698175906
transform 1 0 5152 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_113
timestamp 1698175906
transform 1 0 7000 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_117
timestamp 1698175906
transform 1 0 7224 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_125
timestamp 1698175906
transform 1 0 7672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_127
timestamp 1698175906
transform 1 0 7784 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_150
timestamp 1698175906
transform 1 0 9072 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_207
timestamp 1698175906
transform 1 0 12264 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 12376 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_222
timestamp 1698175906
transform 1 0 13104 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_224
timestamp 1698175906
transform 1 0 13216 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_254
timestamp 1698175906
transform 1 0 14896 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_270
timestamp 1698175906
transform 1 0 15792 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 16240 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 20048 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 20160 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_123
timestamp 1698175906
transform 1 0 7560 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698175906
transform 1 0 14168 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_88
timestamp 1698175906
transform 1 0 5600 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_96
timestamp 1698175906
transform 1 0 6048 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_98
timestamp 1698175906
transform 1 0 6160 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_128
timestamp 1698175906
transform 1 0 7840 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_132
timestamp 1698175906
transform 1 0 8064 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_148
timestamp 1698175906
transform 1 0 8960 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_160
timestamp 1698175906
transform 1 0 9632 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_164
timestamp 1698175906
transform 1 0 9856 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_172
timestamp 1698175906
transform 1 0 10304 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_185
timestamp 1698175906
transform 1 0 11032 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_187
timestamp 1698175906
transform 1 0 11144 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_205
timestamp 1698175906
transform 1 0 12152 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 12376 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_219
timestamp 1698175906
transform 1 0 12936 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_221
timestamp 1698175906
transform 1 0 13048 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_248
timestamp 1698175906
transform 1 0 14560 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_69
timestamp 1698175906
transform 1 0 4536 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_85
timestamp 1698175906
transform 1 0 5432 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_97
timestamp 1698175906
transform 1 0 6104 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_113
timestamp 1698175906
transform 1 0 7000 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_121
timestamp 1698175906
transform 1 0 7448 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_125
timestamp 1698175906
transform 1 0 7672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_127
timestamp 1698175906
transform 1 0 7784 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_146
timestamp 1698175906
transform 1 0 8848 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_162
timestamp 1698175906
transform 1 0 9744 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_170
timestamp 1698175906
transform 1 0 10192 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 10416 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_188
timestamp 1698175906
transform 1 0 11200 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_190
timestamp 1698175906
transform 1 0 11312 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_213
timestamp 1698175906
transform 1 0 12600 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_217
timestamp 1698175906
transform 1 0 12824 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_233
timestamp 1698175906
transform 1 0 13720 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_241
timestamp 1698175906
transform 1 0 14168 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 2240 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 4032 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 4480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_102
timestamp 1698175906
transform 1 0 6384 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_108
timestamp 1698175906
transform 1 0 6720 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_112
timestamp 1698175906
transform 1 0 6944 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_128
timestamp 1698175906
transform 1 0 7840 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_132
timestamp 1698175906
transform 1 0 8064 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 8456 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_158
timestamp 1698175906
transform 1 0 9520 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_162
timestamp 1698175906
transform 1 0 9744 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_173
timestamp 1698175906
transform 1 0 10360 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_216
timestamp 1698175906
transform 1 0 12768 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_246
timestamp 1698175906
transform 1 0 14448 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_250
timestamp 1698175906
transform 1 0 14672 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_266
timestamp 1698175906
transform 1 0 15568 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_274
timestamp 1698175906
transform 1 0 16016 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698175906
transform 1 0 16240 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_330
timestamp 1698175906
transform 1 0 19152 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_338
timestamp 1698175906
transform 1 0 19600 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_342
timestamp 1698175906
transform 1 0 19824 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_344
timestamp 1698175906
transform 1 0 19936 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_69
timestamp 1698175906
transform 1 0 4536 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_85
timestamp 1698175906
transform 1 0 5432 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_93
timestamp 1698175906
transform 1 0 5880 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_115
timestamp 1698175906
transform 1 0 7112 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_123
timestamp 1698175906
transform 1 0 7560 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_127
timestamp 1698175906
transform 1 0 7784 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_145
timestamp 1698175906
transform 1 0 8792 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_153
timestamp 1698175906
transform 1 0 9240 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_170
timestamp 1698175906
transform 1 0 10192 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 10416 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698175906
transform 1 0 14168 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 2240 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 4032 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 4480 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_76
timestamp 1698175906
transform 1 0 4928 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_106
timestamp 1698175906
transform 1 0 6608 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_110
timestamp 1698175906
transform 1 0 6832 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_146
timestamp 1698175906
transform 1 0 8848 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_150
timestamp 1698175906
transform 1 0 9072 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_183
timestamp 1698175906
transform 1 0 10920 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_199
timestamp 1698175906
transform 1 0 11816 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_207
timestamp 1698175906
transform 1 0 12264 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698175906
transform 1 0 12376 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_216
timestamp 1698175906
transform 1 0 12768 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_246
timestamp 1698175906
transform 1 0 14448 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_250
timestamp 1698175906
transform 1 0 14672 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_266
timestamp 1698175906
transform 1 0 15568 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_274
timestamp 1698175906
transform 1 0 16016 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698175906
transform 1 0 16240 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 2240 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 2464 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_69
timestamp 1698175906
transform 1 0 4536 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_85
timestamp 1698175906
transform 1 0 5432 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_93
timestamp 1698175906
transform 1 0 5880 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_95
timestamp 1698175906
transform 1 0 5992 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_111
timestamp 1698175906
transform 1 0 6888 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_121
timestamp 1698175906
transform 1 0 7448 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_129
timestamp 1698175906
transform 1 0 7896 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_131
timestamp 1698175906
transform 1 0 8008 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_144
timestamp 1698175906
transform 1 0 8736 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_152
timestamp 1698175906
transform 1 0 9184 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_154
timestamp 1698175906
transform 1 0 9296 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_168
timestamp 1698175906
transform 1 0 10080 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698175906
transform 1 0 10304 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 10416 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_185
timestamp 1698175906
transform 1 0 11032 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_189
timestamp 1698175906
transform 1 0 11256 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_191
timestamp 1698175906
transform 1 0 11368 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_233
timestamp 1698175906
transform 1 0 13720 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698175906
transform 1 0 14168 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_88
timestamp 1698175906
transform 1 0 5600 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_96
timestamp 1698175906
transform 1 0 6048 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_100
timestamp 1698175906
transform 1 0 6272 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_135
timestamp 1698175906
transform 1 0 8232 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 8456 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_176
timestamp 1698175906
transform 1 0 10528 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_180
timestamp 1698175906
transform 1 0 10752 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_188
timestamp 1698175906
transform 1 0 11200 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_195
timestamp 1698175906
transform 1 0 11592 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_204
timestamp 1698175906
transform 1 0 12096 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698175906
transform 1 0 12320 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_217
timestamp 1698175906
transform 1 0 12824 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_221
timestamp 1698175906
transform 1 0 13048 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_225
timestamp 1698175906
transform 1 0 13272 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_257
timestamp 1698175906
transform 1 0 15064 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_273
timestamp 1698175906
transform 1 0 15960 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 16184 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 16296 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_139
timestamp 1698175906
transform 1 0 8456 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_143
timestamp 1698175906
transform 1 0 8680 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_210
timestamp 1698175906
transform 1 0 12432 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_226
timestamp 1698175906
transform 1 0 13328 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 14224 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_174
timestamp 1698175906
transform 1 0 10416 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_190
timestamp 1698175906
transform 1 0 11312 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_198
timestamp 1698175906
transform 1 0 11760 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_204
timestamp 1698175906
transform 1 0 12096 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698175906
transform 1 0 12320 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_203
timestamp 1698175906
transform 1 0 12040 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_211
timestamp 1698175906
transform 1 0 12488 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_215
timestamp 1698175906
transform 1 0 12712 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_243
timestamp 1698175906
transform 1 0 14280 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_174
timestamp 1698175906
transform 1 0 10416 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_201
timestamp 1698175906
transform 1 0 11928 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 14000 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 15792 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 16240 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_164
timestamp 1698175906
transform 1 0 9856 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_168
timestamp 1698175906
transform 1 0 10080 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_266
timestamp 1698175906
transform 1 0 15568 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_270
timestamp 1698175906
transform 1 0 15792 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita17_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19992 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita17_26
timestamp 1698175906
transform -1 0 7672 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 2240 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 18760 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 9464 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 10472 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 18760 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 10472 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 8736 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 12824 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 2240 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform -1 0 2240 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 10640 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13104 400 13160 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 11424 400 11480 0 FreeSans 224 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 11760 0 11816 400 0 FreeSans 224 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 20600 9072 21000 9128 0 FreeSans 224 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 12096 0 12152 400 0 FreeSans 224 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 13104 20600 13160 21000 0 FreeSans 224 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 9408 0 9464 400 0 FreeSans 224 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 12432 20600 12488 21000 0 FreeSans 224 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 7392 0 7448 400 0 FreeSans 224 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 10416 0 10472 400 0 FreeSans 224 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 20600 10416 21000 10472 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 20600 7728 21000 7784 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 20600 8400 21000 8456 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 10416 20600 10472 21000 0 FreeSans 224 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 12096 20600 12152 21000 0 FreeSans 224 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 12768 20600 12824 21000 0 FreeSans 224 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 0 12096 400 12152 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 12432 400 12488 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 7728 20600 7784 21000 0 FreeSans 224 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 8400 400 8456 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 10080 20600 10136 21000 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 10752 20600 10808 21000 0 FreeSans 224 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal3 9268 12068 9268 12068 0 _000_
rlabel metal2 7140 12936 7140 12936 0 _001_
rlabel metal2 6412 12152 6412 12152 0 _002_
rlabel metal2 9940 11676 9940 11676 0 _003_
rlabel metal2 5880 9996 5880 9996 0 _004_
rlabel metal2 6692 10948 6692 10948 0 _005_
rlabel metal2 6580 7728 6580 7728 0 _006_
rlabel metal2 6916 8932 6916 8932 0 _007_
rlabel metal2 8708 12012 8708 12012 0 _008_
rlabel metal2 11928 12796 11928 12796 0 _009_
rlabel metal2 13328 12404 13328 12404 0 _010_
rlabel metal2 11312 13468 11312 13468 0 _011_
rlabel metal2 9548 13468 9548 13468 0 _012_
rlabel metal2 13524 9016 13524 9016 0 _013_
rlabel metal2 12236 11396 12236 11396 0 _014_
rlabel metal2 13412 10080 13412 10080 0 _015_
rlabel metal2 13160 7700 13160 7700 0 _016_
rlabel metal2 13356 8876 13356 8876 0 _017_
rlabel metal2 5936 11228 5936 11228 0 _018_
rlabel metal2 6132 8680 6132 8680 0 _019_
rlabel metal2 13020 11368 13020 11368 0 _020_
rlabel metal2 7700 6636 7700 6636 0 _021_
rlabel metal3 8540 7924 8540 7924 0 _022_
rlabel metal3 9576 6412 9576 6412 0 _023_
rlabel metal2 11200 6524 11200 6524 0 _024_
rlabel metal2 11368 6916 11368 6916 0 _025_
rlabel metal2 7532 9184 7532 9184 0 _026_
rlabel metal3 7084 8820 7084 8820 0 _027_
rlabel metal2 8148 12068 8148 12068 0 _028_
rlabel metal3 12292 13132 12292 13132 0 _029_
rlabel metal2 13580 12712 13580 12712 0 _030_
rlabel metal2 13524 12544 13524 12544 0 _031_
rlabel metal2 11900 11256 11900 11256 0 _032_
rlabel metal2 11480 13804 11480 13804 0 _033_
rlabel metal2 10052 12880 10052 12880 0 _034_
rlabel metal2 12908 8792 12908 8792 0 _035_
rlabel metal2 9324 8820 9324 8820 0 _036_
rlabel metal2 12796 8848 12796 8848 0 _037_
rlabel metal2 13692 10640 13692 10640 0 _038_
rlabel metal2 12964 8876 12964 8876 0 _039_
rlabel metal2 11564 9464 11564 9464 0 _040_
rlabel metal2 11676 10892 11676 10892 0 _041_
rlabel metal2 10892 10920 10892 10920 0 _042_
rlabel metal2 12460 9828 12460 9828 0 _043_
rlabel metal3 13020 10108 13020 10108 0 _044_
rlabel metal3 13860 10892 13860 10892 0 _045_
rlabel metal3 13972 10780 13972 10780 0 _046_
rlabel metal2 13524 10430 13524 10430 0 _047_
rlabel metal3 13678 7924 13678 7924 0 _048_
rlabel metal2 13608 8036 13608 8036 0 _049_
rlabel metal2 5796 11284 5796 11284 0 _050_
rlabel metal3 6916 8764 6916 8764 0 _051_
rlabel metal2 13300 11228 13300 11228 0 _052_
rlabel metal3 9828 6972 9828 6972 0 _053_
rlabel metal2 9100 6468 9100 6468 0 _054_
rlabel metal2 9100 8512 9100 8512 0 _055_
rlabel metal2 9156 8204 9156 8204 0 _056_
rlabel metal2 11508 7056 11508 7056 0 _057_
rlabel metal3 10024 6860 10024 6860 0 _058_
rlabel metal2 10108 7056 10108 7056 0 _059_
rlabel metal2 10752 8148 10752 8148 0 _060_
rlabel metal2 11508 7756 11508 7756 0 _061_
rlabel metal2 11900 7336 11900 7336 0 _062_
rlabel metal2 11228 8232 11228 8232 0 _063_
rlabel metal2 8988 10108 8988 10108 0 _064_
rlabel metal2 11844 11144 11844 11144 0 _065_
rlabel metal2 8456 8820 8456 8820 0 _066_
rlabel metal2 13468 8876 13468 8876 0 _067_
rlabel metal3 8932 7644 8932 7644 0 _068_
rlabel metal3 10472 9548 10472 9548 0 _069_
rlabel metal3 8400 9548 8400 9548 0 _070_
rlabel metal2 11172 9520 11172 9520 0 _071_
rlabel metal2 10052 11312 10052 11312 0 _072_
rlabel metal2 13804 10668 13804 10668 0 _073_
rlabel metal2 8120 11900 8120 11900 0 _074_
rlabel metal2 6636 11928 6636 11928 0 _075_
rlabel metal2 9380 12348 9380 12348 0 _076_
rlabel metal2 11060 8764 11060 8764 0 _077_
rlabel metal2 10220 9940 10220 9940 0 _078_
rlabel metal2 12516 9744 12516 9744 0 _079_
rlabel metal2 6860 11032 6860 11032 0 _080_
rlabel metal2 8316 10500 8316 10500 0 _081_
rlabel metal3 8400 11172 8400 11172 0 _082_
rlabel metal2 8344 11452 8344 11452 0 _083_
rlabel metal3 6412 11060 6412 11060 0 _084_
rlabel metal2 12012 13678 12012 13678 0 _085_
rlabel metal2 7420 12880 7420 12880 0 _086_
rlabel metal2 10500 10472 10500 10472 0 _087_
rlabel metal2 10556 8568 10556 8568 0 _088_
rlabel metal2 6468 11480 6468 11480 0 _089_
rlabel metal2 6104 11956 6104 11956 0 _090_
rlabel metal2 9268 8792 9268 8792 0 _091_
rlabel metal2 10052 12180 10052 12180 0 _092_
rlabel metal2 9604 10584 9604 10584 0 _093_
rlabel metal2 10164 11704 10164 11704 0 _094_
rlabel metal2 7308 8568 7308 8568 0 _095_
rlabel metal2 10276 11256 10276 11256 0 _096_
rlabel metal2 9016 6636 9016 6636 0 _097_
rlabel metal2 9156 9352 9156 9352 0 _098_
rlabel metal2 7028 8708 7028 8708 0 _099_
rlabel metal3 11004 8484 11004 8484 0 _100_
rlabel metal2 11956 9632 11956 9632 0 _101_
rlabel metal3 12656 10836 12656 10836 0 _102_
rlabel metal2 12096 11116 12096 11116 0 _103_
rlabel metal3 1239 13132 1239 13132 0 clk
rlabel metal2 11760 10388 11760 10388 0 clknet_0_clk
rlabel metal2 6356 10864 6356 10864 0 clknet_1_0__leaf_clk
rlabel metal2 11536 13524 11536 13524 0 clknet_1_1__leaf_clk
rlabel metal2 6916 9828 6916 9828 0 dut17.count\[0\]
rlabel metal2 7756 10752 7756 10752 0 dut17.count\[1\]
rlabel metal3 8176 7588 8176 7588 0 dut17.count\[2\]
rlabel metal2 7196 9380 7196 9380 0 dut17.count\[3\]
rlabel metal3 3178 11564 3178 11564 0 net1
rlabel metal2 14812 10388 14812 10388 0 net10
rlabel metal2 14028 7756 14028 7756 0 net11
rlabel metal2 13748 8176 13748 8176 0 net12
rlabel metal2 10388 14770 10388 14770 0 net13
rlabel metal2 14364 11564 14364 11564 0 net14
rlabel metal2 8820 2982 8820 2982 0 net15
rlabel metal2 12348 13804 12348 13804 0 net16
rlabel metal2 14364 12712 14364 12712 0 net17
rlabel metal2 12908 15848 12908 15848 0 net18
rlabel metal2 6972 12320 6972 12320 0 net19
rlabel metal2 12264 6524 12264 6524 0 net2
rlabel metal2 5068 12516 5068 12516 0 net20
rlabel metal3 8288 13244 8288 13244 0 net21
rlabel metal3 3178 8820 3178 8820 0 net22
rlabel metal3 10416 18228 10416 18228 0 net23
rlabel metal2 10836 12264 10836 12264 0 net24
rlabel metal2 20132 11536 20132 11536 0 net25
rlabel metal2 7420 1015 7420 1015 0 net26
rlabel metal2 14588 9352 14588 9352 0 net3
rlabel metal2 18844 11312 18844 11312 0 net4
rlabel metal2 12404 6804 12404 6804 0 net5
rlabel metal3 13776 13468 13776 13468 0 net6
rlabel metal2 9268 7280 9268 7280 0 net7
rlabel metal2 12740 16072 12740 16072 0 net8
rlabel metal2 10556 2982 10556 2982 0 net9
rlabel metal3 679 11452 679 11452 0 segm[0]
rlabel metal2 11788 1099 11788 1099 0 segm[10]
rlabel metal3 20321 9100 20321 9100 0 segm[11]
rlabel metal2 20020 11172 20020 11172 0 segm[12]
rlabel metal2 12124 1211 12124 1211 0 segm[13]
rlabel metal2 13132 19873 13132 19873 0 segm[1]
rlabel metal2 9436 1211 9436 1211 0 segm[3]
rlabel metal2 12460 19677 12460 19677 0 segm[4]
rlabel metal2 10444 1099 10444 1099 0 segm[6]
rlabel metal2 20020 10556 20020 10556 0 segm[7]
rlabel metal2 20020 7924 20020 7924 0 segm[8]
rlabel metal2 20020 8652 20020 8652 0 segm[9]
rlabel metal2 10444 19677 10444 19677 0 sel[0]
rlabel metal2 20020 11900 20020 11900 0 sel[10]
rlabel metal2 9100 1099 9100 1099 0 sel[11]
rlabel metal2 12124 19873 12124 19873 0 sel[1]
rlabel metal2 20020 12908 20020 12908 0 sel[2]
rlabel metal2 12796 20573 12796 20573 0 sel[3]
rlabel metal3 679 12124 679 12124 0 sel[4]
rlabel metal3 679 12460 679 12460 0 sel[5]
rlabel metal2 7756 19873 7756 19873 0 sel[6]
rlabel metal3 679 8428 679 8428 0 sel[7]
rlabel metal2 10108 19481 10108 19481 0 sel[8]
rlabel metal2 10780 19873 10780 19873 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
