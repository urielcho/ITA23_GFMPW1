magic
tech gf180mcuD
magscale 1 10
timestamp 1699641766
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 19182 38274 19234 38286
rect 19182 38210 19234 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 22194 38110 22206 38162
rect 22258 38110 22270 38162
rect 19730 37998 19742 38050
rect 19794 37998 19806 38050
rect 23874 37998 23886 38050
rect 23938 37998 23950 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 18398 37490 18450 37502
rect 18398 37426 18450 37438
rect 21422 37490 21474 37502
rect 21422 37426 21474 37438
rect 26798 37490 26850 37502
rect 26798 37426 26850 37438
rect 17378 37214 17390 37266
rect 17442 37214 17454 37266
rect 20402 37214 20414 37266
rect 20466 37214 20478 37266
rect 25778 37214 25790 37266
rect 25842 37214 25854 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 24782 36706 24834 36718
rect 24782 36642 24834 36654
rect 24210 36430 24222 36482
rect 24274 36430 24286 36482
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 24210 28702 24222 28754
rect 24274 28702 24286 28754
rect 24670 28642 24722 28654
rect 21410 28590 21422 28642
rect 21474 28590 21486 28642
rect 24670 28578 24722 28590
rect 22082 28478 22094 28530
rect 22146 28478 22158 28530
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 22094 28082 22146 28094
rect 22094 28018 22146 28030
rect 21982 27970 22034 27982
rect 21982 27906 22034 27918
rect 22206 27858 22258 27870
rect 17490 27806 17502 27858
rect 17554 27806 17566 27858
rect 22206 27794 22258 27806
rect 23214 27858 23266 27870
rect 23426 27806 23438 27858
rect 23490 27806 23502 27858
rect 23214 27794 23266 27806
rect 20862 27746 20914 27758
rect 18162 27694 18174 27746
rect 18226 27694 18238 27746
rect 20290 27694 20302 27746
rect 20354 27694 20366 27746
rect 20862 27682 20914 27694
rect 23102 27634 23154 27646
rect 23102 27570 23154 27582
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 26238 27186 26290 27198
rect 16370 27134 16382 27186
rect 16434 27134 16446 27186
rect 19618 27134 19630 27186
rect 19682 27134 19694 27186
rect 25778 27134 25790 27186
rect 25842 27134 25854 27186
rect 26238 27122 26290 27134
rect 40014 27186 40066 27198
rect 40014 27122 40066 27134
rect 19854 27074 19906 27086
rect 13570 27022 13582 27074
rect 13634 27022 13646 27074
rect 16818 27022 16830 27074
rect 16882 27022 16894 27074
rect 19854 27010 19906 27022
rect 20190 27074 20242 27086
rect 22866 27022 22878 27074
rect 22930 27022 22942 27074
rect 26898 27022 26910 27074
rect 26962 27022 26974 27074
rect 37650 27022 37662 27074
rect 37714 27022 37726 27074
rect 20190 27010 20242 27022
rect 20078 26962 20130 26974
rect 14242 26910 14254 26962
rect 14306 26910 14318 26962
rect 17490 26910 17502 26962
rect 17554 26910 17566 26962
rect 20078 26898 20130 26910
rect 20526 26962 20578 26974
rect 26574 26962 26626 26974
rect 23650 26910 23662 26962
rect 23714 26910 23726 26962
rect 20526 26898 20578 26910
rect 26574 26898 26626 26910
rect 26686 26850 26738 26862
rect 26686 26786 26738 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 16606 26514 16658 26526
rect 16606 26450 16658 26462
rect 17502 26514 17554 26526
rect 17502 26450 17554 26462
rect 18622 26514 18674 26526
rect 18622 26450 18674 26462
rect 19518 26514 19570 26526
rect 19518 26450 19570 26462
rect 19742 26514 19794 26526
rect 19742 26450 19794 26462
rect 19854 26514 19906 26526
rect 19854 26450 19906 26462
rect 20078 26514 20130 26526
rect 20078 26450 20130 26462
rect 23662 26514 23714 26526
rect 23662 26450 23714 26462
rect 24558 26514 24610 26526
rect 24558 26450 24610 26462
rect 18846 26402 18898 26414
rect 18846 26338 18898 26350
rect 17614 26290 17666 26302
rect 17614 26226 17666 26238
rect 18062 26290 18114 26302
rect 18062 26226 18114 26238
rect 18398 26290 18450 26302
rect 18398 26226 18450 26238
rect 19070 26290 19122 26302
rect 19070 26226 19122 26238
rect 19406 26290 19458 26302
rect 19406 26226 19458 26238
rect 20190 26290 20242 26302
rect 23550 26290 23602 26302
rect 23314 26238 23326 26290
rect 23378 26238 23390 26290
rect 20190 26226 20242 26238
rect 23550 26226 23602 26238
rect 23774 26290 23826 26302
rect 24334 26290 24386 26302
rect 23986 26238 23998 26290
rect 24050 26238 24062 26290
rect 23774 26226 23826 26238
rect 24334 26226 24386 26238
rect 24670 26290 24722 26302
rect 25666 26238 25678 26290
rect 25730 26238 25742 26290
rect 24670 26226 24722 26238
rect 20638 26178 20690 26190
rect 28926 26178 28978 26190
rect 26338 26126 26350 26178
rect 26402 26126 26414 26178
rect 28466 26126 28478 26178
rect 28530 26126 28542 26178
rect 20638 26114 20690 26126
rect 28926 26114 28978 26126
rect 17502 26066 17554 26078
rect 17502 26002 17554 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 1934 25618 1986 25630
rect 1934 25554 1986 25566
rect 16718 25618 16770 25630
rect 24110 25618 24162 25630
rect 18722 25566 18734 25618
rect 18786 25566 18798 25618
rect 16718 25554 16770 25566
rect 24110 25554 24162 25566
rect 40014 25618 40066 25630
rect 40014 25554 40066 25566
rect 16606 25506 16658 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 16606 25442 16658 25454
rect 19070 25506 19122 25518
rect 21534 25506 21586 25518
rect 21298 25454 21310 25506
rect 21362 25454 21374 25506
rect 19070 25442 19122 25454
rect 21534 25442 21586 25454
rect 21758 25506 21810 25518
rect 26126 25506 26178 25518
rect 22754 25454 22766 25506
rect 22818 25454 22830 25506
rect 21758 25442 21810 25454
rect 26126 25442 26178 25454
rect 26350 25506 26402 25518
rect 26562 25454 26574 25506
rect 26626 25454 26638 25506
rect 37650 25454 37662 25506
rect 37714 25454 37726 25506
rect 26350 25442 26402 25454
rect 16942 25394 16994 25406
rect 16942 25330 16994 25342
rect 17166 25394 17218 25406
rect 22978 25342 22990 25394
rect 23042 25342 23054 25394
rect 17166 25330 17218 25342
rect 18510 25282 18562 25294
rect 18510 25218 18562 25230
rect 18734 25282 18786 25294
rect 18734 25218 18786 25230
rect 21422 25282 21474 25294
rect 21422 25218 21474 25230
rect 26462 25282 26514 25294
rect 26462 25218 26514 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 15710 24946 15762 24958
rect 23214 24946 23266 24958
rect 17938 24894 17950 24946
rect 18002 24894 18014 24946
rect 15710 24882 15762 24894
rect 23214 24882 23266 24894
rect 26350 24946 26402 24958
rect 26350 24882 26402 24894
rect 23662 24834 23714 24846
rect 23662 24770 23714 24782
rect 30158 24834 30210 24846
rect 30158 24770 30210 24782
rect 15486 24722 15538 24734
rect 14354 24670 14366 24722
rect 14418 24670 14430 24722
rect 15138 24670 15150 24722
rect 15202 24670 15214 24722
rect 15486 24658 15538 24670
rect 15822 24722 15874 24734
rect 15822 24658 15874 24670
rect 17950 24722 18002 24734
rect 17950 24658 18002 24670
rect 18174 24722 18226 24734
rect 18174 24658 18226 24670
rect 18398 24722 18450 24734
rect 18398 24658 18450 24670
rect 18622 24722 18674 24734
rect 22990 24722 23042 24734
rect 19842 24670 19854 24722
rect 19906 24670 19918 24722
rect 18622 24658 18674 24670
rect 22990 24658 23042 24670
rect 23438 24722 23490 24734
rect 26226 24670 26238 24722
rect 26290 24670 26302 24722
rect 26898 24670 26910 24722
rect 26962 24670 26974 24722
rect 23438 24658 23490 24670
rect 16270 24610 16322 24622
rect 12226 24558 12238 24610
rect 12290 24558 12302 24610
rect 16270 24546 16322 24558
rect 19518 24610 19570 24622
rect 25902 24610 25954 24622
rect 20626 24558 20638 24610
rect 20690 24558 20702 24610
rect 22754 24558 22766 24610
rect 22818 24558 22830 24610
rect 27570 24558 27582 24610
rect 27634 24558 27646 24610
rect 29698 24558 29710 24610
rect 29762 24558 29774 24610
rect 19518 24546 19570 24558
rect 25902 24546 25954 24558
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 24882 24110 24894 24162
rect 24946 24110 24958 24162
rect 1934 24050 1986 24062
rect 14030 24050 14082 24062
rect 9986 23998 9998 24050
rect 10050 23998 10062 24050
rect 1934 23986 1986 23998
rect 14030 23986 14082 23998
rect 15710 24050 15762 24062
rect 15710 23986 15762 23998
rect 23662 24050 23714 24062
rect 23662 23986 23714 23998
rect 26574 24050 26626 24062
rect 26574 23986 26626 23998
rect 15486 23938 15538 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 12898 23886 12910 23938
rect 12962 23886 12974 23938
rect 14802 23886 14814 23938
rect 14866 23886 14878 23938
rect 15486 23874 15538 23886
rect 15598 23938 15650 23950
rect 15598 23874 15650 23886
rect 17726 23938 17778 23950
rect 17726 23874 17778 23886
rect 23774 23938 23826 23950
rect 23774 23874 23826 23886
rect 24110 23938 24162 23950
rect 25118 23938 25170 23950
rect 24658 23886 24670 23938
rect 24722 23886 24734 23938
rect 24110 23874 24162 23886
rect 25118 23874 25170 23886
rect 27134 23938 27186 23950
rect 27134 23874 27186 23886
rect 28142 23938 28194 23950
rect 28142 23874 28194 23886
rect 28478 23938 28530 23950
rect 28478 23874 28530 23886
rect 13470 23826 13522 23838
rect 12114 23774 12126 23826
rect 12178 23774 12190 23826
rect 13470 23762 13522 23774
rect 13582 23826 13634 23838
rect 13582 23762 13634 23774
rect 16046 23826 16098 23838
rect 16046 23762 16098 23774
rect 17390 23826 17442 23838
rect 17390 23762 17442 23774
rect 23550 23826 23602 23838
rect 23550 23762 23602 23774
rect 25454 23826 25506 23838
rect 25454 23762 25506 23774
rect 28366 23826 28418 23838
rect 28366 23762 28418 23774
rect 15038 23714 15090 23726
rect 15038 23650 15090 23662
rect 15822 23714 15874 23726
rect 15822 23650 15874 23662
rect 16718 23714 16770 23726
rect 16718 23650 16770 23662
rect 17502 23714 17554 23726
rect 17502 23650 17554 23662
rect 25342 23714 25394 23726
rect 25342 23650 25394 23662
rect 26462 23714 26514 23726
rect 26462 23650 26514 23662
rect 26686 23714 26738 23726
rect 26686 23650 26738 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 21646 23378 21698 23390
rect 26462 23378 26514 23390
rect 17378 23326 17390 23378
rect 17442 23326 17454 23378
rect 24546 23326 24558 23378
rect 24610 23326 24622 23378
rect 21646 23314 21698 23326
rect 26462 23314 26514 23326
rect 30830 23378 30882 23390
rect 30830 23314 30882 23326
rect 20974 23266 21026 23278
rect 15698 23214 15710 23266
rect 15762 23214 15774 23266
rect 20974 23202 21026 23214
rect 22206 23266 22258 23278
rect 22206 23202 22258 23214
rect 22654 23266 22706 23278
rect 23650 23214 23662 23266
rect 23714 23214 23726 23266
rect 22654 23202 22706 23214
rect 17726 23154 17778 23166
rect 4274 23102 4286 23154
rect 4338 23102 4350 23154
rect 16482 23102 16494 23154
rect 16546 23102 16558 23154
rect 17726 23090 17778 23102
rect 20862 23154 20914 23166
rect 20862 23090 20914 23102
rect 21198 23154 21250 23166
rect 22094 23154 22146 23166
rect 21410 23102 21422 23154
rect 21474 23102 21486 23154
rect 21198 23090 21250 23102
rect 22094 23090 22146 23102
rect 23214 23154 23266 23166
rect 26238 23154 26290 23166
rect 23538 23102 23550 23154
rect 23602 23102 23614 23154
rect 24546 23102 24558 23154
rect 24610 23102 24622 23154
rect 26002 23102 26014 23154
rect 26066 23102 26078 23154
rect 23214 23090 23266 23102
rect 26238 23090 26290 23102
rect 26574 23154 26626 23166
rect 27010 23102 27022 23154
rect 27074 23102 27086 23154
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 26574 23090 26626 23102
rect 26350 23042 26402 23054
rect 30382 23042 30434 23054
rect 13570 22990 13582 23042
rect 13634 22990 13646 23042
rect 27794 22990 27806 23042
rect 27858 22990 27870 23042
rect 29922 22990 29934 23042
rect 29986 22990 29998 23042
rect 26350 22978 26402 22990
rect 30382 22978 30434 22990
rect 1934 22930 1986 22942
rect 1934 22866 1986 22878
rect 21758 22930 21810 22942
rect 21758 22866 21810 22878
rect 22206 22930 22258 22942
rect 22206 22866 22258 22878
rect 30270 22930 30322 22942
rect 30270 22866 30322 22878
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 26910 22594 26962 22606
rect 26910 22530 26962 22542
rect 40014 22482 40066 22494
rect 14466 22430 14478 22482
rect 14530 22430 14542 22482
rect 16818 22430 16830 22482
rect 16882 22430 16894 22482
rect 28466 22430 28478 22482
rect 28530 22430 28542 22482
rect 29922 22430 29934 22482
rect 29986 22430 29998 22482
rect 32050 22430 32062 22482
rect 32114 22430 32126 22482
rect 40014 22418 40066 22430
rect 14590 22370 14642 22382
rect 19294 22370 19346 22382
rect 16482 22318 16494 22370
rect 16546 22318 16558 22370
rect 17602 22318 17614 22370
rect 17666 22318 17678 22370
rect 14590 22306 14642 22318
rect 19294 22306 19346 22318
rect 19518 22370 19570 22382
rect 28030 22370 28082 22382
rect 20738 22318 20750 22370
rect 20802 22318 20814 22370
rect 21746 22318 21758 22370
rect 21810 22318 21822 22370
rect 23986 22318 23998 22370
rect 24050 22318 24062 22370
rect 27234 22318 27246 22370
rect 27298 22318 27310 22370
rect 19518 22306 19570 22318
rect 28030 22306 28082 22318
rect 28366 22370 28418 22382
rect 28578 22318 28590 22370
rect 28642 22318 28654 22370
rect 29250 22318 29262 22370
rect 29314 22318 29326 22370
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 28366 22306 28418 22318
rect 15038 22258 15090 22270
rect 16034 22206 16046 22258
rect 16098 22206 16110 22258
rect 17490 22206 17502 22258
rect 17554 22206 17566 22258
rect 19842 22206 19854 22258
rect 19906 22206 19918 22258
rect 20402 22206 20414 22258
rect 20466 22206 20478 22258
rect 21410 22206 21422 22258
rect 21474 22206 21486 22258
rect 23874 22206 23886 22258
rect 23938 22206 23950 22258
rect 25218 22206 25230 22258
rect 25282 22206 25294 22258
rect 26562 22206 26574 22258
rect 26626 22206 26638 22258
rect 15038 22194 15090 22206
rect 14478 22146 14530 22158
rect 14478 22082 14530 22094
rect 14814 22146 14866 22158
rect 14814 22082 14866 22094
rect 18734 22146 18786 22158
rect 24894 22146 24946 22158
rect 23314 22094 23326 22146
rect 23378 22094 23390 22146
rect 18734 22082 18786 22094
rect 24894 22082 24946 22094
rect 25566 22146 25618 22158
rect 26238 22146 26290 22158
rect 25890 22094 25902 22146
rect 25954 22094 25966 22146
rect 25566 22082 25618 22094
rect 26238 22082 26290 22094
rect 27022 22146 27074 22158
rect 27022 22082 27074 22094
rect 28142 22146 28194 22158
rect 28142 22082 28194 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 13134 21810 13186 21822
rect 13134 21746 13186 21758
rect 16382 21810 16434 21822
rect 16382 21746 16434 21758
rect 23550 21810 23602 21822
rect 23550 21746 23602 21758
rect 23662 21810 23714 21822
rect 23662 21746 23714 21758
rect 28814 21810 28866 21822
rect 28814 21746 28866 21758
rect 29038 21810 29090 21822
rect 29038 21746 29090 21758
rect 29598 21810 29650 21822
rect 29598 21746 29650 21758
rect 30046 21810 30098 21822
rect 30046 21746 30098 21758
rect 15934 21698 15986 21710
rect 18498 21646 18510 21698
rect 18562 21646 18574 21698
rect 24098 21646 24110 21698
rect 24162 21646 24174 21698
rect 15934 21634 15986 21646
rect 16270 21586 16322 21598
rect 4274 21534 4286 21586
rect 4338 21534 4350 21586
rect 16270 21522 16322 21534
rect 16606 21586 16658 21598
rect 23774 21586 23826 21598
rect 22642 21534 22654 21586
rect 22706 21534 22718 21586
rect 22978 21534 22990 21586
rect 23042 21534 23054 21586
rect 23314 21534 23326 21586
rect 23378 21534 23390 21586
rect 16606 21522 16658 21534
rect 23774 21522 23826 21534
rect 24446 21586 24498 21598
rect 29150 21586 29202 21598
rect 25666 21534 25678 21586
rect 25730 21534 25742 21586
rect 24446 21522 24498 21534
rect 29150 21522 29202 21534
rect 26450 21422 26462 21474
rect 26514 21422 26526 21474
rect 28578 21422 28590 21474
rect 28642 21422 28654 21474
rect 1934 21362 1986 21374
rect 1934 21298 1986 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 13806 21026 13858 21038
rect 13806 20962 13858 20974
rect 30158 21026 30210 21038
rect 30158 20962 30210 20974
rect 18846 20914 18898 20926
rect 40014 20914 40066 20926
rect 2034 20862 2046 20914
rect 2098 20862 2110 20914
rect 9986 20862 9998 20914
rect 10050 20862 10062 20914
rect 18162 20862 18174 20914
rect 18226 20862 18238 20914
rect 20290 20862 20302 20914
rect 20354 20862 20366 20914
rect 18846 20850 18898 20862
rect 40014 20850 40066 20862
rect 13918 20802 13970 20814
rect 4274 20750 4286 20802
rect 4338 20750 4350 20802
rect 12898 20750 12910 20802
rect 12962 20750 12974 20802
rect 13458 20750 13470 20802
rect 13522 20750 13534 20802
rect 13918 20738 13970 20750
rect 14254 20802 14306 20814
rect 14254 20738 14306 20750
rect 14814 20802 14866 20814
rect 14814 20738 14866 20750
rect 15038 20802 15090 20814
rect 17950 20802 18002 20814
rect 15250 20750 15262 20802
rect 15314 20750 15326 20802
rect 15038 20738 15090 20750
rect 17950 20738 18002 20750
rect 18734 20802 18786 20814
rect 29822 20802 29874 20814
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 21410 20750 21422 20802
rect 21474 20750 21486 20802
rect 37650 20750 37662 20802
rect 37714 20750 37726 20802
rect 18734 20738 18786 20750
rect 29822 20738 29874 20750
rect 14590 20690 14642 20702
rect 17278 20690 17330 20702
rect 26910 20690 26962 20702
rect 12114 20638 12126 20690
rect 12178 20638 12190 20690
rect 16930 20638 16942 20690
rect 16994 20638 17006 20690
rect 19730 20638 19742 20690
rect 19794 20638 19806 20690
rect 25106 20638 25118 20690
rect 25170 20638 25182 20690
rect 14590 20626 14642 20638
rect 17278 20626 17330 20638
rect 26910 20626 26962 20638
rect 27134 20690 27186 20702
rect 27134 20626 27186 20638
rect 30046 20690 30098 20702
rect 30046 20626 30098 20638
rect 14926 20578 14978 20590
rect 13794 20526 13806 20578
rect 13858 20526 13870 20578
rect 14926 20514 14978 20526
rect 18286 20578 18338 20590
rect 18286 20514 18338 20526
rect 18958 20578 19010 20590
rect 18958 20514 19010 20526
rect 19182 20578 19234 20590
rect 19182 20514 19234 20526
rect 20862 20578 20914 20590
rect 20862 20514 20914 20526
rect 27022 20578 27074 20590
rect 27022 20514 27074 20526
rect 29150 20578 29202 20590
rect 29150 20514 29202 20526
rect 29262 20578 29314 20590
rect 29262 20514 29314 20526
rect 29374 20578 29426 20590
rect 29374 20514 29426 20526
rect 30158 20578 30210 20590
rect 30158 20514 30210 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 14478 20242 14530 20254
rect 23438 20242 23490 20254
rect 15586 20190 15598 20242
rect 15650 20190 15662 20242
rect 14478 20178 14530 20190
rect 23438 20178 23490 20190
rect 13470 20130 13522 20142
rect 12226 20078 12238 20130
rect 12290 20078 12302 20130
rect 13470 20066 13522 20078
rect 14366 20130 14418 20142
rect 14366 20066 14418 20078
rect 14590 20130 14642 20142
rect 14590 20066 14642 20078
rect 16718 20130 16770 20142
rect 17602 20078 17614 20130
rect 17666 20078 17678 20130
rect 30034 20078 30046 20130
rect 30098 20078 30110 20130
rect 16718 20066 16770 20078
rect 16606 20018 16658 20030
rect 4274 19966 4286 20018
rect 4338 19966 4350 20018
rect 12898 19966 12910 20018
rect 12962 19966 12974 20018
rect 15810 19966 15822 20018
rect 15874 19966 15886 20018
rect 16606 19954 16658 19966
rect 16942 20018 16994 20030
rect 16942 19954 16994 19966
rect 17390 20018 17442 20030
rect 20974 20018 21026 20030
rect 17938 19966 17950 20018
rect 18002 19966 18014 20018
rect 18610 19966 18622 20018
rect 18674 19966 18686 20018
rect 19394 19966 19406 20018
rect 19458 19966 19470 20018
rect 20514 19966 20526 20018
rect 20578 19966 20590 20018
rect 21858 19966 21870 20018
rect 21922 19966 21934 20018
rect 22194 19966 22206 20018
rect 22258 19966 22270 20018
rect 22418 19966 22430 20018
rect 22482 19966 22494 20018
rect 23538 19966 23550 20018
rect 23602 19966 23614 20018
rect 23986 19966 23998 20018
rect 24050 19966 24062 20018
rect 25218 19966 25230 20018
rect 25282 19966 25294 20018
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 17390 19954 17442 19966
rect 20974 19954 21026 19966
rect 13694 19906 13746 19918
rect 10098 19854 10110 19906
rect 10162 19854 10174 19906
rect 13346 19854 13358 19906
rect 13410 19854 13422 19906
rect 19282 19854 19294 19906
rect 19346 19854 19358 19906
rect 13694 19842 13746 19854
rect 1934 19794 1986 19806
rect 40014 19794 40066 19806
rect 17714 19742 17726 19794
rect 17778 19742 17790 19794
rect 19842 19742 19854 19794
rect 19906 19742 19918 19794
rect 21410 19742 21422 19794
rect 21474 19742 21486 19794
rect 22194 19742 22206 19794
rect 22258 19791 22270 19794
rect 22418 19791 22430 19794
rect 22258 19745 22430 19791
rect 22258 19742 22270 19745
rect 22418 19742 22430 19745
rect 22482 19742 22494 19794
rect 1934 19730 1986 19742
rect 40014 19730 40066 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 13582 19458 13634 19470
rect 26574 19458 26626 19470
rect 19170 19406 19182 19458
rect 19234 19406 19246 19458
rect 13582 19394 13634 19406
rect 26574 19394 26626 19406
rect 14030 19346 14082 19358
rect 17278 19346 17330 19358
rect 20750 19346 20802 19358
rect 16482 19294 16494 19346
rect 16546 19294 16558 19346
rect 18834 19294 18846 19346
rect 18898 19294 18910 19346
rect 14030 19282 14082 19294
rect 17278 19282 17330 19294
rect 20750 19282 20802 19294
rect 23774 19346 23826 19358
rect 29922 19294 29934 19346
rect 29986 19294 29998 19346
rect 32050 19294 32062 19346
rect 32114 19294 32126 19346
rect 23774 19282 23826 19294
rect 13470 19234 13522 19246
rect 17390 19234 17442 19246
rect 19630 19234 19682 19246
rect 12786 19182 12798 19234
rect 12850 19182 12862 19234
rect 16146 19182 16158 19234
rect 16210 19182 16222 19234
rect 18610 19182 18622 19234
rect 18674 19182 18686 19234
rect 18946 19182 18958 19234
rect 19010 19182 19022 19234
rect 13470 19170 13522 19182
rect 17390 19170 17442 19182
rect 19630 19170 19682 19182
rect 19966 19234 20018 19246
rect 25790 19234 25842 19246
rect 26462 19234 26514 19246
rect 20290 19182 20302 19234
rect 20354 19182 20366 19234
rect 21746 19182 21758 19234
rect 21810 19182 21822 19234
rect 24882 19182 24894 19234
rect 24946 19182 24958 19234
rect 25554 19182 25566 19234
rect 25618 19182 25630 19234
rect 25890 19182 25902 19234
rect 25954 19182 25966 19234
rect 19966 19170 20018 19182
rect 25790 19170 25842 19182
rect 26462 19170 26514 19182
rect 27022 19234 27074 19246
rect 27022 19170 27074 19182
rect 28030 19234 28082 19246
rect 28030 19170 28082 19182
rect 28590 19234 28642 19246
rect 29250 19182 29262 19234
rect 29314 19182 29326 19234
rect 28590 19170 28642 19182
rect 17614 19122 17666 19134
rect 26238 19122 26290 19134
rect 12562 19070 12574 19122
rect 12626 19070 12638 19122
rect 16706 19070 16718 19122
rect 16770 19070 16782 19122
rect 21410 19070 21422 19122
rect 21474 19070 21486 19122
rect 24658 19070 24670 19122
rect 24722 19070 24734 19122
rect 17614 19058 17666 19070
rect 26238 19058 26290 19070
rect 27694 19122 27746 19134
rect 27694 19058 27746 19070
rect 27918 19122 27970 19134
rect 27918 19058 27970 19070
rect 17166 19010 17218 19022
rect 17166 18946 17218 18958
rect 19742 19010 19794 19022
rect 24334 19010 24386 19022
rect 21970 18958 21982 19010
rect 22034 18958 22046 19010
rect 19742 18946 19794 18958
rect 24334 18946 24386 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 15598 18674 15650 18686
rect 15598 18610 15650 18622
rect 20638 18674 20690 18686
rect 21634 18622 21646 18674
rect 21698 18622 21710 18674
rect 22866 18622 22878 18674
rect 22930 18622 22942 18674
rect 20638 18610 20690 18622
rect 15374 18562 15426 18574
rect 15374 18498 15426 18510
rect 19070 18562 19122 18574
rect 25342 18562 25394 18574
rect 19730 18510 19742 18562
rect 19794 18510 19806 18562
rect 20178 18510 20190 18562
rect 20242 18510 20254 18562
rect 21298 18510 21310 18562
rect 21362 18510 21374 18562
rect 21746 18510 21758 18562
rect 21810 18510 21822 18562
rect 19070 18498 19122 18510
rect 25342 18498 25394 18510
rect 25454 18562 25506 18574
rect 25454 18498 25506 18510
rect 27134 18562 27186 18574
rect 27134 18498 27186 18510
rect 27246 18562 27298 18574
rect 27246 18498 27298 18510
rect 15262 18450 15314 18462
rect 15262 18386 15314 18398
rect 16158 18450 16210 18462
rect 16158 18386 16210 18398
rect 17950 18450 18002 18462
rect 17950 18386 18002 18398
rect 18286 18450 18338 18462
rect 18286 18386 18338 18398
rect 19294 18450 19346 18462
rect 19294 18386 19346 18398
rect 22094 18450 22146 18462
rect 22094 18386 22146 18398
rect 22542 18450 22594 18462
rect 22542 18386 22594 18398
rect 23326 18450 23378 18462
rect 23326 18386 23378 18398
rect 23886 18450 23938 18462
rect 23886 18386 23938 18398
rect 25790 18450 25842 18462
rect 25790 18386 25842 18398
rect 27470 18450 27522 18462
rect 27470 18386 27522 18398
rect 27806 18450 27858 18462
rect 27806 18386 27858 18398
rect 16046 18338 16098 18350
rect 16046 18274 16098 18286
rect 17390 18338 17442 18350
rect 17390 18274 17442 18286
rect 18846 18338 18898 18350
rect 18846 18274 18898 18286
rect 20750 18338 20802 18350
rect 20750 18274 20802 18286
rect 25902 18338 25954 18350
rect 25902 18274 25954 18286
rect 25342 18226 25394 18238
rect 25342 18162 25394 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 24222 17890 24274 17902
rect 24222 17826 24274 17838
rect 15262 17778 15314 17790
rect 17726 17778 17778 17790
rect 17378 17726 17390 17778
rect 17442 17726 17454 17778
rect 15262 17714 15314 17726
rect 17726 17714 17778 17726
rect 20190 17778 20242 17790
rect 20190 17714 20242 17726
rect 20414 17778 20466 17790
rect 20414 17714 20466 17726
rect 22990 17778 23042 17790
rect 40014 17778 40066 17790
rect 24658 17726 24670 17778
rect 24722 17726 24734 17778
rect 26786 17726 26798 17778
rect 26850 17726 26862 17778
rect 22990 17714 23042 17726
rect 40014 17714 40066 17726
rect 19070 17666 19122 17678
rect 21646 17666 21698 17678
rect 16930 17614 16942 17666
rect 16994 17614 17006 17666
rect 19842 17614 19854 17666
rect 19906 17614 19918 17666
rect 21410 17614 21422 17666
rect 21474 17614 21486 17666
rect 19070 17602 19122 17614
rect 21646 17602 21698 17614
rect 22430 17666 22482 17678
rect 28142 17666 28194 17678
rect 27458 17614 27470 17666
rect 27522 17614 27534 17666
rect 22430 17602 22482 17614
rect 28142 17602 28194 17614
rect 28366 17666 28418 17678
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 28366 17602 28418 17614
rect 14814 17554 14866 17566
rect 24222 17554 24274 17566
rect 16034 17502 16046 17554
rect 16098 17502 16110 17554
rect 14814 17490 14866 17502
rect 24222 17490 24274 17502
rect 24334 17554 24386 17566
rect 24334 17490 24386 17502
rect 27918 17554 27970 17566
rect 27918 17490 27970 17502
rect 14478 17442 14530 17454
rect 14478 17378 14530 17390
rect 15710 17442 15762 17454
rect 19182 17442 19234 17454
rect 16706 17390 16718 17442
rect 16770 17390 16782 17442
rect 15710 17378 15762 17390
rect 19182 17378 19234 17390
rect 19406 17442 19458 17454
rect 19406 17378 19458 17390
rect 21982 17442 22034 17454
rect 21982 17378 22034 17390
rect 28030 17442 28082 17454
rect 28030 17378 28082 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 17950 17106 18002 17118
rect 17950 17042 18002 17054
rect 20078 17106 20130 17118
rect 20078 17042 20130 17054
rect 20302 17106 20354 17118
rect 20302 17042 20354 17054
rect 21198 17106 21250 17118
rect 21198 17042 21250 17054
rect 21310 17106 21362 17118
rect 21310 17042 21362 17054
rect 21870 17106 21922 17118
rect 21870 17042 21922 17054
rect 22654 17106 22706 17118
rect 22654 17042 22706 17054
rect 23326 17106 23378 17118
rect 24334 17106 24386 17118
rect 23650 17054 23662 17106
rect 23714 17054 23726 17106
rect 23326 17042 23378 17054
rect 24334 17042 24386 17054
rect 24558 17106 24610 17118
rect 24558 17042 24610 17054
rect 30270 17106 30322 17118
rect 30270 17042 30322 17054
rect 15262 16994 15314 17006
rect 12786 16942 12798 16994
rect 12850 16942 12862 16994
rect 15262 16930 15314 16942
rect 20414 16994 20466 17006
rect 24222 16994 24274 17006
rect 22306 16942 22318 16994
rect 22370 16942 22382 16994
rect 27682 16942 27694 16994
rect 27746 16942 27758 16994
rect 20414 16930 20466 16942
rect 24222 16930 24274 16942
rect 15374 16882 15426 16894
rect 18510 16882 18562 16894
rect 12114 16830 12126 16882
rect 12178 16830 12190 16882
rect 15922 16830 15934 16882
rect 15986 16830 15998 16882
rect 15374 16818 15426 16830
rect 18510 16818 18562 16830
rect 20638 16882 20690 16894
rect 20638 16818 20690 16830
rect 21086 16882 21138 16894
rect 27010 16830 27022 16882
rect 27074 16830 27086 16882
rect 21086 16818 21138 16830
rect 14914 16718 14926 16770
rect 14978 16718 14990 16770
rect 21970 16718 21982 16770
rect 22034 16718 22046 16770
rect 29810 16718 29822 16770
rect 29874 16718 29886 16770
rect 21646 16658 21698 16670
rect 21646 16594 21698 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 14242 16158 14254 16210
rect 14306 16158 14318 16210
rect 16370 16158 16382 16210
rect 16434 16158 16446 16210
rect 16830 16098 16882 16110
rect 13458 16046 13470 16098
rect 13522 16046 13534 16098
rect 16830 16034 16882 16046
rect 21870 16098 21922 16110
rect 21870 16034 21922 16046
rect 22206 16098 22258 16110
rect 22206 16034 22258 16046
rect 19518 15986 19570 15998
rect 19518 15922 19570 15934
rect 21534 15986 21586 15998
rect 21534 15922 21586 15934
rect 19182 15874 19234 15886
rect 19182 15810 19234 15822
rect 19406 15874 19458 15886
rect 19406 15810 19458 15822
rect 21982 15874 22034 15886
rect 21982 15810 22034 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 18062 15538 18114 15550
rect 18062 15474 18114 15486
rect 18174 15538 18226 15550
rect 18174 15474 18226 15486
rect 19854 15538 19906 15550
rect 20526 15538 20578 15550
rect 20178 15486 20190 15538
rect 20242 15486 20254 15538
rect 19854 15474 19906 15486
rect 20526 15474 20578 15486
rect 20862 15538 20914 15550
rect 20862 15474 20914 15486
rect 21646 15538 21698 15550
rect 21646 15474 21698 15486
rect 25678 15538 25730 15550
rect 25678 15474 25730 15486
rect 17502 15426 17554 15438
rect 17502 15362 17554 15374
rect 19294 15426 19346 15438
rect 19294 15362 19346 15374
rect 21198 15426 21250 15438
rect 21198 15362 21250 15374
rect 21758 15426 21810 15438
rect 21758 15362 21810 15374
rect 17950 15314 18002 15326
rect 17950 15250 18002 15262
rect 18398 15314 18450 15326
rect 18398 15250 18450 15262
rect 18622 15314 18674 15326
rect 18622 15250 18674 15262
rect 18846 15314 18898 15326
rect 18846 15250 18898 15262
rect 19070 15314 19122 15326
rect 19070 15250 19122 15262
rect 19406 15314 19458 15326
rect 19406 15250 19458 15262
rect 21422 15314 21474 15326
rect 21422 15250 21474 15262
rect 25566 15314 25618 15326
rect 26686 15314 26738 15326
rect 25778 15262 25790 15314
rect 25842 15262 25854 15314
rect 26898 15262 26910 15314
rect 26962 15262 26974 15314
rect 37650 15262 37662 15314
rect 37714 15262 37726 15314
rect 25566 15250 25618 15262
rect 26686 15250 26738 15262
rect 17390 15202 17442 15214
rect 17390 15138 17442 15150
rect 40014 15202 40066 15214
rect 40014 15138 40066 15150
rect 25342 15090 25394 15102
rect 25342 15026 25394 15038
rect 26574 15090 26626 15102
rect 26574 15026 26626 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 22206 14754 22258 14766
rect 22206 14690 22258 14702
rect 24670 14642 24722 14654
rect 16146 14590 16158 14642
rect 16210 14590 16222 14642
rect 18274 14590 18286 14642
rect 18338 14590 18350 14642
rect 26114 14590 26126 14642
rect 26178 14590 26190 14642
rect 28242 14590 28254 14642
rect 28306 14590 28318 14642
rect 24670 14578 24722 14590
rect 18846 14530 18898 14542
rect 15474 14478 15486 14530
rect 15538 14478 15550 14530
rect 18846 14466 18898 14478
rect 19182 14530 19234 14542
rect 19182 14466 19234 14478
rect 19406 14530 19458 14542
rect 19406 14466 19458 14478
rect 20078 14530 20130 14542
rect 20078 14466 20130 14478
rect 21982 14530 22034 14542
rect 23886 14530 23938 14542
rect 22530 14478 22542 14530
rect 22594 14478 22606 14530
rect 21982 14466 22034 14478
rect 23886 14466 23938 14478
rect 24334 14530 24386 14542
rect 24334 14466 24386 14478
rect 24446 14530 24498 14542
rect 25330 14478 25342 14530
rect 25394 14478 25406 14530
rect 24446 14466 24498 14478
rect 24894 14418 24946 14430
rect 24894 14354 24946 14366
rect 18958 14306 19010 14318
rect 18958 14242 19010 14254
rect 19742 14306 19794 14318
rect 19742 14242 19794 14254
rect 19966 14306 20018 14318
rect 19966 14242 20018 14254
rect 25006 14306 25058 14318
rect 25006 14242 25058 14254
rect 29262 14306 29314 14318
rect 29262 14242 29314 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 18510 13970 18562 13982
rect 18510 13906 18562 13918
rect 28590 13970 28642 13982
rect 28590 13906 28642 13918
rect 24110 13858 24162 13870
rect 19730 13806 19742 13858
rect 19794 13806 19806 13858
rect 24110 13794 24162 13806
rect 24334 13858 24386 13870
rect 24334 13794 24386 13806
rect 24446 13858 24498 13870
rect 26002 13806 26014 13858
rect 26066 13806 26078 13858
rect 24446 13794 24498 13806
rect 23438 13746 23490 13758
rect 18946 13694 18958 13746
rect 19010 13694 19022 13746
rect 23438 13682 23490 13694
rect 23662 13746 23714 13758
rect 23662 13682 23714 13694
rect 23998 13746 24050 13758
rect 25218 13694 25230 13746
rect 25282 13694 25294 13746
rect 23998 13682 24050 13694
rect 22318 13634 22370 13646
rect 21858 13582 21870 13634
rect 21922 13582 21934 13634
rect 22318 13570 22370 13582
rect 23774 13634 23826 13646
rect 28130 13582 28142 13634
rect 28194 13582 28206 13634
rect 23774 13570 23826 13582
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 26238 13186 26290 13198
rect 26238 13122 26290 13134
rect 19742 13074 19794 13086
rect 17042 13022 17054 13074
rect 17106 13022 17118 13074
rect 19170 13022 19182 13074
rect 19234 13022 19246 13074
rect 22978 13022 22990 13074
rect 23042 13022 23054 13074
rect 25106 13022 25118 13074
rect 25170 13022 25182 13074
rect 19742 13010 19794 13022
rect 16258 12910 16270 12962
rect 16322 12910 16334 12962
rect 22306 12910 22318 12962
rect 22370 12910 22382 12962
rect 26350 12850 26402 12862
rect 26350 12786 26402 12798
rect 25454 12738 25506 12750
rect 25778 12686 25790 12738
rect 25842 12686 25854 12738
rect 25454 12674 25506 12686
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 25454 12402 25506 12414
rect 25454 12338 25506 12350
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 19058 4286 19070 4338
rect 19122 4286 19134 4338
rect 25778 4286 25790 4338
rect 25842 4286 25854 4338
rect 20078 4114 20130 4126
rect 20078 4050 20130 4062
rect 26798 4114 26850 4126
rect 26798 4050 26850 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 18622 3666 18674 3678
rect 18622 3602 18674 3614
rect 26126 3666 26178 3678
rect 26126 3602 26178 3614
rect 29374 3666 29426 3678
rect 29374 3602 29426 3614
rect 17602 3502 17614 3554
rect 17666 3502 17678 3554
rect 25218 3502 25230 3554
rect 25282 3502 25294 3554
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 19182 38222 19234 38274
rect 25566 38222 25618 38274
rect 22206 38110 22258 38162
rect 19742 37998 19794 38050
rect 23886 37998 23938 38050
rect 24558 37998 24610 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 18398 37438 18450 37490
rect 21422 37438 21474 37490
rect 26798 37438 26850 37490
rect 17390 37214 17442 37266
rect 20414 37214 20466 37266
rect 25790 37214 25842 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 24782 36654 24834 36706
rect 24222 36430 24274 36482
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 24222 28702 24274 28754
rect 21422 28590 21474 28642
rect 24670 28590 24722 28642
rect 22094 28478 22146 28530
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 22094 28030 22146 28082
rect 21982 27918 22034 27970
rect 17502 27806 17554 27858
rect 22206 27806 22258 27858
rect 23214 27806 23266 27858
rect 23438 27806 23490 27858
rect 18174 27694 18226 27746
rect 20302 27694 20354 27746
rect 20862 27694 20914 27746
rect 23102 27582 23154 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 16382 27134 16434 27186
rect 19630 27134 19682 27186
rect 25790 27134 25842 27186
rect 26238 27134 26290 27186
rect 40014 27134 40066 27186
rect 13582 27022 13634 27074
rect 16830 27022 16882 27074
rect 19854 27022 19906 27074
rect 20190 27022 20242 27074
rect 22878 27022 22930 27074
rect 26910 27022 26962 27074
rect 37662 27022 37714 27074
rect 14254 26910 14306 26962
rect 17502 26910 17554 26962
rect 20078 26910 20130 26962
rect 20526 26910 20578 26962
rect 23662 26910 23714 26962
rect 26574 26910 26626 26962
rect 26686 26798 26738 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 16606 26462 16658 26514
rect 17502 26462 17554 26514
rect 18622 26462 18674 26514
rect 19518 26462 19570 26514
rect 19742 26462 19794 26514
rect 19854 26462 19906 26514
rect 20078 26462 20130 26514
rect 23662 26462 23714 26514
rect 24558 26462 24610 26514
rect 18846 26350 18898 26402
rect 17614 26238 17666 26290
rect 18062 26238 18114 26290
rect 18398 26238 18450 26290
rect 19070 26238 19122 26290
rect 19406 26238 19458 26290
rect 20190 26238 20242 26290
rect 23326 26238 23378 26290
rect 23550 26238 23602 26290
rect 23774 26238 23826 26290
rect 23998 26238 24050 26290
rect 24334 26238 24386 26290
rect 24670 26238 24722 26290
rect 25678 26238 25730 26290
rect 20638 26126 20690 26178
rect 26350 26126 26402 26178
rect 28478 26126 28530 26178
rect 28926 26126 28978 26178
rect 17502 26014 17554 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 1934 25566 1986 25618
rect 16718 25566 16770 25618
rect 18734 25566 18786 25618
rect 24110 25566 24162 25618
rect 40014 25566 40066 25618
rect 4286 25454 4338 25506
rect 16606 25454 16658 25506
rect 19070 25454 19122 25506
rect 21310 25454 21362 25506
rect 21534 25454 21586 25506
rect 21758 25454 21810 25506
rect 22766 25454 22818 25506
rect 26126 25454 26178 25506
rect 26350 25454 26402 25506
rect 26574 25454 26626 25506
rect 37662 25454 37714 25506
rect 16942 25342 16994 25394
rect 17166 25342 17218 25394
rect 22990 25342 23042 25394
rect 18510 25230 18562 25282
rect 18734 25230 18786 25282
rect 21422 25230 21474 25282
rect 26462 25230 26514 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 15710 24894 15762 24946
rect 17950 24894 18002 24946
rect 23214 24894 23266 24946
rect 26350 24894 26402 24946
rect 23662 24782 23714 24834
rect 30158 24782 30210 24834
rect 14366 24670 14418 24722
rect 15150 24670 15202 24722
rect 15486 24670 15538 24722
rect 15822 24670 15874 24722
rect 17950 24670 18002 24722
rect 18174 24670 18226 24722
rect 18398 24670 18450 24722
rect 18622 24670 18674 24722
rect 19854 24670 19906 24722
rect 22990 24670 23042 24722
rect 23438 24670 23490 24722
rect 26238 24670 26290 24722
rect 26910 24670 26962 24722
rect 12238 24558 12290 24610
rect 16270 24558 16322 24610
rect 19518 24558 19570 24610
rect 20638 24558 20690 24610
rect 22766 24558 22818 24610
rect 25902 24558 25954 24610
rect 27582 24558 27634 24610
rect 29710 24558 29762 24610
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 24894 24110 24946 24162
rect 1934 23998 1986 24050
rect 9998 23998 10050 24050
rect 14030 23998 14082 24050
rect 15710 23998 15762 24050
rect 23662 23998 23714 24050
rect 26574 23998 26626 24050
rect 4286 23886 4338 23938
rect 12910 23886 12962 23938
rect 14814 23886 14866 23938
rect 15486 23886 15538 23938
rect 15598 23886 15650 23938
rect 17726 23886 17778 23938
rect 23774 23886 23826 23938
rect 24110 23886 24162 23938
rect 24670 23886 24722 23938
rect 25118 23886 25170 23938
rect 27134 23886 27186 23938
rect 28142 23886 28194 23938
rect 28478 23886 28530 23938
rect 12126 23774 12178 23826
rect 13470 23774 13522 23826
rect 13582 23774 13634 23826
rect 16046 23774 16098 23826
rect 17390 23774 17442 23826
rect 23550 23774 23602 23826
rect 25454 23774 25506 23826
rect 28366 23774 28418 23826
rect 15038 23662 15090 23714
rect 15822 23662 15874 23714
rect 16718 23662 16770 23714
rect 17502 23662 17554 23714
rect 25342 23662 25394 23714
rect 26462 23662 26514 23714
rect 26686 23662 26738 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 17390 23326 17442 23378
rect 21646 23326 21698 23378
rect 24558 23326 24610 23378
rect 26462 23326 26514 23378
rect 30830 23326 30882 23378
rect 15710 23214 15762 23266
rect 20974 23214 21026 23266
rect 22206 23214 22258 23266
rect 22654 23214 22706 23266
rect 23662 23214 23714 23266
rect 4286 23102 4338 23154
rect 16494 23102 16546 23154
rect 17726 23102 17778 23154
rect 20862 23102 20914 23154
rect 21198 23102 21250 23154
rect 21422 23102 21474 23154
rect 22094 23102 22146 23154
rect 23214 23102 23266 23154
rect 23550 23102 23602 23154
rect 24558 23102 24610 23154
rect 26014 23102 26066 23154
rect 26238 23102 26290 23154
rect 26574 23102 26626 23154
rect 27022 23102 27074 23154
rect 37662 23102 37714 23154
rect 13582 22990 13634 23042
rect 26350 22990 26402 23042
rect 27806 22990 27858 23042
rect 29934 22990 29986 23042
rect 30382 22990 30434 23042
rect 1934 22878 1986 22930
rect 21758 22878 21810 22930
rect 22206 22878 22258 22930
rect 30270 22878 30322 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 26910 22542 26962 22594
rect 14478 22430 14530 22482
rect 16830 22430 16882 22482
rect 28478 22430 28530 22482
rect 29934 22430 29986 22482
rect 32062 22430 32114 22482
rect 40014 22430 40066 22482
rect 14590 22318 14642 22370
rect 16494 22318 16546 22370
rect 17614 22318 17666 22370
rect 19294 22318 19346 22370
rect 19518 22318 19570 22370
rect 20750 22318 20802 22370
rect 21758 22318 21810 22370
rect 23998 22318 24050 22370
rect 27246 22318 27298 22370
rect 28030 22318 28082 22370
rect 28366 22318 28418 22370
rect 28590 22318 28642 22370
rect 29262 22318 29314 22370
rect 37662 22318 37714 22370
rect 15038 22206 15090 22258
rect 16046 22206 16098 22258
rect 17502 22206 17554 22258
rect 19854 22206 19906 22258
rect 20414 22206 20466 22258
rect 21422 22206 21474 22258
rect 23886 22206 23938 22258
rect 25230 22206 25282 22258
rect 26574 22206 26626 22258
rect 14478 22094 14530 22146
rect 14814 22094 14866 22146
rect 18734 22094 18786 22146
rect 23326 22094 23378 22146
rect 24894 22094 24946 22146
rect 25566 22094 25618 22146
rect 25902 22094 25954 22146
rect 26238 22094 26290 22146
rect 27022 22094 27074 22146
rect 28142 22094 28194 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 13134 21758 13186 21810
rect 16382 21758 16434 21810
rect 23550 21758 23602 21810
rect 23662 21758 23714 21810
rect 28814 21758 28866 21810
rect 29038 21758 29090 21810
rect 29598 21758 29650 21810
rect 30046 21758 30098 21810
rect 15934 21646 15986 21698
rect 18510 21646 18562 21698
rect 24110 21646 24162 21698
rect 4286 21534 4338 21586
rect 16270 21534 16322 21586
rect 16606 21534 16658 21586
rect 22654 21534 22706 21586
rect 22990 21534 23042 21586
rect 23326 21534 23378 21586
rect 23774 21534 23826 21586
rect 24446 21534 24498 21586
rect 25678 21534 25730 21586
rect 29150 21534 29202 21586
rect 26462 21422 26514 21474
rect 28590 21422 28642 21474
rect 1934 21310 1986 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 13806 20974 13858 21026
rect 30158 20974 30210 21026
rect 2046 20862 2098 20914
rect 9998 20862 10050 20914
rect 18174 20862 18226 20914
rect 18846 20862 18898 20914
rect 20302 20862 20354 20914
rect 40014 20862 40066 20914
rect 4286 20750 4338 20802
rect 12910 20750 12962 20802
rect 13470 20750 13522 20802
rect 13918 20750 13970 20802
rect 14254 20750 14306 20802
rect 14814 20750 14866 20802
rect 15038 20750 15090 20802
rect 15262 20750 15314 20802
rect 17950 20750 18002 20802
rect 18734 20750 18786 20802
rect 20078 20750 20130 20802
rect 21422 20750 21474 20802
rect 29822 20750 29874 20802
rect 37662 20750 37714 20802
rect 12126 20638 12178 20690
rect 14590 20638 14642 20690
rect 16942 20638 16994 20690
rect 17278 20638 17330 20690
rect 19742 20638 19794 20690
rect 25118 20638 25170 20690
rect 26910 20638 26962 20690
rect 27134 20638 27186 20690
rect 30046 20638 30098 20690
rect 13806 20526 13858 20578
rect 14926 20526 14978 20578
rect 18286 20526 18338 20578
rect 18958 20526 19010 20578
rect 19182 20526 19234 20578
rect 20862 20526 20914 20578
rect 27022 20526 27074 20578
rect 29150 20526 29202 20578
rect 29262 20526 29314 20578
rect 29374 20526 29426 20578
rect 30158 20526 30210 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 14478 20190 14530 20242
rect 15598 20190 15650 20242
rect 23438 20190 23490 20242
rect 12238 20078 12290 20130
rect 13470 20078 13522 20130
rect 14366 20078 14418 20130
rect 14590 20078 14642 20130
rect 16718 20078 16770 20130
rect 17614 20078 17666 20130
rect 30046 20078 30098 20130
rect 4286 19966 4338 20018
rect 12910 19966 12962 20018
rect 15822 19966 15874 20018
rect 16606 19966 16658 20018
rect 16942 19966 16994 20018
rect 17390 19966 17442 20018
rect 17950 19966 18002 20018
rect 18622 19966 18674 20018
rect 19406 19966 19458 20018
rect 20526 19966 20578 20018
rect 20974 19966 21026 20018
rect 21870 19966 21922 20018
rect 22206 19966 22258 20018
rect 22430 19966 22482 20018
rect 23550 19966 23602 20018
rect 23998 19966 24050 20018
rect 25230 19966 25282 20018
rect 37662 19966 37714 20018
rect 10110 19854 10162 19906
rect 13358 19854 13410 19906
rect 13694 19854 13746 19906
rect 19294 19854 19346 19906
rect 1934 19742 1986 19794
rect 17726 19742 17778 19794
rect 19854 19742 19906 19794
rect 21422 19742 21474 19794
rect 22206 19742 22258 19794
rect 22430 19742 22482 19794
rect 40014 19742 40066 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 13582 19406 13634 19458
rect 19182 19406 19234 19458
rect 26574 19406 26626 19458
rect 14030 19294 14082 19346
rect 16494 19294 16546 19346
rect 17278 19294 17330 19346
rect 18846 19294 18898 19346
rect 20750 19294 20802 19346
rect 23774 19294 23826 19346
rect 29934 19294 29986 19346
rect 32062 19294 32114 19346
rect 12798 19182 12850 19234
rect 13470 19182 13522 19234
rect 16158 19182 16210 19234
rect 17390 19182 17442 19234
rect 18622 19182 18674 19234
rect 18958 19182 19010 19234
rect 19630 19182 19682 19234
rect 19966 19182 20018 19234
rect 20302 19182 20354 19234
rect 21758 19182 21810 19234
rect 24894 19182 24946 19234
rect 25566 19182 25618 19234
rect 25790 19182 25842 19234
rect 25902 19182 25954 19234
rect 26462 19182 26514 19234
rect 27022 19182 27074 19234
rect 28030 19182 28082 19234
rect 28590 19182 28642 19234
rect 29262 19182 29314 19234
rect 12574 19070 12626 19122
rect 16718 19070 16770 19122
rect 17614 19070 17666 19122
rect 21422 19070 21474 19122
rect 24670 19070 24722 19122
rect 26238 19070 26290 19122
rect 27694 19070 27746 19122
rect 27918 19070 27970 19122
rect 17166 18958 17218 19010
rect 19742 18958 19794 19010
rect 21982 18958 22034 19010
rect 24334 18958 24386 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 15598 18622 15650 18674
rect 20638 18622 20690 18674
rect 21646 18622 21698 18674
rect 22878 18622 22930 18674
rect 15374 18510 15426 18562
rect 19070 18510 19122 18562
rect 19742 18510 19794 18562
rect 20190 18510 20242 18562
rect 21310 18510 21362 18562
rect 21758 18510 21810 18562
rect 25342 18510 25394 18562
rect 25454 18510 25506 18562
rect 27134 18510 27186 18562
rect 27246 18510 27298 18562
rect 15262 18398 15314 18450
rect 16158 18398 16210 18450
rect 17950 18398 18002 18450
rect 18286 18398 18338 18450
rect 19294 18398 19346 18450
rect 22094 18398 22146 18450
rect 22542 18398 22594 18450
rect 23326 18398 23378 18450
rect 23886 18398 23938 18450
rect 25790 18398 25842 18450
rect 27470 18398 27522 18450
rect 27806 18398 27858 18450
rect 16046 18286 16098 18338
rect 17390 18286 17442 18338
rect 18846 18286 18898 18338
rect 20750 18286 20802 18338
rect 25902 18286 25954 18338
rect 25342 18174 25394 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 24222 17838 24274 17890
rect 15262 17726 15314 17778
rect 17390 17726 17442 17778
rect 17726 17726 17778 17778
rect 20190 17726 20242 17778
rect 20414 17726 20466 17778
rect 22990 17726 23042 17778
rect 24670 17726 24722 17778
rect 26798 17726 26850 17778
rect 40014 17726 40066 17778
rect 16942 17614 16994 17666
rect 19070 17614 19122 17666
rect 19854 17614 19906 17666
rect 21422 17614 21474 17666
rect 21646 17614 21698 17666
rect 22430 17614 22482 17666
rect 27470 17614 27522 17666
rect 28142 17614 28194 17666
rect 28366 17614 28418 17666
rect 37662 17614 37714 17666
rect 14814 17502 14866 17554
rect 16046 17502 16098 17554
rect 24222 17502 24274 17554
rect 24334 17502 24386 17554
rect 27918 17502 27970 17554
rect 14478 17390 14530 17442
rect 15710 17390 15762 17442
rect 16718 17390 16770 17442
rect 19182 17390 19234 17442
rect 19406 17390 19458 17442
rect 21982 17390 22034 17442
rect 28030 17390 28082 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 17950 17054 18002 17106
rect 20078 17054 20130 17106
rect 20302 17054 20354 17106
rect 21198 17054 21250 17106
rect 21310 17054 21362 17106
rect 21870 17054 21922 17106
rect 22654 17054 22706 17106
rect 23326 17054 23378 17106
rect 23662 17054 23714 17106
rect 24334 17054 24386 17106
rect 24558 17054 24610 17106
rect 30270 17054 30322 17106
rect 12798 16942 12850 16994
rect 15262 16942 15314 16994
rect 20414 16942 20466 16994
rect 22318 16942 22370 16994
rect 24222 16942 24274 16994
rect 27694 16942 27746 16994
rect 12126 16830 12178 16882
rect 15374 16830 15426 16882
rect 15934 16830 15986 16882
rect 18510 16830 18562 16882
rect 20638 16830 20690 16882
rect 21086 16830 21138 16882
rect 27022 16830 27074 16882
rect 14926 16718 14978 16770
rect 21982 16718 22034 16770
rect 29822 16718 29874 16770
rect 21646 16606 21698 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 14254 16158 14306 16210
rect 16382 16158 16434 16210
rect 13470 16046 13522 16098
rect 16830 16046 16882 16098
rect 21870 16046 21922 16098
rect 22206 16046 22258 16098
rect 19518 15934 19570 15986
rect 21534 15934 21586 15986
rect 19182 15822 19234 15874
rect 19406 15822 19458 15874
rect 21982 15822 22034 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 18062 15486 18114 15538
rect 18174 15486 18226 15538
rect 19854 15486 19906 15538
rect 20190 15486 20242 15538
rect 20526 15486 20578 15538
rect 20862 15486 20914 15538
rect 21646 15486 21698 15538
rect 25678 15486 25730 15538
rect 17502 15374 17554 15426
rect 19294 15374 19346 15426
rect 21198 15374 21250 15426
rect 21758 15374 21810 15426
rect 17950 15262 18002 15314
rect 18398 15262 18450 15314
rect 18622 15262 18674 15314
rect 18846 15262 18898 15314
rect 19070 15262 19122 15314
rect 19406 15262 19458 15314
rect 21422 15262 21474 15314
rect 25566 15262 25618 15314
rect 25790 15262 25842 15314
rect 26686 15262 26738 15314
rect 26910 15262 26962 15314
rect 37662 15262 37714 15314
rect 17390 15150 17442 15202
rect 40014 15150 40066 15202
rect 25342 15038 25394 15090
rect 26574 15038 26626 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 22206 14702 22258 14754
rect 16158 14590 16210 14642
rect 18286 14590 18338 14642
rect 24670 14590 24722 14642
rect 26126 14590 26178 14642
rect 28254 14590 28306 14642
rect 15486 14478 15538 14530
rect 18846 14478 18898 14530
rect 19182 14478 19234 14530
rect 19406 14478 19458 14530
rect 20078 14478 20130 14530
rect 21982 14478 22034 14530
rect 22542 14478 22594 14530
rect 23886 14478 23938 14530
rect 24334 14478 24386 14530
rect 24446 14478 24498 14530
rect 25342 14478 25394 14530
rect 24894 14366 24946 14418
rect 18958 14254 19010 14306
rect 19742 14254 19794 14306
rect 19966 14254 20018 14306
rect 25006 14254 25058 14306
rect 29262 14254 29314 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 18510 13918 18562 13970
rect 28590 13918 28642 13970
rect 19742 13806 19794 13858
rect 24110 13806 24162 13858
rect 24334 13806 24386 13858
rect 24446 13806 24498 13858
rect 26014 13806 26066 13858
rect 18958 13694 19010 13746
rect 23438 13694 23490 13746
rect 23662 13694 23714 13746
rect 23998 13694 24050 13746
rect 25230 13694 25282 13746
rect 21870 13582 21922 13634
rect 22318 13582 22370 13634
rect 23774 13582 23826 13634
rect 28142 13582 28194 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 26238 13134 26290 13186
rect 17054 13022 17106 13074
rect 19182 13022 19234 13074
rect 19742 13022 19794 13074
rect 22990 13022 23042 13074
rect 25118 13022 25170 13074
rect 16270 12910 16322 12962
rect 22318 12910 22370 12962
rect 26350 12798 26402 12850
rect 25454 12686 25506 12738
rect 25790 12686 25842 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 25454 12350 25506 12402
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 19070 4286 19122 4338
rect 25790 4286 25842 4338
rect 20078 4062 20130 4114
rect 26798 4062 26850 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18622 3614 18674 3666
rect 26126 3614 26178 3666
rect 29374 3614 29426 3666
rect 17614 3502 17666 3554
rect 25230 3502 25282 3554
rect 28590 3502 28642 3554
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 16800 41200 16912 42000
rect 19488 41200 19600 42000
rect 20160 41200 20272 42000
rect 22176 41200 22288 42000
rect 22848 41200 22960 42000
rect 23520 41200 23632 42000
rect 25536 41200 25648 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 16828 37492 16884 41200
rect 19180 38276 19236 38286
rect 19516 38276 19572 41200
rect 19180 38274 19572 38276
rect 19180 38222 19182 38274
rect 19234 38222 19572 38274
rect 19180 38220 19572 38222
rect 19180 38210 19236 38220
rect 19740 38052 19796 38062
rect 19628 38050 19796 38052
rect 19628 37998 19742 38050
rect 19794 37998 19796 38050
rect 19628 37996 19796 37998
rect 16828 37426 16884 37436
rect 18396 37492 18452 37502
rect 18396 37398 18452 37436
rect 17388 37266 17444 37278
rect 17388 37214 17390 37266
rect 17442 37214 17444 37266
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4172 28308 4228 28318
rect 1932 25618 1988 25630
rect 1932 25566 1934 25618
rect 1986 25566 1988 25618
rect 1932 24948 1988 25566
rect 1932 24882 1988 24892
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 1932 23538 1988 23548
rect 1932 22932 1988 22942
rect 1932 22838 1988 22876
rect 1932 21362 1988 21374
rect 1932 21310 1934 21362
rect 1986 21310 1988 21362
rect 1932 20916 1988 21310
rect 1932 20850 1988 20860
rect 2044 20914 2100 20926
rect 2044 20862 2046 20914
rect 2098 20862 2100 20914
rect 2044 20244 2100 20862
rect 4172 20580 4228 28252
rect 16828 27748 16884 27758
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 16380 27188 16436 27198
rect 16380 27094 16436 27132
rect 13580 27076 13636 27086
rect 13580 26982 13636 27020
rect 16604 27076 16660 27086
rect 16828 27076 16884 27692
rect 16660 27074 16884 27076
rect 16660 27022 16830 27074
rect 16882 27022 16884 27074
rect 16660 27020 16884 27022
rect 14252 26962 14308 26974
rect 14252 26910 14254 26962
rect 14306 26910 14308 26962
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 14252 25620 14308 26910
rect 16604 26514 16660 27020
rect 16828 27010 16884 27020
rect 17388 27188 17444 37214
rect 17500 27858 17556 27870
rect 17500 27806 17502 27858
rect 17554 27806 17556 27858
rect 17500 27748 17556 27806
rect 17500 27682 17556 27692
rect 18172 27748 18228 27758
rect 18172 27746 18452 27748
rect 18172 27694 18174 27746
rect 18226 27694 18452 27746
rect 18172 27692 18452 27694
rect 18172 27682 18228 27692
rect 16604 26462 16606 26514
rect 16658 26462 16660 26514
rect 16604 26450 16660 26462
rect 17388 26516 17444 27132
rect 17500 26964 17556 26974
rect 17500 26870 17556 26908
rect 18396 26908 18452 27692
rect 19628 27188 19684 37996
rect 19740 37986 19796 37996
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20188 37492 20244 41200
rect 22204 38162 22260 41200
rect 22876 38276 22932 41200
rect 22876 38210 22932 38220
rect 22204 38110 22206 38162
rect 22258 38110 22260 38162
rect 22204 38098 22260 38110
rect 20188 37426 20244 37436
rect 21420 37492 21476 37502
rect 21420 37398 21476 37436
rect 20412 37266 20468 37278
rect 20412 37214 20414 37266
rect 20466 37214 20468 37266
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20412 31948 20468 37214
rect 23548 36708 23604 41200
rect 25564 38612 25620 41200
rect 25564 38546 25620 38556
rect 26796 38612 26852 38622
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 23548 36642 23604 36652
rect 23884 38050 23940 38062
rect 23884 37998 23886 38050
rect 23938 37998 23940 38050
rect 20300 31892 20468 31948
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19516 27186 19684 27188
rect 19516 27134 19630 27186
rect 19682 27134 19684 27186
rect 19516 27132 19684 27134
rect 18844 27076 18900 27086
rect 18732 27020 18844 27076
rect 18396 26852 18676 26908
rect 17500 26516 17556 26526
rect 17388 26514 17556 26516
rect 17388 26462 17502 26514
rect 17554 26462 17556 26514
rect 17388 26460 17556 26462
rect 17500 26450 17556 26460
rect 18620 26514 18676 26852
rect 18620 26462 18622 26514
rect 18674 26462 18676 26514
rect 18620 26450 18676 26462
rect 17612 26292 17668 26302
rect 18060 26292 18116 26302
rect 18396 26292 18452 26302
rect 17612 26290 18116 26292
rect 17612 26238 17614 26290
rect 17666 26238 18062 26290
rect 18114 26238 18116 26290
rect 17612 26236 18116 26238
rect 17612 26226 17668 26236
rect 18060 26180 18116 26236
rect 18060 26114 18116 26124
rect 18172 26290 18452 26292
rect 18172 26238 18398 26290
rect 18450 26238 18452 26290
rect 18172 26236 18452 26238
rect 14252 25554 14308 25564
rect 16604 26068 16660 26078
rect 4284 25508 4340 25518
rect 4284 25414 4340 25452
rect 12236 25508 12292 25518
rect 12236 24610 12292 25452
rect 16604 25506 16660 26012
rect 17500 26068 17556 26078
rect 17500 25974 17556 26012
rect 16716 25620 16772 25630
rect 16716 25526 16772 25564
rect 16604 25454 16606 25506
rect 16658 25454 16660 25506
rect 16604 25442 16660 25454
rect 16940 25394 16996 25406
rect 16940 25342 16942 25394
rect 16994 25342 16996 25394
rect 16940 25284 16996 25342
rect 16940 25218 16996 25228
rect 17164 25394 17220 25406
rect 17164 25342 17166 25394
rect 17218 25342 17220 25394
rect 15708 25172 15764 25182
rect 15708 24946 15764 25116
rect 15708 24894 15710 24946
rect 15762 24894 15764 24946
rect 15708 24882 15764 24894
rect 14364 24724 14420 24734
rect 14364 24630 14420 24668
rect 15148 24722 15204 24734
rect 15148 24670 15150 24722
rect 15202 24670 15204 24722
rect 12236 24558 12238 24610
rect 12290 24558 12292 24610
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 9996 24050 10052 24062
rect 9996 23998 9998 24050
rect 10050 23998 10052 24050
rect 4284 23940 4340 23950
rect 4284 23846 4340 23884
rect 9996 23940 10052 23998
rect 9996 23604 10052 23884
rect 12236 23940 12292 24558
rect 14028 24612 14084 24622
rect 13132 24052 13188 24062
rect 12236 23874 12292 23884
rect 12908 23940 12964 23950
rect 13132 23940 13188 23996
rect 14028 24052 14084 24556
rect 15148 24612 15204 24670
rect 15484 24724 15540 24734
rect 15484 24630 15540 24668
rect 15820 24722 15876 24734
rect 15820 24670 15822 24722
rect 15874 24670 15876 24722
rect 15148 24546 15204 24556
rect 14028 23958 14084 23996
rect 14700 24052 14756 24062
rect 12908 23938 13188 23940
rect 12908 23886 12910 23938
rect 12962 23886 13188 23938
rect 12908 23884 13188 23886
rect 12908 23874 12964 23884
rect 12124 23828 12180 23838
rect 12124 23734 12180 23772
rect 9996 23538 10052 23548
rect 4284 23156 4340 23166
rect 4284 23062 4340 23100
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 13132 21812 13188 23884
rect 13468 23828 13524 23838
rect 13468 23734 13524 23772
rect 13580 23828 13636 23838
rect 13580 23826 14532 23828
rect 13580 23774 13582 23826
rect 13634 23774 14532 23826
rect 13580 23772 14532 23774
rect 13580 23762 13636 23772
rect 13580 23156 13636 23166
rect 13580 23042 13636 23100
rect 13580 22990 13582 23042
rect 13634 22990 13636 23042
rect 13580 22978 13636 22990
rect 14476 22482 14532 23772
rect 14476 22430 14478 22482
rect 14530 22430 14532 22482
rect 14476 22418 14532 22430
rect 14588 23604 14644 23614
rect 14588 22370 14644 23548
rect 14588 22318 14590 22370
rect 14642 22318 14644 22370
rect 14588 22306 14644 22318
rect 14476 22148 14532 22158
rect 14700 22148 14756 23996
rect 15484 24052 15540 24062
rect 14812 23938 14868 23950
rect 14812 23886 14814 23938
rect 14866 23886 14868 23938
rect 14812 22484 14868 23886
rect 15484 23938 15540 23996
rect 15708 24052 15764 24062
rect 15820 24052 15876 24670
rect 15708 24050 15876 24052
rect 15708 23998 15710 24050
rect 15762 23998 15876 24050
rect 15708 23996 15876 23998
rect 16268 24612 16324 24622
rect 15708 23986 15764 23996
rect 15484 23886 15486 23938
rect 15538 23886 15540 23938
rect 15484 23874 15540 23886
rect 15596 23940 15652 23950
rect 15596 23846 15652 23884
rect 16044 23826 16100 23838
rect 16044 23774 16046 23826
rect 16098 23774 16100 23826
rect 15036 23714 15092 23726
rect 15036 23662 15038 23714
rect 15090 23662 15092 23714
rect 15036 23268 15092 23662
rect 15820 23716 15876 23726
rect 16044 23716 16100 23774
rect 15820 23714 15988 23716
rect 15820 23662 15822 23714
rect 15874 23662 15988 23714
rect 15820 23660 15988 23662
rect 15820 23650 15876 23660
rect 15036 23202 15092 23212
rect 15708 23268 15764 23278
rect 15708 23174 15764 23212
rect 14812 22418 14868 22428
rect 15820 23156 15876 23166
rect 14924 22260 14980 22270
rect 14476 22146 14756 22148
rect 14476 22094 14478 22146
rect 14530 22094 14756 22146
rect 14476 22092 14756 22094
rect 14812 22204 14924 22260
rect 14812 22146 14868 22204
rect 14924 22194 14980 22204
rect 15036 22258 15092 22270
rect 15036 22206 15038 22258
rect 15090 22206 15092 22258
rect 14812 22094 14814 22146
rect 14866 22094 14868 22146
rect 14476 22082 14532 22092
rect 14812 22082 14868 22094
rect 15036 21924 15092 22206
rect 15036 21858 15092 21868
rect 15596 22260 15652 22270
rect 12908 21810 13188 21812
rect 12908 21758 13134 21810
rect 13186 21758 13188 21810
rect 12908 21756 13188 21758
rect 4284 21588 4340 21598
rect 4284 21494 4340 21532
rect 9996 21588 10052 21598
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 9996 20914 10052 21532
rect 9996 20862 9998 20914
rect 10050 20862 10052 20914
rect 4284 20804 4340 20814
rect 4284 20710 4340 20748
rect 9996 20692 10052 20862
rect 12572 20804 12628 20814
rect 9996 20626 10052 20636
rect 12124 20690 12180 20702
rect 12124 20638 12126 20690
rect 12178 20638 12180 20690
rect 4172 20514 4228 20524
rect 2044 20178 2100 20188
rect 4284 20020 4340 20030
rect 4284 19926 4340 19964
rect 10108 20020 10164 20030
rect 10108 19906 10164 19964
rect 10108 19854 10110 19906
rect 10162 19854 10164 19906
rect 10108 19842 10164 19854
rect 12124 19908 12180 20638
rect 12236 20356 12292 20366
rect 12236 20130 12292 20300
rect 12236 20078 12238 20130
rect 12290 20078 12292 20130
rect 12236 20066 12292 20078
rect 12124 19842 12180 19852
rect 1932 19796 1988 19806
rect 1932 19702 1988 19740
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 12124 19348 12180 19358
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 12124 16882 12180 19292
rect 12572 19122 12628 20748
rect 12908 20802 12964 21756
rect 13132 21746 13188 21756
rect 13804 21476 13860 21486
rect 13804 21026 13860 21420
rect 13804 20974 13806 21026
rect 13858 20974 13860 21026
rect 13804 20962 13860 20974
rect 15036 21028 15092 21038
rect 14252 20860 14756 20916
rect 12908 20750 12910 20802
rect 12962 20750 12964 20802
rect 12796 20020 12852 20030
rect 12796 19236 12852 19964
rect 12908 20018 12964 20750
rect 12908 19966 12910 20018
rect 12962 19966 12964 20018
rect 12908 19348 12964 19966
rect 13468 20802 13524 20814
rect 13468 20750 13470 20802
rect 13522 20750 13524 20802
rect 13468 20130 13524 20750
rect 13916 20802 13972 20814
rect 13916 20750 13918 20802
rect 13970 20750 13972 20802
rect 13804 20578 13860 20590
rect 13804 20526 13806 20578
rect 13858 20526 13860 20578
rect 13804 20356 13860 20526
rect 13804 20290 13860 20300
rect 13916 20188 13972 20750
rect 14252 20802 14308 20860
rect 14252 20750 14254 20802
rect 14306 20750 14308 20802
rect 14252 20738 14308 20750
rect 13468 20078 13470 20130
rect 13522 20078 13524 20130
rect 13356 19908 13412 19918
rect 13356 19814 13412 19852
rect 13468 19796 13524 20078
rect 13468 19730 13524 19740
rect 13580 20132 13972 20188
rect 14476 20242 14532 20860
rect 14700 20804 14756 20860
rect 14812 20804 14868 20814
rect 14700 20802 14868 20804
rect 14700 20750 14814 20802
rect 14866 20750 14868 20802
rect 14700 20748 14868 20750
rect 14812 20738 14868 20748
rect 15036 20802 15092 20972
rect 15036 20750 15038 20802
rect 15090 20750 15092 20802
rect 15036 20738 15092 20750
rect 15260 20802 15316 20814
rect 15260 20750 15262 20802
rect 15314 20750 15316 20802
rect 14588 20692 14644 20702
rect 14588 20598 14644 20636
rect 14476 20190 14478 20242
rect 14530 20190 14532 20242
rect 14476 20178 14532 20190
rect 14924 20578 14980 20590
rect 14924 20526 14926 20578
rect 14978 20526 14980 20578
rect 14924 20188 14980 20526
rect 14364 20132 14420 20142
rect 13580 19458 13636 20132
rect 14364 20038 14420 20076
rect 14588 20132 14644 20142
rect 14588 20038 14644 20076
rect 14700 20132 14980 20188
rect 13692 19908 13748 19918
rect 14700 19908 14756 20132
rect 15260 20020 15316 20750
rect 15596 20242 15652 22204
rect 15820 21700 15876 23100
rect 15932 22484 15988 23660
rect 16044 23650 16100 23660
rect 16268 23604 16324 24556
rect 16716 23714 16772 23726
rect 16716 23662 16718 23714
rect 16770 23662 16772 23714
rect 16492 23604 16548 23614
rect 16716 23604 16772 23662
rect 16268 23548 16492 23604
rect 16548 23548 16772 23604
rect 16940 23716 16996 23726
rect 16492 23154 16548 23548
rect 16492 23102 16494 23154
rect 16546 23102 16548 23154
rect 16492 23090 16548 23102
rect 16828 22484 16884 22494
rect 15932 22428 16212 22484
rect 16044 22258 16100 22270
rect 16044 22206 16046 22258
rect 16098 22206 16100 22258
rect 15932 21700 15988 21710
rect 15820 21698 15988 21700
rect 15820 21646 15934 21698
rect 15986 21646 15988 21698
rect 15820 21644 15988 21646
rect 15932 21634 15988 21644
rect 16044 20916 16100 22206
rect 16156 21700 16212 22428
rect 16828 22390 16884 22428
rect 16492 22372 16548 22382
rect 16380 22370 16548 22372
rect 16380 22318 16494 22370
rect 16546 22318 16548 22370
rect 16380 22316 16548 22318
rect 16156 21634 16212 21644
rect 16268 22260 16324 22270
rect 16268 21924 16324 22204
rect 16268 21586 16324 21868
rect 16380 21810 16436 22316
rect 16492 22306 16548 22316
rect 16380 21758 16382 21810
rect 16434 21758 16436 21810
rect 16380 21746 16436 21758
rect 16268 21534 16270 21586
rect 16322 21534 16324 21586
rect 16268 21522 16324 21534
rect 16604 21586 16660 21598
rect 16604 21534 16606 21586
rect 16658 21534 16660 21586
rect 16044 20850 16100 20860
rect 16492 21476 16548 21486
rect 15596 20190 15598 20242
rect 15650 20190 15652 20242
rect 15596 20132 15652 20190
rect 15596 20066 15652 20076
rect 15260 19954 15316 19964
rect 15820 20018 15876 20030
rect 15820 19966 15822 20018
rect 15874 19966 15876 20018
rect 13692 19906 14756 19908
rect 13692 19854 13694 19906
rect 13746 19854 14756 19906
rect 13692 19852 14756 19854
rect 13692 19842 13748 19852
rect 13580 19406 13582 19458
rect 13634 19406 13636 19458
rect 13580 19394 13636 19406
rect 12908 19282 12964 19292
rect 13356 19348 13412 19358
rect 12796 19142 12852 19180
rect 12572 19070 12574 19122
rect 12626 19070 12628 19122
rect 12572 19058 12628 19070
rect 12796 16996 12852 17006
rect 12796 16902 12852 16940
rect 12124 16830 12126 16882
rect 12178 16830 12180 16882
rect 12124 16818 12180 16830
rect 13356 16772 13412 19292
rect 14028 19348 14084 19358
rect 14028 19254 14084 19292
rect 15036 19348 15092 19358
rect 15820 19348 15876 19966
rect 13468 19236 13524 19246
rect 13468 19142 13524 19180
rect 14476 18452 14532 18462
rect 15036 18452 15092 19292
rect 15484 19292 15876 19348
rect 16492 19346 16548 21420
rect 16604 20804 16660 21534
rect 16604 20738 16660 20748
rect 16940 21028 16996 23660
rect 17164 22372 17220 25342
rect 17948 25284 18004 25294
rect 17836 25228 17948 25284
rect 17836 24724 17892 25228
rect 17948 25218 18004 25228
rect 17948 24948 18004 24958
rect 18172 24948 18228 26236
rect 18396 26226 18452 26236
rect 18732 25618 18788 27020
rect 18844 27010 18900 27020
rect 18844 26516 18900 26526
rect 18844 26402 18900 26460
rect 19516 26514 19572 27132
rect 19628 27122 19684 27132
rect 20300 27746 20356 31892
rect 23436 28756 23492 28766
rect 21420 28642 21476 28654
rect 21420 28590 21422 28642
rect 21474 28590 21476 28642
rect 20300 27694 20302 27746
rect 20354 27694 20356 27746
rect 19852 27074 19908 27086
rect 19852 27022 19854 27074
rect 19906 27022 19908 27074
rect 19852 26908 19908 27022
rect 20188 27076 20244 27086
rect 20188 26982 20244 27020
rect 19516 26462 19518 26514
rect 19570 26462 19572 26514
rect 19516 26450 19572 26462
rect 19628 26852 19908 26908
rect 20076 26964 20132 26974
rect 20300 26908 20356 27694
rect 20636 27748 20692 27758
rect 20860 27748 20916 27758
rect 20692 27746 20916 27748
rect 20692 27694 20862 27746
rect 20914 27694 20916 27746
rect 20692 27692 20916 27694
rect 20076 26870 20132 26908
rect 20188 26852 20356 26908
rect 20524 26962 20580 26974
rect 20524 26910 20526 26962
rect 20578 26910 20580 26962
rect 19628 26516 19684 26852
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19740 26516 19796 26526
rect 19628 26514 19796 26516
rect 19628 26462 19742 26514
rect 19794 26462 19796 26514
rect 19628 26460 19796 26462
rect 19740 26450 19796 26460
rect 19852 26516 19908 26526
rect 19852 26422 19908 26460
rect 20076 26516 20132 26526
rect 20188 26516 20244 26852
rect 20076 26514 20244 26516
rect 20076 26462 20078 26514
rect 20130 26462 20244 26514
rect 20076 26460 20244 26462
rect 20076 26450 20132 26460
rect 18844 26350 18846 26402
rect 18898 26350 18900 26402
rect 18844 26338 18900 26350
rect 19180 26404 19236 26414
rect 19068 26292 19124 26302
rect 19180 26292 19236 26348
rect 20524 26404 20580 26910
rect 20524 26338 20580 26348
rect 19068 26290 19236 26292
rect 19068 26238 19070 26290
rect 19122 26238 19236 26290
rect 19068 26236 19236 26238
rect 19068 26226 19124 26236
rect 18732 25566 18734 25618
rect 18786 25566 18788 25618
rect 18732 25554 18788 25566
rect 19068 25506 19124 25518
rect 19068 25454 19070 25506
rect 19122 25454 19124 25506
rect 18508 25284 18564 25294
rect 18508 25190 18564 25228
rect 18732 25282 18788 25294
rect 18732 25230 18734 25282
rect 18786 25230 18788 25282
rect 18732 25060 18788 25230
rect 17948 24946 18228 24948
rect 17948 24894 17950 24946
rect 18002 24894 18228 24946
rect 17948 24892 18228 24894
rect 18396 25004 18788 25060
rect 17948 24882 18004 24892
rect 17948 24724 18004 24734
rect 17612 24722 18004 24724
rect 17612 24670 17950 24722
rect 18002 24670 18004 24722
rect 17612 24668 18004 24670
rect 17388 23828 17444 23838
rect 17164 22306 17220 22316
rect 17276 23826 17444 23828
rect 17276 23774 17390 23826
rect 17442 23774 17444 23826
rect 17276 23772 17444 23774
rect 17276 21924 17332 23772
rect 17388 23762 17444 23772
rect 17500 23716 17556 23726
rect 17500 23622 17556 23660
rect 17612 23492 17668 24668
rect 17948 24658 18004 24668
rect 18172 24722 18228 24734
rect 18172 24670 18174 24722
rect 18226 24670 18228 24722
rect 18172 24276 18228 24670
rect 17724 24220 18228 24276
rect 18396 24722 18452 25004
rect 18396 24670 18398 24722
rect 18450 24670 18452 24722
rect 17724 23938 17780 24220
rect 18284 24164 18340 24174
rect 17724 23886 17726 23938
rect 17778 23886 17780 23938
rect 17724 23874 17780 23886
rect 17836 24108 18284 24164
rect 17388 23436 17668 23492
rect 17388 23378 17444 23436
rect 17836 23380 17892 24108
rect 18284 24098 18340 24108
rect 18396 23828 18452 24670
rect 18620 24724 18676 24734
rect 18620 24630 18676 24668
rect 19068 24724 19124 25454
rect 19068 24658 19124 24668
rect 18396 23772 18676 23828
rect 17388 23326 17390 23378
rect 17442 23326 17444 23378
rect 17388 23314 17444 23326
rect 17500 23324 17892 23380
rect 18508 23604 18564 23614
rect 17276 21858 17332 21868
rect 17500 22258 17556 23324
rect 17724 23154 17780 23166
rect 17724 23102 17726 23154
rect 17778 23102 17780 23154
rect 17612 22372 17668 22382
rect 17612 22278 17668 22316
rect 17500 22206 17502 22258
rect 17554 22206 17556 22258
rect 17500 21476 17556 22206
rect 17500 21410 17556 21420
rect 16940 20690 16996 20972
rect 16940 20638 16942 20690
rect 16994 20638 16996 20690
rect 16940 20626 16996 20638
rect 17276 20692 17332 20702
rect 17276 20598 17332 20636
rect 16716 20132 16772 20142
rect 17612 20132 17668 20142
rect 16716 20038 16772 20076
rect 17500 20130 17668 20132
rect 17500 20078 17614 20130
rect 17666 20078 17668 20130
rect 17500 20076 17668 20078
rect 16604 20018 16660 20030
rect 16604 19966 16606 20018
rect 16658 19966 16660 20018
rect 16604 19684 16660 19966
rect 16604 19618 16660 19628
rect 16940 20018 16996 20030
rect 16940 19966 16942 20018
rect 16994 19966 16996 20018
rect 16492 19294 16494 19346
rect 16546 19294 16548 19346
rect 15372 18564 15428 18574
rect 15484 18564 15540 19292
rect 16492 19282 16548 19294
rect 16156 19236 16212 19246
rect 15596 19234 16212 19236
rect 15596 19182 16158 19234
rect 16210 19182 16212 19234
rect 15596 19180 16212 19182
rect 15596 18674 15652 19180
rect 16156 19170 16212 19180
rect 16716 19124 16772 19134
rect 16716 19030 16772 19068
rect 16940 19012 16996 19966
rect 17388 20018 17444 20030
rect 17388 19966 17390 20018
rect 17442 19966 17444 20018
rect 17388 19908 17444 19966
rect 17276 19796 17332 19806
rect 17276 19346 17332 19740
rect 17276 19294 17278 19346
rect 17330 19294 17332 19346
rect 17276 19282 17332 19294
rect 17388 19234 17444 19852
rect 17388 19182 17390 19234
rect 17442 19182 17444 19234
rect 17164 19012 17220 19022
rect 16940 19010 17220 19012
rect 16940 18958 17166 19010
rect 17218 18958 17220 19010
rect 16940 18956 17220 18958
rect 15596 18622 15598 18674
rect 15650 18622 15652 18674
rect 15596 18610 15652 18622
rect 15372 18562 15540 18564
rect 15372 18510 15374 18562
rect 15426 18510 15540 18562
rect 15372 18508 15540 18510
rect 15260 18452 15316 18462
rect 15036 18396 15204 18452
rect 14252 17444 14308 17454
rect 13356 16716 13524 16772
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 13468 16098 13524 16716
rect 14252 16210 14308 17388
rect 14476 17442 14532 18396
rect 15148 17780 15204 18396
rect 15260 18358 15316 18396
rect 15372 17892 15428 18508
rect 16156 18452 16212 18462
rect 16156 18358 16212 18396
rect 16940 18452 16996 18462
rect 16044 18340 16100 18350
rect 15932 18284 16044 18340
rect 15596 17892 15652 17902
rect 15372 17836 15596 17892
rect 15596 17826 15652 17836
rect 15260 17780 15316 17790
rect 15148 17778 15540 17780
rect 15148 17726 15262 17778
rect 15314 17726 15540 17778
rect 15148 17724 15540 17726
rect 15260 17714 15316 17724
rect 14812 17556 14868 17566
rect 14812 17462 14868 17500
rect 15260 17556 15316 17566
rect 14476 17390 14478 17442
rect 14530 17390 14532 17442
rect 14476 16996 14532 17390
rect 14476 16930 14532 16940
rect 15260 16994 15316 17500
rect 15260 16942 15262 16994
rect 15314 16942 15316 16994
rect 15260 16930 15316 16942
rect 15372 16882 15428 16894
rect 15372 16830 15374 16882
rect 15426 16830 15428 16882
rect 14924 16772 14980 16782
rect 14924 16678 14980 16716
rect 15372 16772 15428 16830
rect 15372 16706 15428 16716
rect 14252 16158 14254 16210
rect 14306 16158 14308 16210
rect 14252 16146 14308 16158
rect 15484 16212 15540 17724
rect 15708 17444 15764 17454
rect 15596 17442 15764 17444
rect 15596 17390 15710 17442
rect 15762 17390 15764 17442
rect 15596 17388 15764 17390
rect 15596 16772 15652 17388
rect 15708 17378 15764 17388
rect 15932 16884 15988 18284
rect 16044 18246 16100 18284
rect 16044 17780 16100 17790
rect 16044 17554 16100 17724
rect 16940 17666 16996 18396
rect 16940 17614 16942 17666
rect 16994 17614 16996 17666
rect 16940 17602 16996 17614
rect 17164 17668 17220 18956
rect 17388 18564 17444 19182
rect 17276 18508 17444 18564
rect 17276 17780 17332 18508
rect 17500 18452 17556 20076
rect 17612 20066 17668 20076
rect 17724 19794 17780 23102
rect 18172 22148 18228 22158
rect 18172 20914 18228 22092
rect 18508 21698 18564 23548
rect 18620 22484 18676 23772
rect 18732 22484 18788 22494
rect 18620 22428 18732 22484
rect 18732 22418 18788 22428
rect 18732 22148 18788 22158
rect 19180 22148 19236 26236
rect 19404 26292 19460 26302
rect 19404 26198 19460 26236
rect 20188 26292 20244 26302
rect 20188 26198 20244 26236
rect 20636 26178 20692 27692
rect 20860 27682 20916 27692
rect 21420 27188 21476 28590
rect 22092 28530 22148 28542
rect 22092 28478 22094 28530
rect 22146 28478 22148 28530
rect 22092 28082 22148 28478
rect 22092 28030 22094 28082
rect 22146 28030 22148 28082
rect 22092 28018 22148 28030
rect 21420 27122 21476 27132
rect 21980 27970 22036 27982
rect 21980 27918 21982 27970
rect 22034 27918 22036 27970
rect 20636 26126 20638 26178
rect 20690 26126 20692 26178
rect 20524 25284 20580 25294
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19852 24836 19908 24846
rect 19852 24722 19908 24780
rect 19852 24670 19854 24722
rect 19906 24670 19908 24722
rect 19516 24612 19572 24622
rect 19852 24612 19908 24670
rect 19516 24610 19908 24612
rect 19516 24558 19518 24610
rect 19570 24558 19908 24610
rect 19516 24556 19908 24558
rect 20524 24612 20580 25228
rect 20636 24836 20692 26126
rect 21308 26404 21364 26414
rect 21308 25506 21364 26348
rect 21308 25454 21310 25506
rect 21362 25454 21364 25506
rect 21308 25442 21364 25454
rect 21532 25506 21588 25518
rect 21532 25454 21534 25506
rect 21586 25454 21588 25506
rect 21420 25284 21476 25294
rect 21420 25190 21476 25228
rect 21532 24948 21588 25454
rect 21532 24882 21588 24892
rect 21756 25508 21812 25518
rect 20636 24770 20692 24780
rect 20636 24612 20692 24622
rect 20524 24610 20692 24612
rect 20524 24558 20638 24610
rect 20690 24558 20692 24610
rect 20524 24556 20692 24558
rect 19516 23604 19572 24556
rect 20636 24546 20692 24556
rect 21644 23716 21700 23726
rect 19516 23538 19572 23548
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 21644 23378 21700 23660
rect 21644 23326 21646 23378
rect 21698 23326 21700 23378
rect 21644 23314 21700 23326
rect 20972 23268 21028 23278
rect 20972 23174 21028 23212
rect 20860 23156 20916 23166
rect 20860 23062 20916 23100
rect 21196 23156 21252 23166
rect 21196 23062 21252 23100
rect 21420 23154 21476 23166
rect 21756 23156 21812 25452
rect 21980 24724 22036 27918
rect 22204 27860 22260 27870
rect 23212 27860 23268 27870
rect 22204 27858 23268 27860
rect 22204 27806 22206 27858
rect 22258 27806 23214 27858
rect 23266 27806 23268 27858
rect 22204 27804 23268 27806
rect 22204 27794 22260 27804
rect 23212 27794 23268 27804
rect 23436 27858 23492 28700
rect 23436 27806 23438 27858
rect 23490 27806 23492 27858
rect 23436 27794 23492 27806
rect 23100 27634 23156 27646
rect 23100 27582 23102 27634
rect 23154 27582 23156 27634
rect 22876 27188 22932 27198
rect 22876 27074 22932 27132
rect 22876 27022 22878 27074
rect 22930 27022 22932 27074
rect 22876 27010 22932 27022
rect 23100 26964 23156 27582
rect 23436 26964 23492 26974
rect 23100 26908 23436 26964
rect 23324 26290 23380 26302
rect 23324 26238 23326 26290
rect 23378 26238 23380 26290
rect 21420 23102 21422 23154
rect 21474 23102 21476 23154
rect 20300 23044 20356 23054
rect 19292 22372 19348 22382
rect 19516 22372 19572 22382
rect 19292 22370 19460 22372
rect 19292 22318 19294 22370
rect 19346 22318 19460 22370
rect 19292 22316 19460 22318
rect 19292 22306 19348 22316
rect 19404 22148 19460 22316
rect 19516 22278 19572 22316
rect 19852 22260 19908 22270
rect 19628 22258 19908 22260
rect 19628 22206 19854 22258
rect 19906 22206 19908 22258
rect 19628 22204 19908 22206
rect 19516 22148 19572 22158
rect 19180 22092 19348 22148
rect 19404 22092 19516 22148
rect 18732 22054 18788 22092
rect 18508 21646 18510 21698
rect 18562 21646 18564 21698
rect 18508 21634 18564 21646
rect 18172 20862 18174 20914
rect 18226 20862 18228 20914
rect 17948 20802 18004 20814
rect 17948 20750 17950 20802
rect 18002 20750 18004 20802
rect 17948 20692 18004 20750
rect 17948 20468 18004 20636
rect 17724 19742 17726 19794
rect 17778 19742 17780 19794
rect 17612 19348 17668 19358
rect 17612 19122 17668 19292
rect 17612 19070 17614 19122
rect 17666 19070 17668 19122
rect 17612 19058 17668 19070
rect 17724 19124 17780 19742
rect 17724 19058 17780 19068
rect 17836 20412 18004 20468
rect 17500 18386 17556 18396
rect 17388 18338 17444 18350
rect 17388 18286 17390 18338
rect 17442 18286 17444 18338
rect 17388 18228 17444 18286
rect 17836 18228 17892 20412
rect 17948 20018 18004 20030
rect 17948 19966 17950 20018
rect 18002 19966 18004 20018
rect 17948 19684 18004 19966
rect 17948 19618 18004 19628
rect 18172 19460 18228 20862
rect 18844 20916 18900 20926
rect 18844 20822 18900 20860
rect 18284 20804 18340 20814
rect 18284 20578 18340 20748
rect 18732 20804 18788 20814
rect 18732 20710 18788 20748
rect 18284 20526 18286 20578
rect 18338 20526 18340 20578
rect 18284 20514 18340 20526
rect 18956 20578 19012 20590
rect 19180 20580 19236 20590
rect 18956 20526 18958 20578
rect 19010 20526 19012 20578
rect 18620 20132 18676 20142
rect 18956 20132 19012 20526
rect 18620 20018 18676 20076
rect 18620 19966 18622 20018
rect 18674 19966 18676 20018
rect 18620 19684 18676 19966
rect 18620 19618 18676 19628
rect 18844 20076 18956 20132
rect 18172 19404 18340 19460
rect 17388 18172 17892 18228
rect 17948 18450 18004 18462
rect 17948 18398 17950 18450
rect 18002 18398 18004 18450
rect 17948 18340 18004 18398
rect 17388 17780 17444 17790
rect 17276 17778 17444 17780
rect 17276 17726 17390 17778
rect 17442 17726 17444 17778
rect 17276 17724 17444 17726
rect 17388 17714 17444 17724
rect 17724 17780 17780 17790
rect 17724 17686 17780 17724
rect 17164 17602 17220 17612
rect 16044 17502 16046 17554
rect 16098 17502 16100 17554
rect 16044 17490 16100 17502
rect 16716 17444 16772 17454
rect 16716 17350 16772 17388
rect 17948 17106 18004 18284
rect 18284 18450 18340 19404
rect 18844 19348 18900 20076
rect 18956 20066 19012 20076
rect 19068 20578 19236 20580
rect 19068 20526 19182 20578
rect 19234 20526 19236 20578
rect 19068 20524 19236 20526
rect 18844 19254 18900 19292
rect 18956 19908 19012 19918
rect 18620 19234 18676 19246
rect 18620 19182 18622 19234
rect 18674 19182 18676 19234
rect 18284 18398 18286 18450
rect 18338 18398 18340 18450
rect 18284 17780 18340 18398
rect 18284 17714 18340 17724
rect 18508 18564 18564 18574
rect 17948 17054 17950 17106
rect 18002 17054 18004 17106
rect 17948 17042 18004 17054
rect 15932 16882 16436 16884
rect 15932 16830 15934 16882
rect 15986 16830 16436 16882
rect 15932 16828 16436 16830
rect 15932 16818 15988 16828
rect 15596 16706 15652 16716
rect 13468 16046 13470 16098
rect 13522 16046 13524 16098
rect 13468 16034 13524 16046
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 15484 14532 15540 16156
rect 16380 16210 16436 16828
rect 18508 16882 18564 18508
rect 18508 16830 18510 16882
rect 18562 16830 18564 16882
rect 18508 16818 18564 16830
rect 18620 17444 18676 19182
rect 18956 19234 19012 19852
rect 18956 19182 18958 19234
rect 19010 19182 19012 19234
rect 18956 19170 19012 19182
rect 19068 18564 19124 20524
rect 19180 20514 19236 20524
rect 19292 20356 19348 22092
rect 19516 22082 19572 22092
rect 19404 21924 19460 21934
rect 19460 21868 19572 21924
rect 19404 21858 19460 21868
rect 19180 20300 19348 20356
rect 19404 20692 19460 20702
rect 19180 19458 19236 20300
rect 19404 20018 19460 20636
rect 19404 19966 19406 20018
rect 19458 19966 19460 20018
rect 19404 19954 19460 19966
rect 19516 20020 19572 21868
rect 19628 20244 19684 22204
rect 19852 22194 19908 22204
rect 20188 22036 20244 22046
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20188 21812 20244 21980
rect 20076 21756 20244 21812
rect 20300 21924 20356 22988
rect 21420 22932 21476 23102
rect 20524 22876 21476 22932
rect 21644 23100 21812 23156
rect 21868 23268 21924 23278
rect 20076 20802 20132 21756
rect 20300 20914 20356 21868
rect 20300 20862 20302 20914
rect 20354 20862 20356 20914
rect 20300 20850 20356 20862
rect 20412 22258 20468 22270
rect 20412 22206 20414 22258
rect 20466 22206 20468 22258
rect 20412 21588 20468 22206
rect 20076 20750 20078 20802
rect 20130 20750 20132 20802
rect 20076 20738 20132 20750
rect 19740 20692 19796 20702
rect 19740 20598 19796 20636
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20412 20244 20468 21532
rect 19628 20178 19684 20188
rect 20076 20188 20468 20244
rect 19516 19964 19908 20020
rect 19292 19908 19348 19918
rect 19292 19814 19348 19852
rect 19852 19908 19908 19964
rect 19180 19406 19182 19458
rect 19234 19406 19236 19458
rect 19180 19394 19236 19406
rect 19628 19796 19684 19806
rect 19628 19234 19684 19740
rect 19852 19794 19908 19852
rect 19852 19742 19854 19794
rect 19906 19742 19908 19794
rect 19852 19730 19908 19742
rect 19628 19182 19630 19234
rect 19682 19182 19684 19234
rect 19628 19170 19684 19182
rect 19964 19236 20020 19246
rect 20076 19236 20132 20188
rect 20524 20020 20580 22876
rect 21644 22820 21700 23100
rect 21196 22764 21700 22820
rect 21756 22930 21812 22942
rect 21756 22878 21758 22930
rect 21810 22878 21812 22930
rect 20748 22372 20804 22382
rect 20748 22278 20804 22316
rect 20860 20580 20916 20590
rect 20860 20486 20916 20524
rect 20972 20020 21028 20030
rect 20524 20018 20916 20020
rect 20524 19966 20526 20018
rect 20578 19966 20916 20018
rect 20524 19964 20916 19966
rect 20524 19954 20580 19964
rect 20748 19348 20804 19358
rect 20748 19254 20804 19292
rect 19964 19234 20132 19236
rect 19964 19182 19966 19234
rect 20018 19182 20132 19234
rect 19964 19180 20132 19182
rect 20300 19234 20356 19246
rect 20300 19182 20302 19234
rect 20354 19182 20356 19234
rect 19964 19170 20020 19180
rect 19740 19012 19796 19022
rect 18956 18562 19124 18564
rect 18956 18510 19070 18562
rect 19122 18510 19124 18562
rect 18956 18508 19124 18510
rect 19628 19010 19796 19012
rect 19628 18958 19742 19010
rect 19794 18958 19796 19010
rect 19628 18956 19796 18958
rect 19628 18564 19684 18956
rect 19740 18946 19796 18956
rect 20300 19012 20356 19182
rect 20300 18956 20692 19012
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19740 18564 19796 18574
rect 19628 18508 19740 18564
rect 18844 18340 18900 18350
rect 18844 18246 18900 18284
rect 16380 16158 16382 16210
rect 16434 16158 16436 16210
rect 16380 16146 16436 16158
rect 16716 16212 16772 16222
rect 16772 16156 16884 16212
rect 16716 16146 16772 16156
rect 16828 16098 16884 16156
rect 16828 16046 16830 16098
rect 16882 16046 16884 16098
rect 16828 16034 16884 16046
rect 18172 15876 18228 15886
rect 18060 15540 18116 15550
rect 17500 15538 18116 15540
rect 17500 15486 18062 15538
rect 18114 15486 18116 15538
rect 17500 15484 18116 15486
rect 17500 15426 17556 15484
rect 18060 15474 18116 15484
rect 18172 15538 18228 15820
rect 18172 15486 18174 15538
rect 18226 15486 18228 15538
rect 18172 15474 18228 15486
rect 17500 15374 17502 15426
rect 17554 15374 17556 15426
rect 17500 15362 17556 15374
rect 17948 15314 18004 15326
rect 17948 15262 17950 15314
rect 18002 15262 18004 15314
rect 16156 15204 16212 15214
rect 16156 14642 16212 15148
rect 17388 15204 17444 15242
rect 17388 15138 17444 15148
rect 16156 14590 16158 14642
rect 16210 14590 16212 14642
rect 16156 14578 16212 14590
rect 17948 14644 18004 15262
rect 18396 15316 18452 15326
rect 18396 15222 18452 15260
rect 18620 15314 18676 17388
rect 18620 15262 18622 15314
rect 18674 15262 18676 15314
rect 18620 15250 18676 15262
rect 18844 16100 18900 16110
rect 18844 15314 18900 16044
rect 18956 15652 19012 18508
rect 19068 18498 19124 18508
rect 19740 18470 19796 18508
rect 20188 18562 20244 18574
rect 20188 18510 20190 18562
rect 20242 18510 20244 18562
rect 19292 18450 19348 18462
rect 19292 18398 19294 18450
rect 19346 18398 19348 18450
rect 19292 17892 19348 18398
rect 19292 17826 19348 17836
rect 20188 18340 20244 18510
rect 20188 17780 20244 18284
rect 20188 17686 20244 17724
rect 19068 17668 19124 17678
rect 19068 17574 19124 17612
rect 19852 17666 19908 17678
rect 19852 17614 19854 17666
rect 19906 17614 19908 17666
rect 19180 17442 19236 17454
rect 19180 17390 19182 17442
rect 19234 17390 19236 17442
rect 19180 17108 19236 17390
rect 19404 17444 19460 17454
rect 19852 17444 19908 17614
rect 19404 17442 19684 17444
rect 19404 17390 19406 17442
rect 19458 17390 19684 17442
rect 19404 17388 19684 17390
rect 19404 17378 19460 17388
rect 19180 17042 19236 17052
rect 19516 15988 19572 15998
rect 19180 15876 19236 15886
rect 19180 15782 19236 15820
rect 19404 15874 19460 15886
rect 19404 15822 19406 15874
rect 19458 15822 19460 15874
rect 18956 15596 19236 15652
rect 18844 15262 18846 15314
rect 18898 15262 18900 15314
rect 18844 15250 18900 15262
rect 19068 15314 19124 15326
rect 19068 15262 19070 15314
rect 19122 15262 19124 15314
rect 19068 15148 19124 15262
rect 18956 15092 19124 15148
rect 18284 14644 18340 14654
rect 17948 14642 18340 14644
rect 17948 14590 18286 14642
rect 18338 14590 18340 14642
rect 17948 14588 18340 14590
rect 15484 14438 15540 14476
rect 16268 14532 16324 14542
rect 16268 13972 16324 14476
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 16268 12962 16324 13916
rect 17052 14308 17108 14318
rect 17052 13074 17108 14252
rect 17052 13022 17054 13074
rect 17106 13022 17108 13074
rect 17052 13010 17108 13022
rect 16268 12910 16270 12962
rect 16322 12910 16324 12962
rect 16268 12898 16324 12910
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 18284 8428 18340 14588
rect 18844 14532 18900 14542
rect 18956 14532 19012 15092
rect 18844 14530 19012 14532
rect 18844 14478 18846 14530
rect 18898 14478 19012 14530
rect 18844 14476 19012 14478
rect 19180 14530 19236 15596
rect 19404 15540 19460 15822
rect 19404 15474 19460 15484
rect 19180 14478 19182 14530
rect 19234 14478 19236 14530
rect 18844 14466 18900 14476
rect 18956 14308 19012 14318
rect 18956 14214 19012 14252
rect 19180 14308 19236 14478
rect 19180 14242 19236 14252
rect 19292 15426 19348 15438
rect 19292 15374 19294 15426
rect 19346 15374 19348 15426
rect 18508 13972 18564 13982
rect 18508 13878 18564 13916
rect 18956 13972 19012 13982
rect 18956 13746 19012 13916
rect 18956 13694 18958 13746
rect 19010 13694 19012 13746
rect 18956 13682 19012 13694
rect 19180 13076 19236 13086
rect 19292 13076 19348 15374
rect 19404 15314 19460 15326
rect 19404 15262 19406 15314
rect 19458 15262 19460 15314
rect 19404 15204 19460 15262
rect 19516 15316 19572 15932
rect 19516 15250 19572 15260
rect 19404 15138 19460 15148
rect 19628 14756 19684 17388
rect 19852 17378 19908 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20076 17108 20132 17118
rect 20076 17014 20132 17052
rect 20300 17106 20356 18956
rect 20412 18788 20468 18798
rect 20412 17778 20468 18732
rect 20636 18674 20692 18956
rect 20636 18622 20638 18674
rect 20690 18622 20692 18674
rect 20636 18610 20692 18622
rect 20748 18340 20804 18350
rect 20748 18246 20804 18284
rect 20412 17726 20414 17778
rect 20466 17726 20468 17778
rect 20412 17714 20468 17726
rect 20300 17054 20302 17106
rect 20354 17054 20356 17106
rect 20300 17042 20356 17054
rect 20412 17444 20468 17454
rect 20412 16994 20468 17388
rect 20860 17108 20916 19964
rect 20972 19926 21028 19964
rect 20860 17042 20916 17052
rect 21196 17106 21252 22764
rect 21420 22484 21476 22494
rect 21420 22258 21476 22428
rect 21756 22372 21812 22878
rect 21420 22206 21422 22258
rect 21474 22206 21476 22258
rect 21420 22194 21476 22206
rect 21644 22370 21812 22372
rect 21644 22318 21758 22370
rect 21810 22318 21812 22370
rect 21644 22316 21812 22318
rect 21532 21924 21588 21934
rect 21420 20802 21476 20814
rect 21420 20750 21422 20802
rect 21474 20750 21476 20802
rect 21420 20580 21476 20750
rect 21420 20514 21476 20524
rect 21420 19796 21476 19806
rect 21420 19702 21476 19740
rect 21420 19122 21476 19134
rect 21420 19070 21422 19122
rect 21474 19070 21476 19122
rect 21196 17054 21198 17106
rect 21250 17054 21252 17106
rect 21196 17042 21252 17054
rect 21308 18562 21364 18574
rect 21308 18510 21310 18562
rect 21362 18510 21364 18562
rect 21308 17780 21364 18510
rect 21308 17106 21364 17724
rect 21420 18452 21476 19070
rect 21420 17666 21476 18396
rect 21420 17614 21422 17666
rect 21474 17614 21476 17666
rect 21420 17444 21476 17614
rect 21420 17378 21476 17388
rect 21308 17054 21310 17106
rect 21362 17054 21364 17106
rect 21308 17042 21364 17054
rect 21532 17108 21588 21868
rect 21644 20804 21700 22316
rect 21756 22306 21812 22316
rect 21868 21924 21924 23212
rect 21980 22932 22036 24668
rect 22764 25506 22820 25518
rect 22764 25454 22766 25506
rect 22818 25454 22820 25506
rect 22764 25172 22820 25454
rect 23324 25508 23380 26238
rect 23324 25442 23380 25452
rect 22988 25396 23044 25406
rect 22988 25302 23044 25340
rect 22764 24610 22820 25116
rect 23212 24948 23268 24958
rect 23436 24948 23492 26908
rect 23660 26962 23716 26974
rect 23660 26910 23662 26962
rect 23714 26910 23716 26962
rect 23660 26514 23716 26910
rect 23660 26462 23662 26514
rect 23714 26462 23716 26514
rect 23660 26450 23716 26462
rect 23212 24854 23268 24892
rect 23324 24892 23492 24948
rect 23548 26290 23604 26302
rect 23548 26238 23550 26290
rect 23602 26238 23604 26290
rect 22764 24558 22766 24610
rect 22818 24558 22820 24610
rect 22764 24546 22820 24558
rect 22988 24722 23044 24734
rect 22988 24670 22990 24722
rect 23042 24670 23044 24722
rect 22204 23268 22260 23278
rect 22652 23268 22708 23278
rect 22204 23266 22372 23268
rect 22204 23214 22206 23266
rect 22258 23214 22372 23266
rect 22204 23212 22372 23214
rect 22204 23202 22260 23212
rect 22092 23156 22148 23166
rect 22092 23062 22148 23100
rect 22204 22932 22260 22942
rect 21980 22930 22260 22932
rect 21980 22878 22206 22930
rect 22258 22878 22260 22930
rect 21980 22876 22260 22878
rect 22204 22866 22260 22876
rect 21644 20738 21700 20748
rect 21756 21868 21924 21924
rect 21644 20244 21700 20254
rect 21644 18676 21700 20188
rect 21756 20020 21812 21868
rect 21868 20020 21924 20030
rect 21756 20018 21924 20020
rect 21756 19966 21870 20018
rect 21922 19966 21924 20018
rect 21756 19964 21924 19966
rect 21756 19348 21812 19964
rect 21868 19954 21924 19964
rect 22204 20020 22260 20030
rect 22316 20020 22372 23212
rect 22652 23174 22708 23212
rect 22988 22484 23044 24670
rect 23324 23380 23380 24892
rect 23436 24722 23492 24734
rect 23436 24670 23438 24722
rect 23490 24670 23492 24722
rect 23436 23940 23492 24670
rect 23548 24052 23604 26238
rect 23772 26292 23828 26302
rect 23772 26198 23828 26236
rect 23884 25172 23940 37998
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 24220 36482 24276 36494
rect 24220 36430 24222 36482
rect 24274 36430 24276 36482
rect 24220 28756 24276 36430
rect 24556 31948 24612 37998
rect 26796 37490 26852 38556
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 26796 37438 26798 37490
rect 26850 37438 26852 37490
rect 26796 37426 26852 37438
rect 25788 37266 25844 37278
rect 25788 37214 25790 37266
rect 25842 37214 25844 37266
rect 24780 36708 24836 36718
rect 24780 36614 24836 36652
rect 24220 28662 24276 28700
rect 24444 31892 24612 31948
rect 23996 26292 24052 26302
rect 24332 26292 24388 26302
rect 23996 26290 24388 26292
rect 23996 26238 23998 26290
rect 24050 26238 24334 26290
rect 24386 26238 24388 26290
rect 23996 26236 24388 26238
rect 23996 26226 24052 26236
rect 24332 26226 24388 26236
rect 24108 26068 24164 26078
rect 24108 25618 24164 26012
rect 24108 25566 24110 25618
rect 24162 25566 24164 25618
rect 24108 25554 24164 25566
rect 24444 25396 24500 31892
rect 24668 28642 24724 28654
rect 24668 28590 24670 28642
rect 24722 28590 24724 28642
rect 24668 27188 24724 28590
rect 24668 27122 24724 27132
rect 25676 27188 25732 27198
rect 24556 26516 24612 26526
rect 24556 26422 24612 26460
rect 24444 25330 24500 25340
rect 24556 26292 24612 26302
rect 23660 24836 23716 24846
rect 23884 24836 23940 25116
rect 23660 24834 23940 24836
rect 23660 24782 23662 24834
rect 23714 24782 23940 24834
rect 23660 24780 23940 24782
rect 23660 24770 23716 24780
rect 24108 24164 24164 24174
rect 23660 24052 23716 24062
rect 23548 24050 23716 24052
rect 23548 23998 23662 24050
rect 23714 23998 23716 24050
rect 23548 23996 23716 23998
rect 23660 23986 23716 23996
rect 23436 23874 23492 23884
rect 23772 23940 23828 23950
rect 23772 23846 23828 23884
rect 24108 23938 24164 24108
rect 24108 23886 24110 23938
rect 24162 23886 24164 23938
rect 24108 23874 24164 23886
rect 23548 23828 23604 23838
rect 23548 23492 23604 23772
rect 24556 23604 24612 26236
rect 24668 26290 24724 26302
rect 24668 26238 24670 26290
rect 24722 26238 24724 26290
rect 24668 26180 24724 26238
rect 25676 26290 25732 27132
rect 25788 27186 25844 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 25788 27134 25790 27186
rect 25842 27134 25844 27186
rect 25788 26516 25844 27134
rect 26236 27188 26292 27198
rect 26236 27094 26292 27132
rect 40012 27186 40068 27198
rect 40012 27134 40014 27186
rect 40066 27134 40068 27186
rect 26908 27074 26964 27086
rect 26908 27022 26910 27074
rect 26962 27022 26964 27074
rect 25788 26450 25844 26460
rect 26236 26964 26292 26974
rect 26572 26964 26628 26974
rect 26292 26962 26628 26964
rect 26292 26910 26574 26962
rect 26626 26910 26628 26962
rect 26292 26908 26628 26910
rect 25676 26238 25678 26290
rect 25730 26238 25732 26290
rect 24724 26124 24836 26180
rect 24668 26114 24724 26124
rect 24668 25172 24724 25182
rect 24668 23938 24724 25116
rect 24668 23886 24670 23938
rect 24722 23886 24724 23938
rect 24668 23716 24724 23886
rect 24668 23650 24724 23660
rect 23548 23436 23828 23492
rect 23324 23324 23716 23380
rect 23212 23156 23268 23166
rect 23324 23156 23380 23324
rect 23660 23266 23716 23324
rect 23660 23214 23662 23266
rect 23714 23214 23716 23266
rect 23660 23202 23716 23214
rect 23212 23154 23380 23156
rect 23212 23102 23214 23154
rect 23266 23102 23380 23154
rect 23212 23100 23380 23102
rect 23548 23154 23604 23166
rect 23548 23102 23550 23154
rect 23602 23102 23604 23154
rect 23212 23090 23268 23100
rect 23548 23044 23604 23102
rect 23548 22978 23604 22988
rect 23772 22820 23828 23436
rect 24556 23378 24612 23548
rect 24556 23326 24558 23378
rect 24610 23326 24612 23378
rect 24556 23314 24612 23326
rect 23548 22764 23828 22820
rect 24556 23154 24612 23166
rect 24556 23102 24558 23154
rect 24610 23102 24612 23154
rect 22988 22418 23044 22428
rect 23436 22484 23492 22494
rect 23324 22372 23380 22382
rect 23324 22146 23380 22316
rect 23324 22094 23326 22146
rect 23378 22094 23380 22146
rect 22204 20018 22372 20020
rect 22204 19966 22206 20018
rect 22258 19966 22372 20018
rect 22204 19964 22372 19966
rect 22204 19954 22260 19964
rect 22204 19794 22260 19806
rect 22204 19742 22206 19794
rect 22258 19742 22260 19794
rect 21756 19234 21812 19292
rect 21756 19182 21758 19234
rect 21810 19182 21812 19234
rect 21756 19170 21812 19182
rect 21868 19684 21924 19694
rect 21644 18582 21700 18620
rect 21756 18564 21812 18574
rect 20412 16942 20414 16994
rect 20466 16942 20468 16994
rect 20412 16930 20468 16942
rect 20636 16882 20692 16894
rect 21084 16884 21140 16894
rect 20636 16830 20638 16882
rect 20690 16830 20692 16882
rect 20188 16772 20244 16782
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19852 15540 19908 15550
rect 20188 15540 20244 16716
rect 20636 15988 20692 16830
rect 20636 15922 20692 15932
rect 20860 16882 21140 16884
rect 20860 16830 21086 16882
rect 21138 16830 21140 16882
rect 20860 16828 21140 16830
rect 19852 15538 20244 15540
rect 19852 15486 19854 15538
rect 19906 15486 20190 15538
rect 20242 15486 20244 15538
rect 19852 15484 20244 15486
rect 19852 15204 19908 15484
rect 20188 15474 20244 15484
rect 20524 15540 20580 15550
rect 20860 15540 20916 16828
rect 21084 16818 21140 16828
rect 21196 16884 21252 16894
rect 20524 15538 20860 15540
rect 20524 15486 20526 15538
rect 20578 15486 20860 15538
rect 20524 15484 20860 15486
rect 20524 15474 20580 15484
rect 20860 15446 20916 15484
rect 21196 15428 21252 16828
rect 21532 16436 21588 17052
rect 21644 18340 21700 18350
rect 21644 17668 21700 18284
rect 21644 16884 21700 17612
rect 21644 16818 21700 16828
rect 21756 16772 21812 18508
rect 21868 17106 21924 19628
rect 21980 19012 22036 19022
rect 21980 19010 22148 19012
rect 21980 18958 21982 19010
rect 22034 18958 22148 19010
rect 21980 18956 22148 18958
rect 21980 18946 22036 18956
rect 21980 18676 22036 18686
rect 21980 18116 22036 18620
rect 22092 18564 22148 18956
rect 22092 18450 22148 18508
rect 22092 18398 22094 18450
rect 22146 18398 22148 18450
rect 22092 18386 22148 18398
rect 21980 18060 22148 18116
rect 21980 17892 22036 17902
rect 21980 17442 22036 17836
rect 22092 17556 22148 18060
rect 22092 17490 22148 17500
rect 21980 17390 21982 17442
rect 22034 17390 22036 17442
rect 21980 17378 22036 17390
rect 21868 17054 21870 17106
rect 21922 17054 21924 17106
rect 21868 17042 21924 17054
rect 21980 17220 22036 17230
rect 21756 16716 21924 16772
rect 21644 16660 21700 16670
rect 21644 16566 21700 16604
rect 21532 16380 21812 16436
rect 21532 15988 21588 15998
rect 21532 15894 21588 15932
rect 21644 15540 21700 15550
rect 21644 15446 21700 15484
rect 21196 15334 21252 15372
rect 21756 15426 21812 16380
rect 21868 16098 21924 16716
rect 21980 16770 22036 17164
rect 21980 16718 21982 16770
rect 22034 16718 22036 16770
rect 21980 16706 22036 16718
rect 22204 16660 22260 19742
rect 22316 19124 22372 19964
rect 22428 22036 22484 22046
rect 22428 20018 22484 21980
rect 22652 21586 22708 21598
rect 22652 21534 22654 21586
rect 22706 21534 22708 21586
rect 22652 20692 22708 21534
rect 22988 21588 23044 21598
rect 22988 21494 23044 21532
rect 23324 21586 23380 22094
rect 23324 21534 23326 21586
rect 23378 21534 23380 21586
rect 23324 21522 23380 21534
rect 23436 21588 23492 22428
rect 23548 21812 23604 22764
rect 23996 22370 24052 22382
rect 23996 22318 23998 22370
rect 24050 22318 24052 22370
rect 23884 22258 23940 22270
rect 23884 22206 23886 22258
rect 23938 22206 23940 22258
rect 23548 21718 23604 21756
rect 23660 21924 23716 21934
rect 23660 21810 23716 21868
rect 23660 21758 23662 21810
rect 23714 21758 23716 21810
rect 23660 21746 23716 21758
rect 23772 21588 23828 21598
rect 23436 21532 23604 21588
rect 22652 20626 22708 20636
rect 23436 20244 23492 20254
rect 23548 20244 23604 21532
rect 23772 21494 23828 21532
rect 23436 20242 23604 20244
rect 23436 20190 23438 20242
rect 23490 20190 23604 20242
rect 23436 20188 23604 20190
rect 23436 20178 23492 20188
rect 22428 19966 22430 20018
rect 22482 19966 22484 20018
rect 22428 19794 22484 19966
rect 22428 19742 22430 19794
rect 22482 19742 22484 19794
rect 22428 19730 22484 19742
rect 23548 20018 23604 20030
rect 23548 19966 23550 20018
rect 23602 19966 23604 20018
rect 22876 19684 22932 19694
rect 23548 19684 23604 19966
rect 23884 19908 23940 22206
rect 23996 22036 24052 22318
rect 24556 22148 24612 23102
rect 23996 21980 24388 22036
rect 23996 21812 24052 21822
rect 23996 21700 24052 21756
rect 24108 21700 24164 21710
rect 23996 21698 24164 21700
rect 23996 21646 24110 21698
rect 24162 21646 24164 21698
rect 23996 21644 24164 21646
rect 24108 21634 24164 21644
rect 24332 21588 24388 21980
rect 24444 21588 24500 21598
rect 24332 21586 24500 21588
rect 24332 21534 24446 21586
rect 24498 21534 24500 21586
rect 24332 21532 24500 21534
rect 23996 20020 24052 20030
rect 23996 20018 24164 20020
rect 23996 19966 23998 20018
rect 24050 19966 24164 20018
rect 23996 19964 24164 19966
rect 23996 19954 24052 19964
rect 23884 19842 23940 19852
rect 22932 19628 23044 19684
rect 22876 19618 22932 19628
rect 22316 19068 22932 19124
rect 22540 18452 22596 18462
rect 22540 18358 22596 18396
rect 22428 17668 22484 17678
rect 22428 17574 22484 17612
rect 22652 17108 22708 19068
rect 22876 18674 22932 19068
rect 22876 18622 22878 18674
rect 22930 18622 22932 18674
rect 22876 18610 22932 18622
rect 22988 17778 23044 19628
rect 23548 19618 23604 19628
rect 23772 19572 23828 19582
rect 23772 19346 23828 19516
rect 23772 19294 23774 19346
rect 23826 19294 23828 19346
rect 23772 19282 23828 19294
rect 23548 19236 23604 19246
rect 23324 18452 23380 18462
rect 23324 18358 23380 18396
rect 22988 17726 22990 17778
rect 23042 17726 23044 17778
rect 22988 17714 23044 17726
rect 23324 17108 23380 17118
rect 22652 17106 23380 17108
rect 22652 17054 22654 17106
rect 22706 17054 23326 17106
rect 23378 17054 23380 17106
rect 22652 17052 23380 17054
rect 22652 17042 22708 17052
rect 23324 17042 23380 17052
rect 22204 16594 22260 16604
rect 22316 16994 22372 17006
rect 22316 16942 22318 16994
rect 22370 16942 22372 16994
rect 21868 16046 21870 16098
rect 21922 16046 21924 16098
rect 21868 16034 21924 16046
rect 22204 16100 22260 16110
rect 22204 16006 22260 16044
rect 22316 15988 22372 16942
rect 23548 16772 23604 19180
rect 24108 19012 24164 19964
rect 24332 19012 24388 19022
rect 24108 19010 24388 19012
rect 24108 18958 24334 19010
rect 24386 18958 24388 19010
rect 24108 18956 24388 18958
rect 24220 18676 24276 18686
rect 24108 18620 24220 18676
rect 23884 18450 23940 18462
rect 23884 18398 23886 18450
rect 23938 18398 23940 18450
rect 23884 18340 23940 18398
rect 23884 18274 23940 18284
rect 24108 17220 24164 18620
rect 24220 18610 24276 18620
rect 24332 18452 24388 18956
rect 24444 18564 24500 21532
rect 24556 19572 24612 22092
rect 24556 19506 24612 19516
rect 24668 21588 24724 21598
rect 24668 19124 24724 21532
rect 24780 20132 24836 26124
rect 25676 24836 25732 26238
rect 24892 24164 24948 24174
rect 24892 24070 24948 24108
rect 25116 23940 25172 23950
rect 25172 23884 25284 23940
rect 25116 23846 25172 23884
rect 25228 22258 25284 23884
rect 25452 23828 25508 23838
rect 25452 23734 25508 23772
rect 25340 23716 25396 23726
rect 25340 23622 25396 23660
rect 25228 22206 25230 22258
rect 25282 22206 25284 22258
rect 25228 22194 25284 22206
rect 24892 22146 24948 22158
rect 24892 22094 24894 22146
rect 24946 22094 24948 22146
rect 24892 22036 24948 22094
rect 25564 22148 25620 22158
rect 25564 22054 25620 22092
rect 24892 21970 24948 21980
rect 25676 21586 25732 24780
rect 26124 25506 26180 25518
rect 26124 25454 26126 25506
rect 26178 25454 26180 25506
rect 25900 24612 25956 24622
rect 26124 24612 26180 25454
rect 26236 24722 26292 26908
rect 26572 26898 26628 26908
rect 26908 26964 26964 27022
rect 37660 27076 37716 27086
rect 37660 26982 37716 27020
rect 26908 26898 26964 26908
rect 28476 26964 28532 26974
rect 26684 26850 26740 26862
rect 26684 26798 26686 26850
rect 26738 26798 26740 26850
rect 26348 26180 26404 26190
rect 26348 26178 26516 26180
rect 26348 26126 26350 26178
rect 26402 26126 26516 26178
rect 26348 26124 26516 26126
rect 26348 26114 26404 26124
rect 26348 25506 26404 25518
rect 26348 25454 26350 25506
rect 26402 25454 26404 25506
rect 26348 25172 26404 25454
rect 26460 25282 26516 26124
rect 26572 25508 26628 25518
rect 26684 25508 26740 26798
rect 28476 26178 28532 26908
rect 40012 26964 40068 27134
rect 40012 26898 40068 26908
rect 28476 26126 28478 26178
rect 28530 26126 28532 26178
rect 28476 26114 28532 26126
rect 28924 26178 28980 26190
rect 28924 26126 28926 26178
rect 28978 26126 28980 26178
rect 26572 25506 26740 25508
rect 26572 25454 26574 25506
rect 26626 25454 26740 25506
rect 26572 25452 26740 25454
rect 26572 25442 26628 25452
rect 26460 25230 26462 25282
rect 26514 25230 26516 25282
rect 26460 25218 26516 25230
rect 26348 25106 26404 25116
rect 26236 24670 26238 24722
rect 26290 24670 26292 24722
rect 26236 24658 26292 24670
rect 26348 24946 26404 24958
rect 26348 24894 26350 24946
rect 26402 24894 26404 24946
rect 25900 24610 26180 24612
rect 25900 24558 25902 24610
rect 25954 24558 26180 24610
rect 25900 24556 26180 24558
rect 25900 22146 25956 24556
rect 26348 24052 26404 24894
rect 26796 24836 26852 24846
rect 28924 24836 28980 26126
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 40012 25618 40068 25630
rect 40012 25566 40014 25618
rect 40066 25566 40068 25618
rect 37660 25506 37716 25518
rect 37660 25454 37662 25506
rect 37714 25454 37716 25506
rect 26852 24780 26964 24836
rect 26796 24770 26852 24780
rect 26908 24724 26964 24780
rect 28924 24770 28980 24780
rect 30156 24836 30212 24846
rect 26908 24722 27076 24724
rect 26908 24670 26910 24722
rect 26962 24670 27076 24722
rect 26908 24668 27076 24670
rect 26908 24658 26964 24668
rect 26348 23986 26404 23996
rect 26572 24612 26628 24622
rect 26572 24050 26628 24556
rect 26572 23998 26574 24050
rect 26626 23998 26628 24050
rect 26572 23986 26628 23998
rect 26236 23940 26292 23950
rect 26236 23380 26292 23884
rect 26908 23828 26964 23838
rect 26460 23716 26516 23726
rect 26460 23622 26516 23660
rect 26684 23714 26740 23726
rect 26684 23662 26686 23714
rect 26738 23662 26740 23714
rect 26684 23604 26740 23662
rect 26684 23538 26740 23548
rect 26460 23380 26516 23390
rect 26236 23378 26516 23380
rect 26236 23326 26462 23378
rect 26514 23326 26516 23378
rect 26236 23324 26516 23326
rect 26460 23314 26516 23324
rect 25900 22094 25902 22146
rect 25954 22094 25956 22146
rect 25900 21700 25956 22094
rect 26012 23154 26068 23166
rect 26012 23102 26014 23154
rect 26066 23102 26068 23154
rect 26012 21924 26068 23102
rect 26236 23154 26292 23166
rect 26236 23102 26238 23154
rect 26290 23102 26292 23154
rect 26124 22484 26180 22494
rect 26124 22148 26180 22428
rect 26236 22372 26292 23102
rect 26572 23154 26628 23166
rect 26572 23102 26574 23154
rect 26626 23102 26628 23154
rect 26348 23044 26404 23054
rect 26348 22950 26404 22988
rect 26236 22316 26404 22372
rect 26236 22148 26292 22158
rect 26124 22146 26292 22148
rect 26124 22094 26238 22146
rect 26290 22094 26292 22146
rect 26124 22092 26292 22094
rect 26236 22082 26292 22092
rect 26012 21858 26068 21868
rect 26348 21812 26404 22316
rect 26572 22260 26628 23102
rect 26908 22594 26964 23772
rect 27020 23154 27076 24668
rect 27580 24612 27636 24622
rect 27580 24518 27636 24556
rect 28364 24612 28420 24622
rect 27132 23940 27188 23950
rect 28140 23940 28196 23950
rect 27132 23938 28196 23940
rect 27132 23886 27134 23938
rect 27186 23886 28142 23938
rect 28194 23886 28196 23938
rect 27132 23884 28196 23886
rect 27132 23874 27188 23884
rect 28140 23874 28196 23884
rect 28364 23826 28420 24556
rect 29708 24612 29764 24622
rect 29708 24518 29764 24556
rect 28476 24052 28532 24062
rect 28476 23940 28532 23996
rect 28476 23938 28644 23940
rect 28476 23886 28478 23938
rect 28530 23886 28644 23938
rect 28476 23884 28644 23886
rect 28476 23874 28532 23884
rect 28364 23774 28366 23826
rect 28418 23774 28420 23826
rect 28364 23762 28420 23774
rect 27020 23102 27022 23154
rect 27074 23102 27076 23154
rect 27020 23090 27076 23102
rect 27804 23044 27860 23054
rect 27804 22950 27860 22988
rect 28476 23044 28532 23054
rect 26908 22542 26910 22594
rect 26962 22542 26964 22594
rect 26908 22530 26964 22542
rect 28364 22484 28420 22494
rect 26572 22166 26628 22204
rect 27244 22370 27300 22382
rect 27244 22318 27246 22370
rect 27298 22318 27300 22370
rect 26348 21746 26404 21756
rect 27020 22146 27076 22158
rect 27020 22094 27022 22146
rect 27074 22094 27076 22146
rect 25900 21634 25956 21644
rect 25676 21534 25678 21586
rect 25730 21534 25732 21586
rect 25676 21522 25732 21534
rect 26460 21476 26516 21486
rect 25788 21474 26516 21476
rect 25788 21422 26462 21474
rect 26514 21422 26516 21474
rect 25788 21420 26516 21422
rect 25116 20692 25172 20702
rect 25172 20636 25284 20692
rect 25116 20598 25172 20636
rect 24780 20066 24836 20076
rect 24892 20468 24948 20478
rect 24892 19234 24948 20412
rect 25228 20018 25284 20636
rect 25228 19966 25230 20018
rect 25282 19966 25284 20018
rect 25228 19954 25284 19966
rect 25564 20132 25620 20142
rect 24892 19182 24894 19234
rect 24946 19182 24948 19234
rect 24668 19122 24836 19124
rect 24668 19070 24670 19122
rect 24722 19070 24836 19122
rect 24668 19068 24836 19070
rect 24668 19058 24724 19068
rect 24444 18498 24500 18508
rect 24332 18386 24388 18396
rect 24668 18340 24724 18350
rect 24220 17890 24276 17902
rect 24220 17838 24222 17890
rect 24274 17838 24276 17890
rect 24220 17780 24276 17838
rect 24220 17714 24276 17724
rect 24668 17778 24724 18284
rect 24668 17726 24670 17778
rect 24722 17726 24724 17778
rect 24668 17714 24724 17726
rect 24220 17556 24276 17566
rect 24220 17462 24276 17500
rect 24332 17556 24388 17566
rect 24332 17554 24612 17556
rect 24332 17502 24334 17554
rect 24386 17502 24612 17554
rect 24332 17500 24612 17502
rect 24332 17490 24388 17500
rect 23660 17164 24388 17220
rect 23660 17106 23716 17164
rect 23660 17054 23662 17106
rect 23714 17054 23716 17106
rect 23660 17042 23716 17054
rect 24332 17108 24388 17164
rect 24332 17106 24500 17108
rect 24332 17054 24334 17106
rect 24386 17054 24500 17106
rect 24332 17052 24500 17054
rect 24332 17042 24388 17052
rect 24220 16996 24276 17006
rect 24220 16902 24276 16940
rect 23548 16706 23604 16716
rect 22316 15922 22372 15932
rect 24332 16660 24388 16670
rect 21980 15876 22036 15886
rect 21980 15782 22036 15820
rect 23884 15876 23940 15886
rect 21756 15374 21758 15426
rect 21810 15374 21812 15426
rect 21756 15362 21812 15374
rect 21868 15428 21924 15438
rect 19852 15138 19908 15148
rect 21420 15314 21476 15326
rect 21420 15262 21422 15314
rect 21474 15262 21476 15314
rect 19404 14532 19460 14542
rect 19628 14532 19684 14700
rect 19404 14530 19684 14532
rect 19404 14478 19406 14530
rect 19458 14478 19684 14530
rect 19404 14476 19684 14478
rect 20076 14532 20132 14542
rect 19404 14466 19460 14476
rect 20076 14438 20132 14476
rect 21420 14532 21476 15262
rect 21420 14466 21476 14476
rect 19740 14308 19796 14318
rect 19628 14306 19796 14308
rect 19628 14254 19742 14306
rect 19794 14254 19796 14306
rect 19628 14252 19796 14254
rect 19628 13972 19684 14252
rect 19740 14242 19796 14252
rect 19964 14308 20020 14346
rect 19964 14242 20020 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19852 13972 19908 13982
rect 19628 13916 19796 13972
rect 19740 13858 19796 13916
rect 19740 13806 19742 13858
rect 19794 13806 19796 13858
rect 19740 13794 19796 13806
rect 19852 13636 19908 13916
rect 17612 8372 18340 8428
rect 19068 13074 19348 13076
rect 19068 13022 19182 13074
rect 19234 13022 19348 13074
rect 19068 13020 19348 13022
rect 19740 13076 19796 13086
rect 19852 13076 19908 13580
rect 21868 13634 21924 15372
rect 23884 15316 23940 15820
rect 22204 15092 22260 15102
rect 22204 14756 22260 15036
rect 22204 14662 22260 14700
rect 21980 14532 22036 14542
rect 21980 14438 22036 14476
rect 22540 14532 22596 14542
rect 22540 14438 22596 14476
rect 23436 14532 23492 14542
rect 23436 13746 23492 14476
rect 23884 14530 23940 15260
rect 24332 14532 24388 16604
rect 24444 15148 24500 17052
rect 24556 17106 24612 17500
rect 24556 17054 24558 17106
rect 24610 17054 24612 17106
rect 24556 17042 24612 17054
rect 24780 16100 24836 19068
rect 24892 17220 24948 19182
rect 25452 19908 25508 19918
rect 25340 18564 25396 18574
rect 25340 18470 25396 18508
rect 25452 18562 25508 19852
rect 25564 19236 25620 20076
rect 25564 19142 25620 19180
rect 25788 19234 25844 21420
rect 26460 21410 26516 21420
rect 27020 21140 27076 22094
rect 27244 22148 27300 22318
rect 28028 22372 28084 22382
rect 28028 22370 28308 22372
rect 28028 22318 28030 22370
rect 28082 22318 28308 22370
rect 28028 22316 28308 22318
rect 28028 22306 28084 22316
rect 27244 22082 27300 22092
rect 28140 22148 28196 22158
rect 26572 21084 27076 21140
rect 27132 21700 27188 21710
rect 25788 19182 25790 19234
rect 25842 19182 25844 19234
rect 25788 19170 25844 19182
rect 25900 21028 25956 21038
rect 25900 19234 25956 20972
rect 26572 19458 26628 21084
rect 26908 20692 26964 20702
rect 26908 20598 26964 20636
rect 27132 20690 27188 21644
rect 27132 20638 27134 20690
rect 27186 20638 27188 20690
rect 27020 20580 27076 20590
rect 27020 20486 27076 20524
rect 27132 20188 27188 20638
rect 26572 19406 26574 19458
rect 26626 19406 26628 19458
rect 26572 19394 26628 19406
rect 26684 20132 27188 20188
rect 27916 20804 27972 20814
rect 25900 19182 25902 19234
rect 25954 19182 25956 19234
rect 25900 19170 25956 19182
rect 26460 19234 26516 19246
rect 26460 19182 26462 19234
rect 26514 19182 26516 19234
rect 26236 19124 26292 19134
rect 26236 19030 26292 19068
rect 26460 18788 26516 19182
rect 26460 18722 26516 18732
rect 25452 18510 25454 18562
rect 25506 18510 25508 18562
rect 25452 18498 25508 18510
rect 25788 18452 25844 18462
rect 25788 18358 25844 18396
rect 25900 18340 25956 18350
rect 25900 18246 25956 18284
rect 24892 17154 24948 17164
rect 25340 18226 25396 18238
rect 25340 18174 25342 18226
rect 25394 18174 25396 18226
rect 25340 16660 25396 18174
rect 26684 17556 26740 20132
rect 27020 19236 27076 19246
rect 27020 19142 27076 19180
rect 27692 19124 27748 19134
rect 27692 19030 27748 19068
rect 27916 19122 27972 20748
rect 28028 20580 28084 20590
rect 28028 19234 28084 20524
rect 28140 20356 28196 22092
rect 28252 20468 28308 22316
rect 28364 22370 28420 22428
rect 28476 22482 28532 22988
rect 28476 22430 28478 22482
rect 28530 22430 28532 22482
rect 28476 22418 28532 22430
rect 28364 22318 28366 22370
rect 28418 22318 28420 22370
rect 28364 22306 28420 22318
rect 28588 22370 28644 23884
rect 29260 23380 29316 23390
rect 28588 22318 28590 22370
rect 28642 22318 28644 22370
rect 28588 22306 28644 22318
rect 29036 22932 29092 22942
rect 28812 21812 28868 21822
rect 28812 21718 28868 21756
rect 29036 21810 29092 22876
rect 29260 22372 29316 23324
rect 30156 23380 30212 24780
rect 37660 24612 37716 25454
rect 40012 24948 40068 25566
rect 40012 24882 40068 24892
rect 37660 24546 37716 24556
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 30156 23314 30212 23324
rect 30828 23380 30884 23390
rect 30828 23286 30884 23324
rect 32060 23156 32116 23166
rect 29932 23042 29988 23054
rect 29932 22990 29934 23042
rect 29986 22990 29988 23042
rect 29932 22932 29988 22990
rect 30380 23044 30436 23054
rect 30380 22950 30436 22988
rect 30268 22932 30324 22942
rect 29932 22866 29988 22876
rect 30044 22930 30324 22932
rect 30044 22878 30270 22930
rect 30322 22878 30324 22930
rect 30044 22876 30324 22878
rect 29932 22484 29988 22494
rect 30044 22484 30100 22876
rect 30268 22866 30324 22876
rect 29932 22482 30100 22484
rect 29932 22430 29934 22482
rect 29986 22430 30100 22482
rect 29932 22428 30100 22430
rect 32060 22484 32116 23100
rect 37660 23156 37716 23194
rect 37660 23090 37716 23100
rect 37660 22932 37716 22942
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 29932 22418 29988 22428
rect 32060 22390 32116 22428
rect 29260 22370 29652 22372
rect 29260 22318 29262 22370
rect 29314 22318 29652 22370
rect 29260 22316 29652 22318
rect 29260 22306 29316 22316
rect 29036 21758 29038 21810
rect 29090 21758 29092 21810
rect 29036 21746 29092 21758
rect 29596 21812 29652 22316
rect 37660 22370 37716 22876
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 37660 22318 37662 22370
rect 37714 22318 37716 22370
rect 37660 22306 37716 22318
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 30044 21812 30100 21822
rect 29596 21810 30100 21812
rect 29596 21758 29598 21810
rect 29650 21758 30046 21810
rect 30098 21758 30100 21810
rect 29596 21756 30100 21758
rect 29596 21746 29652 21756
rect 29148 21588 29204 21598
rect 28924 21586 29204 21588
rect 28924 21534 29150 21586
rect 29202 21534 29204 21586
rect 28924 21532 29204 21534
rect 28588 21474 28644 21486
rect 28588 21422 28590 21474
rect 28642 21422 28644 21474
rect 28588 20804 28644 21422
rect 28588 20738 28644 20748
rect 28924 20580 28980 21532
rect 29148 21522 29204 21532
rect 28924 20514 28980 20524
rect 29036 20748 29428 20804
rect 28476 20468 28532 20478
rect 28252 20412 28476 20468
rect 28140 20300 28420 20356
rect 28028 19182 28030 19234
rect 28082 19182 28084 19234
rect 28028 19170 28084 19182
rect 27916 19070 27918 19122
rect 27970 19070 27972 19122
rect 27916 19058 27972 19070
rect 27132 18676 27188 18686
rect 27132 18562 27188 18620
rect 27132 18510 27134 18562
rect 27186 18510 27188 18562
rect 27132 18498 27188 18510
rect 27244 18564 27300 18574
rect 27244 18470 27300 18508
rect 27356 18452 27412 18462
rect 26796 17780 26852 17790
rect 26796 17686 26852 17724
rect 27356 17668 27412 18396
rect 27468 18450 27524 18462
rect 27468 18398 27470 18450
rect 27522 18398 27524 18450
rect 27468 18004 27524 18398
rect 27804 18452 27860 18462
rect 27804 18358 27860 18396
rect 27468 17948 28196 18004
rect 27468 17668 27524 17678
rect 27020 17666 27524 17668
rect 27020 17614 27470 17666
rect 27522 17614 27524 17666
rect 27020 17612 27524 17614
rect 26684 17500 26852 17556
rect 25340 16594 25396 16604
rect 24780 16034 24836 16044
rect 25676 15538 25732 15550
rect 25676 15486 25678 15538
rect 25730 15486 25732 15538
rect 25564 15316 25620 15326
rect 25564 15222 25620 15260
rect 24444 15092 24724 15148
rect 24668 14644 24724 15092
rect 25340 15092 25396 15102
rect 25340 14998 25396 15036
rect 25676 14868 25732 15486
rect 25788 15316 25844 15326
rect 26684 15316 26740 15326
rect 25788 15314 26740 15316
rect 25788 15262 25790 15314
rect 25842 15262 26686 15314
rect 26738 15262 26740 15314
rect 25788 15260 26740 15262
rect 25788 15250 25844 15260
rect 26684 15250 26740 15260
rect 26572 15092 26628 15102
rect 26796 15092 26852 17500
rect 27020 16882 27076 17612
rect 27468 17602 27524 17612
rect 28140 17666 28196 17948
rect 28140 17614 28142 17666
rect 28194 17614 28196 17666
rect 28140 17602 28196 17614
rect 28364 17666 28420 20300
rect 28476 18788 28532 20412
rect 29036 20020 29092 20748
rect 29148 20578 29204 20590
rect 29148 20526 29150 20578
rect 29202 20526 29204 20578
rect 29148 20468 29204 20526
rect 29148 20402 29204 20412
rect 29260 20578 29316 20590
rect 29260 20526 29262 20578
rect 29314 20526 29316 20578
rect 29036 19954 29092 19964
rect 29260 19908 29316 20526
rect 29372 20578 29428 20748
rect 29372 20526 29374 20578
rect 29426 20526 29428 20578
rect 29372 20514 29428 20526
rect 29708 20468 29764 21756
rect 30044 21746 30100 21756
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 30156 21028 30212 21038
rect 29820 21026 30212 21028
rect 29820 20974 30158 21026
rect 30210 20974 30212 21026
rect 29820 20972 30212 20974
rect 29820 20802 29876 20972
rect 30156 20962 30212 20972
rect 40012 20914 40068 20926
rect 40012 20862 40014 20914
rect 40066 20862 40068 20914
rect 29820 20750 29822 20802
rect 29874 20750 29876 20802
rect 29820 20738 29876 20750
rect 37660 20804 37716 20814
rect 37660 20710 37716 20748
rect 30044 20690 30100 20702
rect 30044 20638 30046 20690
rect 30098 20638 30100 20690
rect 30044 20580 30100 20638
rect 30044 20514 30100 20524
rect 30156 20578 30212 20590
rect 30156 20526 30158 20578
rect 30210 20526 30212 20578
rect 29708 20412 29988 20468
rect 29932 20356 29988 20412
rect 29932 20300 30100 20356
rect 30044 20130 30100 20300
rect 30044 20078 30046 20130
rect 30098 20078 30100 20130
rect 29260 19852 29988 19908
rect 29932 19346 29988 19852
rect 29932 19294 29934 19346
rect 29986 19294 29988 19346
rect 29932 19282 29988 19294
rect 28476 18722 28532 18732
rect 28588 19236 28644 19246
rect 29260 19236 29316 19246
rect 28588 19234 29316 19236
rect 28588 19182 28590 19234
rect 28642 19182 29262 19234
rect 29314 19182 29316 19234
rect 28588 19180 29316 19182
rect 28364 17614 28366 17666
rect 28418 17614 28420 17666
rect 28364 17602 28420 17614
rect 28588 18452 28644 19180
rect 29260 19124 29316 19180
rect 30044 19124 30100 20078
rect 30156 20020 30212 20526
rect 40012 20244 40068 20862
rect 40012 20178 40068 20188
rect 30156 19954 30212 19964
rect 32060 20020 32116 20030
rect 32060 19346 32116 19964
rect 37660 20020 37716 20030
rect 37660 19926 37716 19964
rect 40012 19794 40068 19806
rect 40012 19742 40014 19794
rect 40066 19742 40068 19794
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 40012 19572 40068 19742
rect 40012 19506 40068 19516
rect 32060 19294 32062 19346
rect 32114 19294 32116 19346
rect 32060 19282 32116 19294
rect 29260 19068 30212 19124
rect 27916 17556 27972 17566
rect 27916 17462 27972 17500
rect 28028 17442 28084 17454
rect 28028 17390 28030 17442
rect 28082 17390 28084 17442
rect 28028 17108 28084 17390
rect 27692 17052 28084 17108
rect 27692 16994 27748 17052
rect 27692 16942 27694 16994
rect 27746 16942 27748 16994
rect 27692 16930 27748 16942
rect 27020 16830 27022 16882
rect 27074 16830 27076 16882
rect 27020 16818 27076 16830
rect 26908 15316 26964 15326
rect 26908 15222 26964 15260
rect 28252 15316 28308 15326
rect 26572 15090 26852 15092
rect 26572 15038 26574 15090
rect 26626 15038 26852 15090
rect 26572 15036 26852 15038
rect 26572 15026 26628 15036
rect 25676 14812 26180 14868
rect 24556 14642 24724 14644
rect 24556 14590 24670 14642
rect 24722 14590 24724 14642
rect 24556 14588 24724 14590
rect 23884 14478 23886 14530
rect 23938 14478 23940 14530
rect 23884 14466 23940 14478
rect 23996 14530 24388 14532
rect 23996 14478 24334 14530
rect 24386 14478 24388 14530
rect 23996 14476 24388 14478
rect 23996 14308 24052 14476
rect 24332 14466 24388 14476
rect 24444 14532 24500 14542
rect 24444 14438 24500 14476
rect 23436 13694 23438 13746
rect 23490 13694 23492 13746
rect 23436 13682 23492 13694
rect 23660 14252 24052 14308
rect 23660 13746 23716 14252
rect 24108 13858 24164 13870
rect 24108 13806 24110 13858
rect 24162 13806 24164 13858
rect 23660 13694 23662 13746
rect 23714 13694 23716 13746
rect 23660 13682 23716 13694
rect 23996 13748 24052 13758
rect 24108 13748 24164 13806
rect 23996 13746 24164 13748
rect 23996 13694 23998 13746
rect 24050 13694 24164 13746
rect 23996 13692 24164 13694
rect 24332 13858 24388 13870
rect 24332 13806 24334 13858
rect 24386 13806 24388 13858
rect 23996 13682 24052 13692
rect 21868 13582 21870 13634
rect 21922 13582 21924 13634
rect 21868 13570 21924 13582
rect 22316 13636 22372 13646
rect 22316 13542 22372 13580
rect 22988 13636 23044 13646
rect 19740 13074 19908 13076
rect 19740 13022 19742 13074
rect 19794 13022 19908 13074
rect 19740 13020 19908 13022
rect 22988 13074 23044 13580
rect 23772 13636 23828 13646
rect 23772 13542 23828 13580
rect 22988 13022 22990 13074
rect 23042 13022 23044 13074
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 17612 3554 17668 8372
rect 19068 4338 19124 13020
rect 19180 13010 19236 13020
rect 19740 13010 19796 13020
rect 22988 13010 23044 13022
rect 22316 12964 22372 12974
rect 22316 12870 22372 12908
rect 24332 12740 24388 13806
rect 24444 13860 24500 13870
rect 24556 13860 24612 14588
rect 24668 14578 24724 14588
rect 26124 14642 26180 14812
rect 26124 14590 26126 14642
rect 26178 14590 26180 14642
rect 26124 14578 26180 14590
rect 28252 14642 28308 15260
rect 28252 14590 28254 14642
rect 28306 14590 28308 14642
rect 28252 14578 28308 14590
rect 25340 14530 25396 14542
rect 25340 14478 25342 14530
rect 25394 14478 25396 14530
rect 24444 13858 24612 13860
rect 24444 13806 24446 13858
rect 24498 13806 24612 13858
rect 24444 13804 24612 13806
rect 24892 14418 24948 14430
rect 24892 14366 24894 14418
rect 24946 14366 24948 14418
rect 24444 13794 24500 13804
rect 24892 13188 24948 14366
rect 25004 14308 25060 14318
rect 25004 14214 25060 14252
rect 25340 13972 25396 14478
rect 24892 13122 24948 13132
rect 25228 13748 25284 13758
rect 25340 13748 25396 13916
rect 26012 14308 26068 14318
rect 26012 13858 26068 14252
rect 28588 13972 28644 18396
rect 29820 18564 29876 18574
rect 29820 17668 29876 18508
rect 29820 16770 29876 17612
rect 30156 17108 30212 19068
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 37660 17668 37716 17678
rect 37660 17574 37716 17612
rect 30268 17108 30324 17118
rect 30156 17106 30324 17108
rect 30156 17054 30270 17106
rect 30322 17054 30324 17106
rect 30156 17052 30324 17054
rect 30268 17042 30324 17052
rect 40012 16884 40068 17726
rect 40012 16818 40068 16828
rect 29820 16718 29822 16770
rect 29874 16718 29876 16770
rect 29820 16706 29876 16718
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 37660 15316 37716 15326
rect 37660 15222 37716 15260
rect 40012 15202 40068 15214
rect 40012 15150 40014 15202
rect 40066 15150 40068 15202
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 40012 14868 40068 15150
rect 40012 14802 40068 14812
rect 28588 13878 28644 13916
rect 29260 14306 29316 14318
rect 29260 14254 29262 14306
rect 29314 14254 29316 14306
rect 29260 13972 29316 14254
rect 29260 13906 29316 13916
rect 26012 13806 26014 13858
rect 26066 13806 26068 13858
rect 26012 13794 26068 13806
rect 25228 13746 25396 13748
rect 25228 13694 25230 13746
rect 25282 13694 25396 13746
rect 25228 13692 25396 13694
rect 25116 13074 25172 13086
rect 25116 13022 25118 13074
rect 25170 13022 25172 13074
rect 25116 12740 25172 13022
rect 25228 12964 25284 13692
rect 28140 13634 28196 13646
rect 28140 13582 28142 13634
rect 28194 13582 28196 13634
rect 26236 13188 26292 13198
rect 26236 13094 26292 13132
rect 25284 12908 25396 12964
rect 25228 12898 25284 12908
rect 25228 12740 25284 12750
rect 25116 12684 25228 12740
rect 24332 12674 24388 12684
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19068 4286 19070 4338
rect 19122 4286 19124 4338
rect 19068 4274 19124 4286
rect 18844 4116 18900 4126
rect 18620 3668 18676 3678
rect 17612 3502 17614 3554
rect 17666 3502 17668 3554
rect 17612 3490 17668 3502
rect 18172 3666 18676 3668
rect 18172 3614 18622 3666
rect 18674 3614 18676 3666
rect 18172 3612 18676 3614
rect 18172 800 18228 3612
rect 18620 3602 18676 3612
rect 18844 800 18900 4060
rect 20076 4116 20132 4126
rect 20076 4022 20132 4060
rect 25228 3554 25284 12684
rect 25340 12404 25396 12908
rect 26348 12852 26404 12862
rect 26348 12758 26404 12796
rect 28140 12852 28196 13582
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 25452 12740 25508 12750
rect 25452 12646 25508 12684
rect 25788 12738 25844 12750
rect 25788 12686 25790 12738
rect 25842 12686 25844 12738
rect 25452 12404 25508 12414
rect 25340 12402 25508 12404
rect 25340 12350 25454 12402
rect 25506 12350 25508 12402
rect 25340 12348 25508 12350
rect 25452 12338 25508 12348
rect 25788 4338 25844 12686
rect 28140 11844 28196 12796
rect 28140 11788 28644 11844
rect 25788 4286 25790 4338
rect 25842 4286 25844 4338
rect 25788 4274 25844 4286
rect 25228 3502 25230 3554
rect 25282 3502 25284 3554
rect 25228 3490 25284 3502
rect 25564 4116 25620 4126
rect 24892 3444 24948 3454
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 24892 800 24948 3388
rect 25564 800 25620 4060
rect 26796 4116 26852 4126
rect 26796 4022 26852 4060
rect 26124 3666 26180 3678
rect 26124 3614 26126 3666
rect 26178 3614 26180 3666
rect 26124 3444 26180 3614
rect 26124 3378 26180 3388
rect 26236 3668 26292 3678
rect 26236 800 26292 3612
rect 28588 3554 28644 11788
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 29372 3668 29428 3678
rect 29372 3574 29428 3612
rect 28588 3502 28590 3554
rect 28642 3502 28644 3554
rect 28588 3490 28644 3502
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 24864 0 24976 800
rect 25536 0 25648 800
rect 26208 0 26320 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 16828 37436 16884 37492
rect 18396 37490 18452 37492
rect 18396 37438 18398 37490
rect 18398 37438 18450 37490
rect 18450 37438 18452 37490
rect 18396 37436 18452 37438
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4172 28252 4228 28308
rect 1932 24892 1988 24948
rect 1932 23548 1988 23604
rect 1932 22930 1988 22932
rect 1932 22878 1934 22930
rect 1934 22878 1986 22930
rect 1986 22878 1988 22930
rect 1932 22876 1988 22878
rect 1932 20860 1988 20916
rect 16828 27692 16884 27748
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 16380 27186 16436 27188
rect 16380 27134 16382 27186
rect 16382 27134 16434 27186
rect 16434 27134 16436 27186
rect 16380 27132 16436 27134
rect 13580 27074 13636 27076
rect 13580 27022 13582 27074
rect 13582 27022 13634 27074
rect 13634 27022 13636 27074
rect 13580 27020 13636 27022
rect 16604 27020 16660 27076
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 17500 27692 17556 27748
rect 17388 27132 17444 27188
rect 17500 26962 17556 26964
rect 17500 26910 17502 26962
rect 17502 26910 17554 26962
rect 17554 26910 17556 26962
rect 17500 26908 17556 26910
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 22876 38220 22932 38276
rect 20188 37436 20244 37492
rect 21420 37490 21476 37492
rect 21420 37438 21422 37490
rect 21422 37438 21474 37490
rect 21474 37438 21476 37490
rect 21420 37436 21476 37438
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 25564 38556 25620 38612
rect 26796 38556 26852 38612
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 23548 36652 23604 36708
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 18844 27020 18900 27076
rect 18060 26124 18116 26180
rect 14252 25564 14308 25620
rect 16604 26012 16660 26068
rect 4284 25506 4340 25508
rect 4284 25454 4286 25506
rect 4286 25454 4338 25506
rect 4338 25454 4340 25506
rect 4284 25452 4340 25454
rect 12236 25452 12292 25508
rect 17500 26066 17556 26068
rect 17500 26014 17502 26066
rect 17502 26014 17554 26066
rect 17554 26014 17556 26066
rect 17500 26012 17556 26014
rect 16716 25618 16772 25620
rect 16716 25566 16718 25618
rect 16718 25566 16770 25618
rect 16770 25566 16772 25618
rect 16716 25564 16772 25566
rect 16940 25228 16996 25284
rect 15708 25116 15764 25172
rect 14364 24722 14420 24724
rect 14364 24670 14366 24722
rect 14366 24670 14418 24722
rect 14418 24670 14420 24722
rect 14364 24668 14420 24670
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4284 23938 4340 23940
rect 4284 23886 4286 23938
rect 4286 23886 4338 23938
rect 4338 23886 4340 23938
rect 4284 23884 4340 23886
rect 9996 23884 10052 23940
rect 14028 24556 14084 24612
rect 13132 23996 13188 24052
rect 12236 23884 12292 23940
rect 15484 24722 15540 24724
rect 15484 24670 15486 24722
rect 15486 24670 15538 24722
rect 15538 24670 15540 24722
rect 15484 24668 15540 24670
rect 15148 24556 15204 24612
rect 14028 24050 14084 24052
rect 14028 23998 14030 24050
rect 14030 23998 14082 24050
rect 14082 23998 14084 24050
rect 14028 23996 14084 23998
rect 14700 23996 14756 24052
rect 12124 23826 12180 23828
rect 12124 23774 12126 23826
rect 12126 23774 12178 23826
rect 12178 23774 12180 23826
rect 12124 23772 12180 23774
rect 9996 23548 10052 23604
rect 4284 23154 4340 23156
rect 4284 23102 4286 23154
rect 4286 23102 4338 23154
rect 4338 23102 4340 23154
rect 4284 23100 4340 23102
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 13468 23826 13524 23828
rect 13468 23774 13470 23826
rect 13470 23774 13522 23826
rect 13522 23774 13524 23826
rect 13468 23772 13524 23774
rect 13580 23100 13636 23156
rect 14588 23548 14644 23604
rect 15484 23996 15540 24052
rect 16268 24610 16324 24612
rect 16268 24558 16270 24610
rect 16270 24558 16322 24610
rect 16322 24558 16324 24610
rect 16268 24556 16324 24558
rect 15596 23938 15652 23940
rect 15596 23886 15598 23938
rect 15598 23886 15650 23938
rect 15650 23886 15652 23938
rect 15596 23884 15652 23886
rect 15036 23212 15092 23268
rect 15708 23266 15764 23268
rect 15708 23214 15710 23266
rect 15710 23214 15762 23266
rect 15762 23214 15764 23266
rect 15708 23212 15764 23214
rect 14812 22428 14868 22484
rect 15820 23100 15876 23156
rect 14924 22204 14980 22260
rect 15036 21868 15092 21924
rect 15596 22204 15652 22260
rect 4284 21586 4340 21588
rect 4284 21534 4286 21586
rect 4286 21534 4338 21586
rect 4338 21534 4340 21586
rect 4284 21532 4340 21534
rect 9996 21532 10052 21588
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4284 20802 4340 20804
rect 4284 20750 4286 20802
rect 4286 20750 4338 20802
rect 4338 20750 4340 20802
rect 4284 20748 4340 20750
rect 12572 20748 12628 20804
rect 9996 20636 10052 20692
rect 4172 20524 4228 20580
rect 2044 20188 2100 20244
rect 4284 20018 4340 20020
rect 4284 19966 4286 20018
rect 4286 19966 4338 20018
rect 4338 19966 4340 20018
rect 4284 19964 4340 19966
rect 10108 19964 10164 20020
rect 12236 20300 12292 20356
rect 12124 19852 12180 19908
rect 1932 19794 1988 19796
rect 1932 19742 1934 19794
rect 1934 19742 1986 19794
rect 1986 19742 1988 19794
rect 1932 19740 1988 19742
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 12124 19292 12180 19348
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 13804 21420 13860 21476
rect 15036 20972 15092 21028
rect 12796 19964 12852 20020
rect 13804 20300 13860 20356
rect 13356 19906 13412 19908
rect 13356 19854 13358 19906
rect 13358 19854 13410 19906
rect 13410 19854 13412 19906
rect 13356 19852 13412 19854
rect 13468 19740 13524 19796
rect 14588 20690 14644 20692
rect 14588 20638 14590 20690
rect 14590 20638 14642 20690
rect 14642 20638 14644 20690
rect 14588 20636 14644 20638
rect 14364 20130 14420 20132
rect 14364 20078 14366 20130
rect 14366 20078 14418 20130
rect 14418 20078 14420 20130
rect 14364 20076 14420 20078
rect 14588 20130 14644 20132
rect 14588 20078 14590 20130
rect 14590 20078 14642 20130
rect 14642 20078 14644 20130
rect 14588 20076 14644 20078
rect 16044 23660 16100 23716
rect 16492 23548 16548 23604
rect 16940 23660 16996 23716
rect 16828 22482 16884 22484
rect 16828 22430 16830 22482
rect 16830 22430 16882 22482
rect 16882 22430 16884 22482
rect 16828 22428 16884 22430
rect 16156 21644 16212 21700
rect 16268 22204 16324 22260
rect 16268 21868 16324 21924
rect 16044 20860 16100 20916
rect 16492 21420 16548 21476
rect 15596 20076 15652 20132
rect 15260 19964 15316 20020
rect 12908 19292 12964 19348
rect 13356 19292 13412 19348
rect 12796 19234 12852 19236
rect 12796 19182 12798 19234
rect 12798 19182 12850 19234
rect 12850 19182 12852 19234
rect 12796 19180 12852 19182
rect 12796 16994 12852 16996
rect 12796 16942 12798 16994
rect 12798 16942 12850 16994
rect 12850 16942 12852 16994
rect 12796 16940 12852 16942
rect 14028 19346 14084 19348
rect 14028 19294 14030 19346
rect 14030 19294 14082 19346
rect 14082 19294 14084 19346
rect 14028 19292 14084 19294
rect 15036 19292 15092 19348
rect 13468 19234 13524 19236
rect 13468 19182 13470 19234
rect 13470 19182 13522 19234
rect 13522 19182 13524 19234
rect 13468 19180 13524 19182
rect 14476 18396 14532 18452
rect 16604 20748 16660 20804
rect 17948 25228 18004 25284
rect 18844 26460 18900 26516
rect 23436 28700 23492 28756
rect 20188 27074 20244 27076
rect 20188 27022 20190 27074
rect 20190 27022 20242 27074
rect 20242 27022 20244 27074
rect 20188 27020 20244 27022
rect 20076 26962 20132 26964
rect 20076 26910 20078 26962
rect 20078 26910 20130 26962
rect 20130 26910 20132 26962
rect 20076 26908 20132 26910
rect 20636 27692 20692 27748
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19852 26514 19908 26516
rect 19852 26462 19854 26514
rect 19854 26462 19906 26514
rect 19906 26462 19908 26514
rect 19852 26460 19908 26462
rect 19180 26348 19236 26404
rect 20524 26348 20580 26404
rect 18508 25282 18564 25284
rect 18508 25230 18510 25282
rect 18510 25230 18562 25282
rect 18562 25230 18564 25282
rect 18508 25228 18564 25230
rect 17164 22316 17220 22372
rect 17500 23714 17556 23716
rect 17500 23662 17502 23714
rect 17502 23662 17554 23714
rect 17554 23662 17556 23714
rect 17500 23660 17556 23662
rect 18284 24108 18340 24164
rect 18620 24722 18676 24724
rect 18620 24670 18622 24722
rect 18622 24670 18674 24722
rect 18674 24670 18676 24722
rect 18620 24668 18676 24670
rect 19068 24668 19124 24724
rect 18508 23548 18564 23604
rect 17276 21868 17332 21924
rect 17612 22370 17668 22372
rect 17612 22318 17614 22370
rect 17614 22318 17666 22370
rect 17666 22318 17668 22370
rect 17612 22316 17668 22318
rect 17500 21420 17556 21476
rect 16940 20972 16996 21028
rect 17276 20690 17332 20692
rect 17276 20638 17278 20690
rect 17278 20638 17330 20690
rect 17330 20638 17332 20690
rect 17276 20636 17332 20638
rect 16716 20130 16772 20132
rect 16716 20078 16718 20130
rect 16718 20078 16770 20130
rect 16770 20078 16772 20130
rect 16716 20076 16772 20078
rect 16604 19628 16660 19684
rect 16716 19122 16772 19124
rect 16716 19070 16718 19122
rect 16718 19070 16770 19122
rect 16770 19070 16772 19122
rect 16716 19068 16772 19070
rect 17388 19852 17444 19908
rect 17276 19740 17332 19796
rect 14252 17388 14308 17444
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 15260 18450 15316 18452
rect 15260 18398 15262 18450
rect 15262 18398 15314 18450
rect 15314 18398 15316 18450
rect 15260 18396 15316 18398
rect 16156 18450 16212 18452
rect 16156 18398 16158 18450
rect 16158 18398 16210 18450
rect 16210 18398 16212 18450
rect 16156 18396 16212 18398
rect 16940 18396 16996 18452
rect 16044 18338 16100 18340
rect 16044 18286 16046 18338
rect 16046 18286 16098 18338
rect 16098 18286 16100 18338
rect 16044 18284 16100 18286
rect 15596 17836 15652 17892
rect 14812 17554 14868 17556
rect 14812 17502 14814 17554
rect 14814 17502 14866 17554
rect 14866 17502 14868 17554
rect 14812 17500 14868 17502
rect 15260 17500 15316 17556
rect 14476 16940 14532 16996
rect 14924 16770 14980 16772
rect 14924 16718 14926 16770
rect 14926 16718 14978 16770
rect 14978 16718 14980 16770
rect 14924 16716 14980 16718
rect 15372 16716 15428 16772
rect 16044 17724 16100 17780
rect 18172 22092 18228 22148
rect 18732 22428 18788 22484
rect 18732 22146 18788 22148
rect 18732 22094 18734 22146
rect 18734 22094 18786 22146
rect 18786 22094 18788 22146
rect 18732 22092 18788 22094
rect 19404 26290 19460 26292
rect 19404 26238 19406 26290
rect 19406 26238 19458 26290
rect 19458 26238 19460 26290
rect 19404 26236 19460 26238
rect 20188 26290 20244 26292
rect 20188 26238 20190 26290
rect 20190 26238 20242 26290
rect 20242 26238 20244 26290
rect 20188 26236 20244 26238
rect 21420 27132 21476 27188
rect 20524 25228 20580 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19852 24780 19908 24836
rect 21308 26348 21364 26404
rect 21420 25282 21476 25284
rect 21420 25230 21422 25282
rect 21422 25230 21474 25282
rect 21474 25230 21476 25282
rect 21420 25228 21476 25230
rect 21532 24892 21588 24948
rect 21756 25506 21812 25508
rect 21756 25454 21758 25506
rect 21758 25454 21810 25506
rect 21810 25454 21812 25506
rect 21756 25452 21812 25454
rect 20636 24780 20692 24836
rect 19516 23548 19572 23604
rect 21644 23660 21700 23716
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20972 23266 21028 23268
rect 20972 23214 20974 23266
rect 20974 23214 21026 23266
rect 21026 23214 21028 23266
rect 20972 23212 21028 23214
rect 20860 23154 20916 23156
rect 20860 23102 20862 23154
rect 20862 23102 20914 23154
rect 20914 23102 20916 23154
rect 20860 23100 20916 23102
rect 21196 23154 21252 23156
rect 21196 23102 21198 23154
rect 21198 23102 21250 23154
rect 21250 23102 21252 23154
rect 21196 23100 21252 23102
rect 22876 27132 22932 27188
rect 23436 26908 23492 26964
rect 21980 24668 22036 24724
rect 20300 22988 20356 23044
rect 19516 22370 19572 22372
rect 19516 22318 19518 22370
rect 19518 22318 19570 22370
rect 19570 22318 19572 22370
rect 19516 22316 19572 22318
rect 19516 22092 19572 22148
rect 17948 20636 18004 20692
rect 17612 19292 17668 19348
rect 17724 19068 17780 19124
rect 17500 18396 17556 18452
rect 17948 19628 18004 19684
rect 18844 20914 18900 20916
rect 18844 20862 18846 20914
rect 18846 20862 18898 20914
rect 18898 20862 18900 20914
rect 18844 20860 18900 20862
rect 18284 20748 18340 20804
rect 18732 20802 18788 20804
rect 18732 20750 18734 20802
rect 18734 20750 18786 20802
rect 18786 20750 18788 20802
rect 18732 20748 18788 20750
rect 18620 20076 18676 20132
rect 18620 19628 18676 19684
rect 18956 20076 19012 20132
rect 17948 18284 18004 18340
rect 17724 17778 17780 17780
rect 17724 17726 17726 17778
rect 17726 17726 17778 17778
rect 17778 17726 17780 17778
rect 17724 17724 17780 17726
rect 17164 17612 17220 17668
rect 16716 17442 16772 17444
rect 16716 17390 16718 17442
rect 16718 17390 16770 17442
rect 16770 17390 16772 17442
rect 16716 17388 16772 17390
rect 18844 19346 18900 19348
rect 18844 19294 18846 19346
rect 18846 19294 18898 19346
rect 18898 19294 18900 19346
rect 18844 19292 18900 19294
rect 18956 19852 19012 19908
rect 18284 17724 18340 17780
rect 18508 18508 18564 18564
rect 15596 16716 15652 16772
rect 15484 16156 15540 16212
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 19404 21868 19460 21924
rect 19404 20636 19460 20692
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20188 21980 20244 22036
rect 21868 23212 21924 23268
rect 20300 21868 20356 21924
rect 20412 21532 20468 21588
rect 19740 20690 19796 20692
rect 19740 20638 19742 20690
rect 19742 20638 19794 20690
rect 19794 20638 19796 20690
rect 19740 20636 19796 20638
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19628 20188 19684 20244
rect 19292 19906 19348 19908
rect 19292 19854 19294 19906
rect 19294 19854 19346 19906
rect 19346 19854 19348 19906
rect 19292 19852 19348 19854
rect 19852 19852 19908 19908
rect 19628 19740 19684 19796
rect 20748 22370 20804 22372
rect 20748 22318 20750 22370
rect 20750 22318 20802 22370
rect 20802 22318 20804 22370
rect 20748 22316 20804 22318
rect 20860 20578 20916 20580
rect 20860 20526 20862 20578
rect 20862 20526 20914 20578
rect 20914 20526 20916 20578
rect 20860 20524 20916 20526
rect 20748 19346 20804 19348
rect 20748 19294 20750 19346
rect 20750 19294 20802 19346
rect 20802 19294 20804 19346
rect 20748 19292 20804 19294
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19740 18562 19796 18564
rect 19740 18510 19742 18562
rect 19742 18510 19794 18562
rect 19794 18510 19796 18562
rect 19740 18508 19796 18510
rect 18844 18338 18900 18340
rect 18844 18286 18846 18338
rect 18846 18286 18898 18338
rect 18898 18286 18900 18338
rect 18844 18284 18900 18286
rect 18620 17388 18676 17444
rect 16716 16156 16772 16212
rect 18172 15820 18228 15876
rect 16156 15148 16212 15204
rect 17388 15202 17444 15204
rect 17388 15150 17390 15202
rect 17390 15150 17442 15202
rect 17442 15150 17444 15202
rect 17388 15148 17444 15150
rect 18396 15314 18452 15316
rect 18396 15262 18398 15314
rect 18398 15262 18450 15314
rect 18450 15262 18452 15314
rect 18396 15260 18452 15262
rect 18844 16044 18900 16100
rect 19292 17836 19348 17892
rect 20188 18284 20244 18340
rect 20188 17778 20244 17780
rect 20188 17726 20190 17778
rect 20190 17726 20242 17778
rect 20242 17726 20244 17778
rect 20188 17724 20244 17726
rect 19068 17666 19124 17668
rect 19068 17614 19070 17666
rect 19070 17614 19122 17666
rect 19122 17614 19124 17666
rect 19068 17612 19124 17614
rect 19180 17052 19236 17108
rect 19516 15986 19572 15988
rect 19516 15934 19518 15986
rect 19518 15934 19570 15986
rect 19570 15934 19572 15986
rect 19516 15932 19572 15934
rect 19180 15874 19236 15876
rect 19180 15822 19182 15874
rect 19182 15822 19234 15874
rect 19234 15822 19236 15874
rect 19180 15820 19236 15822
rect 15484 14530 15540 14532
rect 15484 14478 15486 14530
rect 15486 14478 15538 14530
rect 15538 14478 15540 14530
rect 15484 14476 15540 14478
rect 16268 14476 16324 14532
rect 16268 13916 16324 13972
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 17052 14252 17108 14308
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 19404 15484 19460 15540
rect 18956 14306 19012 14308
rect 18956 14254 18958 14306
rect 18958 14254 19010 14306
rect 19010 14254 19012 14306
rect 18956 14252 19012 14254
rect 19180 14252 19236 14308
rect 18508 13970 18564 13972
rect 18508 13918 18510 13970
rect 18510 13918 18562 13970
rect 18562 13918 18564 13970
rect 18508 13916 18564 13918
rect 18956 13916 19012 13972
rect 19516 15260 19572 15316
rect 19404 15148 19460 15204
rect 19852 17388 19908 17444
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20076 17106 20132 17108
rect 20076 17054 20078 17106
rect 20078 17054 20130 17106
rect 20130 17054 20132 17106
rect 20076 17052 20132 17054
rect 20412 18732 20468 18788
rect 20748 18338 20804 18340
rect 20748 18286 20750 18338
rect 20750 18286 20802 18338
rect 20802 18286 20804 18338
rect 20748 18284 20804 18286
rect 20412 17388 20468 17444
rect 20972 20018 21028 20020
rect 20972 19966 20974 20018
rect 20974 19966 21026 20018
rect 21026 19966 21028 20018
rect 20972 19964 21028 19966
rect 20860 17052 20916 17108
rect 21420 22428 21476 22484
rect 21532 21868 21588 21924
rect 21420 20524 21476 20580
rect 21420 19794 21476 19796
rect 21420 19742 21422 19794
rect 21422 19742 21474 19794
rect 21474 19742 21476 19794
rect 21420 19740 21476 19742
rect 21308 17724 21364 17780
rect 21420 18396 21476 18452
rect 21420 17388 21476 17444
rect 23324 25452 23380 25508
rect 22988 25394 23044 25396
rect 22988 25342 22990 25394
rect 22990 25342 23042 25394
rect 23042 25342 23044 25394
rect 22988 25340 23044 25342
rect 22764 25116 22820 25172
rect 23212 24946 23268 24948
rect 23212 24894 23214 24946
rect 23214 24894 23266 24946
rect 23266 24894 23268 24946
rect 23212 24892 23268 24894
rect 22092 23154 22148 23156
rect 22092 23102 22094 23154
rect 22094 23102 22146 23154
rect 22146 23102 22148 23154
rect 22092 23100 22148 23102
rect 21644 20748 21700 20804
rect 21644 20188 21700 20244
rect 22652 23266 22708 23268
rect 22652 23214 22654 23266
rect 22654 23214 22706 23266
rect 22706 23214 22708 23266
rect 22652 23212 22708 23214
rect 23772 26290 23828 26292
rect 23772 26238 23774 26290
rect 23774 26238 23826 26290
rect 23826 26238 23828 26290
rect 23772 26236 23828 26238
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 24780 36706 24836 36708
rect 24780 36654 24782 36706
rect 24782 36654 24834 36706
rect 24834 36654 24836 36706
rect 24780 36652 24836 36654
rect 24220 28754 24276 28756
rect 24220 28702 24222 28754
rect 24222 28702 24274 28754
rect 24274 28702 24276 28754
rect 24220 28700 24276 28702
rect 24108 26012 24164 26068
rect 24668 27132 24724 27188
rect 25676 27132 25732 27188
rect 24556 26514 24612 26516
rect 24556 26462 24558 26514
rect 24558 26462 24610 26514
rect 24610 26462 24612 26514
rect 24556 26460 24612 26462
rect 24444 25340 24500 25396
rect 24556 26236 24612 26292
rect 23884 25116 23940 25172
rect 24108 24108 24164 24164
rect 23436 23884 23492 23940
rect 23772 23938 23828 23940
rect 23772 23886 23774 23938
rect 23774 23886 23826 23938
rect 23826 23886 23828 23938
rect 23772 23884 23828 23886
rect 23548 23826 23604 23828
rect 23548 23774 23550 23826
rect 23550 23774 23602 23826
rect 23602 23774 23604 23826
rect 23548 23772 23604 23774
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 26236 27186 26292 27188
rect 26236 27134 26238 27186
rect 26238 27134 26290 27186
rect 26290 27134 26292 27186
rect 26236 27132 26292 27134
rect 25788 26460 25844 26516
rect 26236 26908 26292 26964
rect 24668 26124 24724 26180
rect 24668 25116 24724 25172
rect 24668 23660 24724 23716
rect 24556 23548 24612 23604
rect 23548 22988 23604 23044
rect 22988 22428 23044 22484
rect 23436 22428 23492 22484
rect 23324 22316 23380 22372
rect 21756 19292 21812 19348
rect 21868 19628 21924 19684
rect 21644 18674 21700 18676
rect 21644 18622 21646 18674
rect 21646 18622 21698 18674
rect 21698 18622 21700 18674
rect 21644 18620 21700 18622
rect 21756 18562 21812 18564
rect 21756 18510 21758 18562
rect 21758 18510 21810 18562
rect 21810 18510 21812 18562
rect 21756 18508 21812 18510
rect 21532 17052 21588 17108
rect 20188 16716 20244 16772
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20636 15932 20692 15988
rect 21196 16828 21252 16884
rect 20860 15538 20916 15540
rect 20860 15486 20862 15538
rect 20862 15486 20914 15538
rect 20914 15486 20916 15538
rect 20860 15484 20916 15486
rect 21644 18284 21700 18340
rect 21644 17666 21700 17668
rect 21644 17614 21646 17666
rect 21646 17614 21698 17666
rect 21698 17614 21700 17666
rect 21644 17612 21700 17614
rect 21644 16828 21700 16884
rect 21980 18620 22036 18676
rect 22092 18508 22148 18564
rect 21980 17836 22036 17892
rect 22092 17500 22148 17556
rect 21980 17164 22036 17220
rect 21644 16658 21700 16660
rect 21644 16606 21646 16658
rect 21646 16606 21698 16658
rect 21698 16606 21700 16658
rect 21644 16604 21700 16606
rect 21532 15986 21588 15988
rect 21532 15934 21534 15986
rect 21534 15934 21586 15986
rect 21586 15934 21588 15986
rect 21532 15932 21588 15934
rect 21644 15538 21700 15540
rect 21644 15486 21646 15538
rect 21646 15486 21698 15538
rect 21698 15486 21700 15538
rect 21644 15484 21700 15486
rect 21196 15426 21252 15428
rect 21196 15374 21198 15426
rect 21198 15374 21250 15426
rect 21250 15374 21252 15426
rect 21196 15372 21252 15374
rect 22428 21980 22484 22036
rect 22988 21586 23044 21588
rect 22988 21534 22990 21586
rect 22990 21534 23042 21586
rect 23042 21534 23044 21586
rect 22988 21532 23044 21534
rect 23548 21810 23604 21812
rect 23548 21758 23550 21810
rect 23550 21758 23602 21810
rect 23602 21758 23604 21810
rect 23548 21756 23604 21758
rect 23660 21868 23716 21924
rect 22652 20636 22708 20692
rect 23772 21586 23828 21588
rect 23772 21534 23774 21586
rect 23774 21534 23826 21586
rect 23826 21534 23828 21586
rect 23772 21532 23828 21534
rect 24556 22092 24612 22148
rect 23996 21756 24052 21812
rect 23884 19852 23940 19908
rect 22876 19628 22932 19684
rect 22540 18450 22596 18452
rect 22540 18398 22542 18450
rect 22542 18398 22594 18450
rect 22594 18398 22596 18450
rect 22540 18396 22596 18398
rect 22428 17666 22484 17668
rect 22428 17614 22430 17666
rect 22430 17614 22482 17666
rect 22482 17614 22484 17666
rect 22428 17612 22484 17614
rect 23548 19628 23604 19684
rect 23772 19516 23828 19572
rect 23548 19180 23604 19236
rect 23324 18450 23380 18452
rect 23324 18398 23326 18450
rect 23326 18398 23378 18450
rect 23378 18398 23380 18450
rect 23324 18396 23380 18398
rect 22204 16604 22260 16660
rect 22204 16098 22260 16100
rect 22204 16046 22206 16098
rect 22206 16046 22258 16098
rect 22258 16046 22260 16098
rect 22204 16044 22260 16046
rect 24220 18620 24276 18676
rect 23884 18284 23940 18340
rect 24556 19516 24612 19572
rect 24668 21532 24724 21588
rect 25676 24780 25732 24836
rect 24892 24162 24948 24164
rect 24892 24110 24894 24162
rect 24894 24110 24946 24162
rect 24946 24110 24948 24162
rect 24892 24108 24948 24110
rect 25116 23938 25172 23940
rect 25116 23886 25118 23938
rect 25118 23886 25170 23938
rect 25170 23886 25172 23938
rect 25116 23884 25172 23886
rect 25452 23826 25508 23828
rect 25452 23774 25454 23826
rect 25454 23774 25506 23826
rect 25506 23774 25508 23826
rect 25452 23772 25508 23774
rect 25340 23714 25396 23716
rect 25340 23662 25342 23714
rect 25342 23662 25394 23714
rect 25394 23662 25396 23714
rect 25340 23660 25396 23662
rect 25564 22146 25620 22148
rect 25564 22094 25566 22146
rect 25566 22094 25618 22146
rect 25618 22094 25620 22146
rect 25564 22092 25620 22094
rect 24892 21980 24948 22036
rect 37660 27074 37716 27076
rect 37660 27022 37662 27074
rect 37662 27022 37714 27074
rect 37714 27022 37716 27074
rect 37660 27020 37716 27022
rect 26908 26908 26964 26964
rect 28476 26908 28532 26964
rect 40012 26908 40068 26964
rect 26348 25116 26404 25172
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 26796 24780 26852 24836
rect 28924 24780 28980 24836
rect 30156 24834 30212 24836
rect 30156 24782 30158 24834
rect 30158 24782 30210 24834
rect 30210 24782 30212 24834
rect 30156 24780 30212 24782
rect 26348 23996 26404 24052
rect 26572 24556 26628 24612
rect 26236 23884 26292 23940
rect 26908 23772 26964 23828
rect 26460 23714 26516 23716
rect 26460 23662 26462 23714
rect 26462 23662 26514 23714
rect 26514 23662 26516 23714
rect 26460 23660 26516 23662
rect 26684 23548 26740 23604
rect 26124 22428 26180 22484
rect 26348 23042 26404 23044
rect 26348 22990 26350 23042
rect 26350 22990 26402 23042
rect 26402 22990 26404 23042
rect 26348 22988 26404 22990
rect 26012 21868 26068 21924
rect 27580 24610 27636 24612
rect 27580 24558 27582 24610
rect 27582 24558 27634 24610
rect 27634 24558 27636 24610
rect 27580 24556 27636 24558
rect 28364 24556 28420 24612
rect 29708 24610 29764 24612
rect 29708 24558 29710 24610
rect 29710 24558 29762 24610
rect 29762 24558 29764 24610
rect 29708 24556 29764 24558
rect 28476 23996 28532 24052
rect 27804 23042 27860 23044
rect 27804 22990 27806 23042
rect 27806 22990 27858 23042
rect 27858 22990 27860 23042
rect 27804 22988 27860 22990
rect 28476 22988 28532 23044
rect 28364 22428 28420 22484
rect 26572 22258 26628 22260
rect 26572 22206 26574 22258
rect 26574 22206 26626 22258
rect 26626 22206 26628 22258
rect 26572 22204 26628 22206
rect 26348 21756 26404 21812
rect 25900 21644 25956 21700
rect 25116 20690 25172 20692
rect 25116 20638 25118 20690
rect 25118 20638 25170 20690
rect 25170 20638 25172 20690
rect 25116 20636 25172 20638
rect 24780 20076 24836 20132
rect 24892 20412 24948 20468
rect 25564 20076 25620 20132
rect 24444 18508 24500 18564
rect 24332 18396 24388 18452
rect 24668 18284 24724 18340
rect 24220 17724 24276 17780
rect 24220 17554 24276 17556
rect 24220 17502 24222 17554
rect 24222 17502 24274 17554
rect 24274 17502 24276 17554
rect 24220 17500 24276 17502
rect 24220 16994 24276 16996
rect 24220 16942 24222 16994
rect 24222 16942 24274 16994
rect 24274 16942 24276 16994
rect 24220 16940 24276 16942
rect 23548 16716 23604 16772
rect 22316 15932 22372 15988
rect 24332 16604 24388 16660
rect 21980 15874 22036 15876
rect 21980 15822 21982 15874
rect 21982 15822 22034 15874
rect 22034 15822 22036 15874
rect 21980 15820 22036 15822
rect 23884 15820 23940 15876
rect 21868 15372 21924 15428
rect 19852 15148 19908 15204
rect 19628 14700 19684 14756
rect 20076 14530 20132 14532
rect 20076 14478 20078 14530
rect 20078 14478 20130 14530
rect 20130 14478 20132 14530
rect 20076 14476 20132 14478
rect 21420 14476 21476 14532
rect 19964 14306 20020 14308
rect 19964 14254 19966 14306
rect 19966 14254 20018 14306
rect 20018 14254 20020 14306
rect 19964 14252 20020 14254
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19852 13916 19908 13972
rect 19852 13580 19908 13636
rect 23884 15260 23940 15316
rect 22204 15036 22260 15092
rect 22204 14754 22260 14756
rect 22204 14702 22206 14754
rect 22206 14702 22258 14754
rect 22258 14702 22260 14754
rect 22204 14700 22260 14702
rect 21980 14530 22036 14532
rect 21980 14478 21982 14530
rect 21982 14478 22034 14530
rect 22034 14478 22036 14530
rect 21980 14476 22036 14478
rect 22540 14530 22596 14532
rect 22540 14478 22542 14530
rect 22542 14478 22594 14530
rect 22594 14478 22596 14530
rect 22540 14476 22596 14478
rect 23436 14476 23492 14532
rect 25452 19852 25508 19908
rect 25340 18562 25396 18564
rect 25340 18510 25342 18562
rect 25342 18510 25394 18562
rect 25394 18510 25396 18562
rect 25340 18508 25396 18510
rect 25564 19234 25620 19236
rect 25564 19182 25566 19234
rect 25566 19182 25618 19234
rect 25618 19182 25620 19234
rect 25564 19180 25620 19182
rect 27244 22092 27300 22148
rect 28140 22146 28196 22148
rect 28140 22094 28142 22146
rect 28142 22094 28194 22146
rect 28194 22094 28196 22146
rect 28140 22092 28196 22094
rect 27132 21644 27188 21700
rect 25900 20972 25956 21028
rect 26908 20690 26964 20692
rect 26908 20638 26910 20690
rect 26910 20638 26962 20690
rect 26962 20638 26964 20690
rect 26908 20636 26964 20638
rect 27020 20578 27076 20580
rect 27020 20526 27022 20578
rect 27022 20526 27074 20578
rect 27074 20526 27076 20578
rect 27020 20524 27076 20526
rect 27916 20748 27972 20804
rect 26236 19122 26292 19124
rect 26236 19070 26238 19122
rect 26238 19070 26290 19122
rect 26290 19070 26292 19122
rect 26236 19068 26292 19070
rect 26460 18732 26516 18788
rect 25788 18450 25844 18452
rect 25788 18398 25790 18450
rect 25790 18398 25842 18450
rect 25842 18398 25844 18450
rect 25788 18396 25844 18398
rect 25900 18338 25956 18340
rect 25900 18286 25902 18338
rect 25902 18286 25954 18338
rect 25954 18286 25956 18338
rect 25900 18284 25956 18286
rect 24892 17164 24948 17220
rect 27020 19234 27076 19236
rect 27020 19182 27022 19234
rect 27022 19182 27074 19234
rect 27074 19182 27076 19234
rect 27020 19180 27076 19182
rect 27692 19122 27748 19124
rect 27692 19070 27694 19122
rect 27694 19070 27746 19122
rect 27746 19070 27748 19122
rect 27692 19068 27748 19070
rect 28028 20524 28084 20580
rect 29260 23324 29316 23380
rect 29036 22876 29092 22932
rect 28812 21810 28868 21812
rect 28812 21758 28814 21810
rect 28814 21758 28866 21810
rect 28866 21758 28868 21810
rect 28812 21756 28868 21758
rect 40012 24892 40068 24948
rect 37660 24556 37716 24612
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 30156 23324 30212 23380
rect 30828 23378 30884 23380
rect 30828 23326 30830 23378
rect 30830 23326 30882 23378
rect 30882 23326 30884 23378
rect 30828 23324 30884 23326
rect 32060 23100 32116 23156
rect 30380 23042 30436 23044
rect 30380 22990 30382 23042
rect 30382 22990 30434 23042
rect 30434 22990 30436 23042
rect 30380 22988 30436 22990
rect 29932 22876 29988 22932
rect 37660 23154 37716 23156
rect 37660 23102 37662 23154
rect 37662 23102 37714 23154
rect 37714 23102 37716 23154
rect 37660 23100 37716 23102
rect 37660 22876 37716 22932
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 32060 22482 32116 22484
rect 32060 22430 32062 22482
rect 32062 22430 32114 22482
rect 32114 22430 32116 22482
rect 32060 22428 32116 22430
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 40012 22204 40068 22260
rect 28588 20748 28644 20804
rect 28924 20524 28980 20580
rect 28476 20412 28532 20468
rect 27132 18620 27188 18676
rect 27244 18562 27300 18564
rect 27244 18510 27246 18562
rect 27246 18510 27298 18562
rect 27298 18510 27300 18562
rect 27244 18508 27300 18510
rect 27356 18396 27412 18452
rect 26796 17778 26852 17780
rect 26796 17726 26798 17778
rect 26798 17726 26850 17778
rect 26850 17726 26852 17778
rect 26796 17724 26852 17726
rect 27804 18450 27860 18452
rect 27804 18398 27806 18450
rect 27806 18398 27858 18450
rect 27858 18398 27860 18450
rect 27804 18396 27860 18398
rect 25340 16604 25396 16660
rect 24780 16044 24836 16100
rect 25564 15314 25620 15316
rect 25564 15262 25566 15314
rect 25566 15262 25618 15314
rect 25618 15262 25620 15314
rect 25564 15260 25620 15262
rect 25340 15090 25396 15092
rect 25340 15038 25342 15090
rect 25342 15038 25394 15090
rect 25394 15038 25396 15090
rect 25340 15036 25396 15038
rect 29148 20412 29204 20468
rect 29036 19964 29092 20020
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 37660 20802 37716 20804
rect 37660 20750 37662 20802
rect 37662 20750 37714 20802
rect 37714 20750 37716 20802
rect 37660 20748 37716 20750
rect 30044 20524 30100 20580
rect 28476 18732 28532 18788
rect 40012 20188 40068 20244
rect 30156 19964 30212 20020
rect 32060 19964 32116 20020
rect 37660 20018 37716 20020
rect 37660 19966 37662 20018
rect 37662 19966 37714 20018
rect 37714 19966 37716 20018
rect 37660 19964 37716 19966
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 40012 19516 40068 19572
rect 28588 18396 28644 18452
rect 27916 17554 27972 17556
rect 27916 17502 27918 17554
rect 27918 17502 27970 17554
rect 27970 17502 27972 17554
rect 27916 17500 27972 17502
rect 26908 15314 26964 15316
rect 26908 15262 26910 15314
rect 26910 15262 26962 15314
rect 26962 15262 26964 15314
rect 26908 15260 26964 15262
rect 28252 15260 28308 15316
rect 24444 14530 24500 14532
rect 24444 14478 24446 14530
rect 24446 14478 24498 14530
rect 24498 14478 24500 14530
rect 24444 14476 24500 14478
rect 22316 13634 22372 13636
rect 22316 13582 22318 13634
rect 22318 13582 22370 13634
rect 22370 13582 22372 13634
rect 22316 13580 22372 13582
rect 22988 13580 23044 13636
rect 23772 13634 23828 13636
rect 23772 13582 23774 13634
rect 23774 13582 23826 13634
rect 23826 13582 23828 13634
rect 23772 13580 23828 13582
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 22316 12962 22372 12964
rect 22316 12910 22318 12962
rect 22318 12910 22370 12962
rect 22370 12910 22372 12962
rect 22316 12908 22372 12910
rect 25004 14306 25060 14308
rect 25004 14254 25006 14306
rect 25006 14254 25058 14306
rect 25058 14254 25060 14306
rect 25004 14252 25060 14254
rect 25340 13916 25396 13972
rect 24892 13132 24948 13188
rect 26012 14252 26068 14308
rect 29820 18508 29876 18564
rect 29820 17612 29876 17668
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 37660 17666 37716 17668
rect 37660 17614 37662 17666
rect 37662 17614 37714 17666
rect 37714 17614 37716 17666
rect 37660 17612 37716 17614
rect 40012 16828 40068 16884
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 37660 15314 37716 15316
rect 37660 15262 37662 15314
rect 37662 15262 37714 15314
rect 37714 15262 37716 15314
rect 37660 15260 37716 15262
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 40012 14812 40068 14868
rect 28588 13970 28644 13972
rect 28588 13918 28590 13970
rect 28590 13918 28642 13970
rect 28642 13918 28644 13970
rect 28588 13916 28644 13918
rect 29260 13916 29316 13972
rect 24332 12684 24388 12740
rect 26236 13186 26292 13188
rect 26236 13134 26238 13186
rect 26238 13134 26290 13186
rect 26290 13134 26292 13186
rect 26236 13132 26292 13134
rect 25228 12908 25284 12964
rect 25228 12684 25284 12740
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 18844 4060 18900 4116
rect 20076 4114 20132 4116
rect 20076 4062 20078 4114
rect 20078 4062 20130 4114
rect 20130 4062 20132 4114
rect 20076 4060 20132 4062
rect 26348 12850 26404 12852
rect 26348 12798 26350 12850
rect 26350 12798 26402 12850
rect 26402 12798 26404 12850
rect 26348 12796 26404 12798
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 28140 12796 28196 12852
rect 25452 12738 25508 12740
rect 25452 12686 25454 12738
rect 25454 12686 25506 12738
rect 25506 12686 25508 12738
rect 25452 12684 25508 12686
rect 25564 4060 25620 4116
rect 24892 3388 24948 3444
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 26796 4114 26852 4116
rect 26796 4062 26798 4114
rect 26798 4062 26850 4114
rect 26850 4062 26852 4114
rect 26796 4060 26852 4062
rect 26124 3388 26180 3444
rect 26236 3612 26292 3668
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 29372 3666 29428 3668
rect 29372 3614 29374 3666
rect 29374 3614 29426 3666
rect 29426 3614 29428 3666
rect 29372 3612 29428 3614
<< metal3 >>
rect 25554 38556 25564 38612
rect 25620 38556 26796 38612
rect 26852 38556 26862 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 22866 38220 22876 38276
rect 22932 38220 25564 38276
rect 25620 38220 25630 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 16818 37436 16828 37492
rect 16884 37436 18396 37492
rect 18452 37436 18462 37492
rect 20178 37436 20188 37492
rect 20244 37436 21420 37492
rect 21476 37436 21486 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 23538 36652 23548 36708
rect 23604 36652 24780 36708
rect 24836 36652 24846 36708
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 23426 28700 23436 28756
rect 23492 28700 24220 28756
rect 24276 28700 24286 28756
rect 0 28308 800 28336
rect 0 28252 4172 28308
rect 4228 28252 4238 28308
rect 0 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 16818 27692 16828 27748
rect 16884 27692 17500 27748
rect 17556 27692 20636 27748
rect 20692 27692 20702 27748
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 16370 27132 16380 27188
rect 16436 27132 17388 27188
rect 17444 27132 17454 27188
rect 21410 27132 21420 27188
rect 21476 27132 22876 27188
rect 22932 27132 24668 27188
rect 24724 27132 25676 27188
rect 25732 27132 26236 27188
rect 26292 27132 26302 27188
rect 13570 27020 13580 27076
rect 13636 27020 16604 27076
rect 16660 27020 16670 27076
rect 18834 27020 18844 27076
rect 18900 27020 20188 27076
rect 20244 27020 20254 27076
rect 31892 27020 37660 27076
rect 37716 27020 37726 27076
rect 31892 26964 31948 27020
rect 41200 26964 42000 26992
rect 17490 26908 17500 26964
rect 17556 26908 20076 26964
rect 20132 26908 20142 26964
rect 23426 26908 23436 26964
rect 23492 26908 26236 26964
rect 26292 26908 26302 26964
rect 26898 26908 26908 26964
rect 26964 26908 28476 26964
rect 28532 26908 31948 26964
rect 40002 26908 40012 26964
rect 40068 26908 42000 26964
rect 41200 26880 42000 26908
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 18834 26460 18844 26516
rect 18900 26460 19852 26516
rect 19908 26460 19918 26516
rect 24546 26460 24556 26516
rect 24612 26460 25788 26516
rect 25844 26460 25854 26516
rect 19170 26348 19180 26404
rect 19236 26348 20524 26404
rect 20580 26348 21308 26404
rect 21364 26348 21374 26404
rect 19394 26236 19404 26292
rect 19460 26236 20188 26292
rect 20244 26236 23772 26292
rect 23828 26236 24556 26292
rect 24612 26236 24622 26292
rect 18050 26124 18060 26180
rect 18116 26124 24668 26180
rect 24724 26124 24734 26180
rect 24108 26068 24164 26124
rect 16594 26012 16604 26068
rect 16660 26012 17500 26068
rect 17556 26012 17566 26068
rect 24098 26012 24108 26068
rect 24164 26012 24174 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 14242 25564 14252 25620
rect 14308 25564 16716 25620
rect 16772 25564 16782 25620
rect 4274 25452 4284 25508
rect 4340 25452 12236 25508
rect 12292 25452 12302 25508
rect 21746 25452 21756 25508
rect 21812 25452 23324 25508
rect 23380 25452 23390 25508
rect 22978 25340 22988 25396
rect 23044 25340 24444 25396
rect 24500 25340 24510 25396
rect 16930 25228 16940 25284
rect 16996 25228 17948 25284
rect 18004 25228 18508 25284
rect 18564 25228 18574 25284
rect 20514 25228 20524 25284
rect 20580 25228 21420 25284
rect 21476 25228 21486 25284
rect 16940 25172 16996 25228
rect 15698 25116 15708 25172
rect 15764 25116 16996 25172
rect 22754 25116 22764 25172
rect 22820 25116 23884 25172
rect 23940 25116 23950 25172
rect 24658 25116 24668 25172
rect 24724 25116 26348 25172
rect 26404 25116 26414 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 0 24948 800 24976
rect 41200 24948 42000 24976
rect 0 24892 1932 24948
rect 1988 24892 1998 24948
rect 21522 24892 21532 24948
rect 21588 24892 23212 24948
rect 23268 24892 23278 24948
rect 40002 24892 40012 24948
rect 40068 24892 42000 24948
rect 0 24864 800 24892
rect 41200 24864 42000 24892
rect 19842 24780 19852 24836
rect 19908 24780 20636 24836
rect 20692 24780 20702 24836
rect 25666 24780 25676 24836
rect 25732 24780 26796 24836
rect 26852 24780 28924 24836
rect 28980 24780 30156 24836
rect 30212 24780 30222 24836
rect 14354 24668 14364 24724
rect 14420 24668 15484 24724
rect 15540 24668 15550 24724
rect 18610 24668 18620 24724
rect 18676 24668 19068 24724
rect 19124 24668 21980 24724
rect 22036 24668 22046 24724
rect 14018 24556 14028 24612
rect 14084 24556 15148 24612
rect 15204 24556 16268 24612
rect 16324 24556 16334 24612
rect 26562 24556 26572 24612
rect 26628 24556 27580 24612
rect 27636 24556 27646 24612
rect 28354 24556 28364 24612
rect 28420 24556 29708 24612
rect 29764 24556 37660 24612
rect 37716 24556 37726 24612
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 18274 24108 18284 24164
rect 18340 24108 24108 24164
rect 24164 24108 24892 24164
rect 24948 24108 24958 24164
rect 13122 23996 13132 24052
rect 13188 23996 14028 24052
rect 14084 23996 14094 24052
rect 14690 23996 14700 24052
rect 14756 23996 15484 24052
rect 15540 23996 26348 24052
rect 26404 23996 28476 24052
rect 28532 23996 28542 24052
rect 4274 23884 4284 23940
rect 4340 23884 9996 23940
rect 10052 23884 10062 23940
rect 12226 23884 12236 23940
rect 12292 23884 15596 23940
rect 15652 23884 15662 23940
rect 23426 23884 23436 23940
rect 23492 23884 23772 23940
rect 23828 23884 25116 23940
rect 25172 23884 26236 23940
rect 26292 23884 26302 23940
rect 12114 23772 12124 23828
rect 12180 23772 13468 23828
rect 13524 23772 13534 23828
rect 23538 23772 23548 23828
rect 23604 23772 25452 23828
rect 25508 23772 26908 23828
rect 26964 23772 26974 23828
rect 16034 23660 16044 23716
rect 16100 23660 16940 23716
rect 16996 23660 17500 23716
rect 17556 23660 17566 23716
rect 21634 23660 21644 23716
rect 21700 23660 24668 23716
rect 24724 23660 24734 23716
rect 25330 23660 25340 23716
rect 25396 23660 26460 23716
rect 26516 23660 26526 23716
rect 0 23604 800 23632
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 9986 23548 9996 23604
rect 10052 23548 14588 23604
rect 14644 23548 14654 23604
rect 16482 23548 16492 23604
rect 16548 23548 18508 23604
rect 18564 23548 19516 23604
rect 19572 23548 19582 23604
rect 24546 23548 24556 23604
rect 24612 23548 26684 23604
rect 26740 23548 26750 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 29250 23324 29260 23380
rect 29316 23324 30156 23380
rect 30212 23324 30828 23380
rect 30884 23324 30894 23380
rect 15026 23212 15036 23268
rect 15092 23212 15708 23268
rect 15764 23212 15774 23268
rect 20962 23212 20972 23268
rect 21028 23212 21868 23268
rect 21924 23212 22652 23268
rect 22708 23212 22718 23268
rect 4274 23100 4284 23156
rect 4340 23100 13580 23156
rect 13636 23100 15820 23156
rect 15876 23100 15886 23156
rect 20850 23100 20860 23156
rect 20916 23100 20926 23156
rect 21186 23100 21196 23156
rect 21252 23100 22092 23156
rect 22148 23100 22158 23156
rect 32050 23100 32060 23156
rect 32116 23100 37660 23156
rect 37716 23100 37726 23156
rect 20860 23044 20916 23100
rect 20290 22988 20300 23044
rect 20356 22988 23548 23044
rect 23604 22988 23614 23044
rect 26338 22988 26348 23044
rect 26404 22988 27804 23044
rect 27860 22988 27870 23044
rect 28466 22988 28476 23044
rect 28532 22988 30380 23044
rect 30436 22988 30446 23044
rect 0 22932 800 22960
rect 41200 22932 42000 22960
rect 0 22876 1932 22932
rect 1988 22876 1998 22932
rect 29026 22876 29036 22932
rect 29092 22876 29932 22932
rect 29988 22876 37660 22932
rect 37716 22876 37726 22932
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 0 22848 800 22876
rect 41200 22848 42000 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 14802 22428 14812 22484
rect 14868 22428 16828 22484
rect 16884 22428 16894 22484
rect 18722 22428 18732 22484
rect 18788 22428 20804 22484
rect 21410 22428 21420 22484
rect 21476 22428 22988 22484
rect 23044 22428 23436 22484
rect 23492 22428 26124 22484
rect 26180 22428 26190 22484
rect 28354 22428 28364 22484
rect 28420 22428 32060 22484
rect 32116 22428 32126 22484
rect 20748 22372 20804 22428
rect 17154 22316 17164 22372
rect 17220 22316 17612 22372
rect 17668 22316 19516 22372
rect 19572 22316 19582 22372
rect 20738 22316 20748 22372
rect 20804 22316 23324 22372
rect 23380 22316 23390 22372
rect 41200 22260 42000 22288
rect 14914 22204 14924 22260
rect 14980 22204 15596 22260
rect 15652 22204 16268 22260
rect 16324 22204 16334 22260
rect 26562 22204 26572 22260
rect 26628 22204 26908 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 26852 22148 26908 22204
rect 41200 22176 42000 22204
rect 18162 22092 18172 22148
rect 18228 22092 18732 22148
rect 18788 22092 18798 22148
rect 19506 22092 19516 22148
rect 19572 22092 20244 22148
rect 24546 22092 24556 22148
rect 24612 22092 25564 22148
rect 25620 22092 25630 22148
rect 26852 22092 27244 22148
rect 27300 22092 28140 22148
rect 28196 22092 28206 22148
rect 20188 22036 20244 22092
rect 15092 21980 19460 22036
rect 20178 21980 20188 22036
rect 20244 21980 22428 22036
rect 22484 21980 24892 22036
rect 24948 21980 24958 22036
rect 15026 21868 15036 21924
rect 15092 21868 15148 21980
rect 19404 21924 19460 21980
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 16258 21868 16268 21924
rect 16324 21868 17276 21924
rect 17332 21868 17342 21924
rect 19394 21868 19404 21924
rect 19460 21868 19470 21924
rect 20290 21868 20300 21924
rect 20356 21868 21532 21924
rect 21588 21868 21598 21924
rect 23650 21868 23660 21924
rect 23716 21868 26012 21924
rect 26068 21868 26078 21924
rect 23538 21756 23548 21812
rect 23604 21756 23996 21812
rect 24052 21756 24062 21812
rect 26338 21756 26348 21812
rect 26404 21756 28812 21812
rect 28868 21756 28878 21812
rect 16146 21644 16156 21700
rect 16212 21644 23828 21700
rect 25890 21644 25900 21700
rect 25956 21644 27132 21700
rect 27188 21644 27198 21700
rect 23772 21588 23828 21644
rect 4274 21532 4284 21588
rect 4340 21532 9996 21588
rect 10052 21532 10062 21588
rect 20402 21532 20412 21588
rect 20468 21532 22988 21588
rect 23044 21532 23054 21588
rect 23762 21532 23772 21588
rect 23828 21532 24668 21588
rect 24724 21532 24734 21588
rect 13794 21420 13804 21476
rect 13860 21420 16492 21476
rect 16548 21420 17500 21476
rect 17556 21420 17566 21476
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 15026 20972 15036 21028
rect 15092 20972 16940 21028
rect 16996 20972 25900 21028
rect 25956 20972 25966 21028
rect 0 20916 800 20944
rect 0 20860 1932 20916
rect 1988 20860 1998 20916
rect 16034 20860 16044 20916
rect 16100 20860 18844 20916
rect 18900 20860 18910 20916
rect 0 20832 800 20860
rect 4274 20748 4284 20804
rect 4340 20748 12572 20804
rect 12628 20748 12638 20804
rect 16594 20748 16604 20804
rect 16660 20748 18284 20804
rect 18340 20748 18732 20804
rect 18788 20748 21644 20804
rect 21700 20748 21710 20804
rect 27906 20748 27916 20804
rect 27972 20748 28588 20804
rect 28644 20748 37660 20804
rect 37716 20748 37726 20804
rect 9986 20636 9996 20692
rect 10052 20636 14588 20692
rect 14644 20636 14654 20692
rect 17266 20636 17276 20692
rect 17332 20636 17948 20692
rect 18004 20636 19404 20692
rect 19460 20636 19740 20692
rect 19796 20636 19806 20692
rect 22642 20636 22652 20692
rect 22708 20636 25116 20692
rect 25172 20636 25182 20692
rect 4162 20524 4172 20580
rect 4228 20524 20860 20580
rect 20916 20524 21420 20580
rect 21476 20524 21486 20580
rect 26852 20468 26908 20692
rect 26964 20636 26974 20692
rect 27010 20524 27020 20580
rect 27076 20524 28028 20580
rect 28084 20524 28924 20580
rect 28980 20524 30044 20580
rect 30100 20524 30110 20580
rect 24882 20412 24892 20468
rect 24948 20412 26908 20468
rect 28466 20412 28476 20468
rect 28532 20412 29148 20468
rect 29204 20412 29214 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 12226 20300 12236 20356
rect 12292 20300 13804 20356
rect 13860 20300 13870 20356
rect 0 20244 800 20272
rect 41200 20244 42000 20272
rect 0 20188 2044 20244
rect 2100 20188 2110 20244
rect 19618 20188 19628 20244
rect 19684 20188 21644 20244
rect 21700 20188 21710 20244
rect 40002 20188 40012 20244
rect 40068 20188 42000 20244
rect 0 20160 800 20188
rect 41200 20160 42000 20188
rect 14354 20076 14364 20132
rect 14420 20076 14430 20132
rect 14578 20076 14588 20132
rect 14644 20076 15596 20132
rect 15652 20076 15662 20132
rect 16706 20076 16716 20132
rect 16772 20076 18620 20132
rect 18676 20076 18686 20132
rect 18946 20076 18956 20132
rect 19012 20076 21028 20132
rect 24770 20076 24780 20132
rect 24836 20076 25564 20132
rect 25620 20076 25630 20132
rect 14364 20020 14420 20076
rect 20972 20020 21028 20076
rect 4274 19964 4284 20020
rect 4340 19964 10108 20020
rect 10164 19964 12796 20020
rect 12852 19964 12862 20020
rect 14364 19964 15260 20020
rect 15316 19964 19684 20020
rect 20962 19964 20972 20020
rect 21028 19964 29036 20020
rect 29092 19964 29102 20020
rect 30146 19964 30156 20020
rect 30212 19964 32060 20020
rect 32116 19964 37660 20020
rect 37716 19964 37726 20020
rect 12114 19852 12124 19908
rect 12180 19852 13356 19908
rect 13412 19852 13422 19908
rect 17378 19852 17388 19908
rect 17444 19852 18956 19908
rect 19012 19852 19292 19908
rect 19348 19852 19358 19908
rect 19628 19796 19684 19964
rect 19842 19852 19852 19908
rect 19908 19852 23884 19908
rect 23940 19852 25452 19908
rect 25508 19852 25518 19908
rect 1922 19740 1932 19796
rect 1988 19740 1998 19796
rect 13458 19740 13468 19796
rect 13524 19740 17276 19796
rect 17332 19740 17342 19796
rect 19618 19740 19628 19796
rect 19684 19740 21420 19796
rect 21476 19740 21486 19796
rect 0 19572 800 19600
rect 1932 19572 1988 19740
rect 16594 19628 16604 19684
rect 16660 19628 17948 19684
rect 18004 19628 18014 19684
rect 18610 19628 18620 19684
rect 18676 19628 21868 19684
rect 21924 19628 22876 19684
rect 22932 19628 23548 19684
rect 23604 19628 23614 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 17948 19572 18004 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 0 19516 1988 19572
rect 17948 19516 23772 19572
rect 23828 19516 24556 19572
rect 24612 19516 24622 19572
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 0 19488 800 19516
rect 41200 19488 42000 19516
rect 12114 19292 12124 19348
rect 12180 19292 12908 19348
rect 12964 19292 13356 19348
rect 13412 19292 14028 19348
rect 14084 19292 15036 19348
rect 15092 19292 15102 19348
rect 17602 19292 17612 19348
rect 17668 19292 18844 19348
rect 18900 19292 18910 19348
rect 20738 19292 20748 19348
rect 20804 19292 21756 19348
rect 21812 19292 21822 19348
rect 12786 19180 12796 19236
rect 12852 19180 13468 19236
rect 13524 19180 13534 19236
rect 23538 19180 23548 19236
rect 23604 19180 25564 19236
rect 25620 19180 27020 19236
rect 27076 19180 27086 19236
rect 16706 19068 16716 19124
rect 16772 19068 17724 19124
rect 17780 19068 17790 19124
rect 26226 19068 26236 19124
rect 26292 19068 27692 19124
rect 27748 19068 27758 19124
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 20402 18732 20412 18788
rect 20468 18732 26460 18788
rect 26516 18732 28476 18788
rect 28532 18732 28542 18788
rect 21634 18620 21644 18676
rect 21700 18620 21980 18676
rect 22036 18620 22046 18676
rect 24210 18620 24220 18676
rect 24276 18620 27132 18676
rect 27188 18620 27198 18676
rect 18498 18508 18508 18564
rect 18564 18508 19740 18564
rect 19796 18508 21756 18564
rect 21812 18508 21822 18564
rect 22082 18508 22092 18564
rect 22148 18508 24444 18564
rect 24500 18508 25340 18564
rect 25396 18508 25406 18564
rect 27234 18508 27244 18564
rect 27300 18508 29820 18564
rect 29876 18508 29886 18564
rect 14466 18396 14476 18452
rect 14532 18396 15260 18452
rect 15316 18396 15326 18452
rect 16146 18396 16156 18452
rect 16212 18396 16940 18452
rect 16996 18396 17500 18452
rect 17556 18396 17566 18452
rect 21410 18396 21420 18452
rect 21476 18396 22540 18452
rect 22596 18396 23324 18452
rect 23380 18396 23390 18452
rect 24322 18396 24332 18452
rect 24388 18396 25788 18452
rect 25844 18396 25854 18452
rect 27346 18396 27356 18452
rect 27412 18396 27804 18452
rect 27860 18396 28588 18452
rect 28644 18396 28654 18452
rect 16034 18284 16044 18340
rect 16100 18284 17948 18340
rect 18004 18284 18014 18340
rect 18834 18284 18844 18340
rect 18900 18284 20188 18340
rect 20244 18284 20254 18340
rect 20738 18284 20748 18340
rect 20804 18284 21644 18340
rect 21700 18284 21710 18340
rect 23874 18284 23884 18340
rect 23940 18284 24668 18340
rect 24724 18284 25900 18340
rect 25956 18284 25966 18340
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 15586 17836 15596 17892
rect 15652 17836 19292 17892
rect 19348 17836 21980 17892
rect 22036 17836 22046 17892
rect 16034 17724 16044 17780
rect 16100 17724 17724 17780
rect 17780 17724 18284 17780
rect 18340 17724 18350 17780
rect 20178 17724 20188 17780
rect 20244 17724 21308 17780
rect 21364 17724 21374 17780
rect 24210 17724 24220 17780
rect 24276 17724 26796 17780
rect 26852 17724 26862 17780
rect 17154 17612 17164 17668
rect 17220 17612 19068 17668
rect 19124 17612 19134 17668
rect 21634 17612 21644 17668
rect 21700 17612 22428 17668
rect 22484 17612 22494 17668
rect 29810 17612 29820 17668
rect 29876 17612 37660 17668
rect 37716 17612 37726 17668
rect 14802 17500 14812 17556
rect 14868 17500 15260 17556
rect 15316 17500 15326 17556
rect 22082 17500 22092 17556
rect 22148 17500 24220 17556
rect 24276 17500 27916 17556
rect 27972 17500 27982 17556
rect 14242 17388 14252 17444
rect 14308 17388 16716 17444
rect 16772 17388 18620 17444
rect 18676 17388 19852 17444
rect 19908 17388 19918 17444
rect 20402 17388 20412 17444
rect 20468 17388 21420 17444
rect 21476 17388 21486 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 21970 17164 21980 17220
rect 22036 17164 24892 17220
rect 24948 17164 24958 17220
rect 19170 17052 19180 17108
rect 19236 17052 20076 17108
rect 20132 17052 20860 17108
rect 20916 17052 20926 17108
rect 21522 17052 21532 17108
rect 21588 17052 24276 17108
rect 24220 16996 24276 17052
rect 12786 16940 12796 16996
rect 12852 16940 14476 16996
rect 14532 16940 14542 16996
rect 24210 16940 24220 16996
rect 24276 16940 24286 16996
rect 41200 16884 42000 16912
rect 21186 16828 21196 16884
rect 21252 16828 21644 16884
rect 21700 16828 21710 16884
rect 40002 16828 40012 16884
rect 40068 16828 42000 16884
rect 41200 16800 42000 16828
rect 14914 16716 14924 16772
rect 14980 16716 15372 16772
rect 15428 16716 15596 16772
rect 15652 16716 15662 16772
rect 20178 16716 20188 16772
rect 20244 16716 23548 16772
rect 23604 16716 23614 16772
rect 21634 16604 21644 16660
rect 21700 16604 22204 16660
rect 22260 16604 22270 16660
rect 24322 16604 24332 16660
rect 24388 16604 25340 16660
rect 25396 16604 25406 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 15474 16156 15484 16212
rect 15540 16156 16716 16212
rect 16772 16156 16782 16212
rect 18834 16044 18844 16100
rect 18900 16044 22204 16100
rect 22260 16044 24780 16100
rect 24836 16044 24846 16100
rect 19506 15932 19516 15988
rect 19572 15932 20636 15988
rect 20692 15932 21532 15988
rect 21588 15932 22316 15988
rect 22372 15932 22382 15988
rect 18162 15820 18172 15876
rect 18228 15820 19180 15876
rect 19236 15820 19246 15876
rect 21970 15820 21980 15876
rect 22036 15820 23884 15876
rect 23940 15820 23950 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 19394 15484 19404 15540
rect 19460 15484 20860 15540
rect 20916 15484 21644 15540
rect 21700 15484 21710 15540
rect 21186 15372 21196 15428
rect 21252 15372 21868 15428
rect 21924 15372 21934 15428
rect 18386 15260 18396 15316
rect 18452 15260 19516 15316
rect 19572 15260 19582 15316
rect 23874 15260 23884 15316
rect 23940 15260 25564 15316
rect 25620 15260 25630 15316
rect 26898 15260 26908 15316
rect 26964 15260 28252 15316
rect 28308 15260 37660 15316
rect 37716 15260 37726 15316
rect 16146 15148 16156 15204
rect 16212 15148 17388 15204
rect 17444 15148 17454 15204
rect 19394 15148 19404 15204
rect 19460 15148 19852 15204
rect 19908 15148 19918 15204
rect 22194 15036 22204 15092
rect 22260 15036 25340 15092
rect 25396 15036 25406 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 41200 14868 42000 14896
rect 40002 14812 40012 14868
rect 40068 14812 42000 14868
rect 41200 14784 42000 14812
rect 19618 14700 19628 14756
rect 19684 14700 22204 14756
rect 22260 14700 22270 14756
rect 15474 14476 15484 14532
rect 15540 14476 16268 14532
rect 16324 14476 16334 14532
rect 20066 14476 20076 14532
rect 20132 14476 21420 14532
rect 21476 14476 21980 14532
rect 22036 14476 22046 14532
rect 22530 14476 22540 14532
rect 22596 14476 23436 14532
rect 23492 14476 24444 14532
rect 24500 14476 24510 14532
rect 17042 14252 17052 14308
rect 17108 14252 18956 14308
rect 19012 14252 19022 14308
rect 19170 14252 19180 14308
rect 19236 14252 19964 14308
rect 20020 14252 20030 14308
rect 24994 14252 25004 14308
rect 25060 14252 26012 14308
rect 26068 14252 26078 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 16258 13916 16268 13972
rect 16324 13916 18508 13972
rect 18564 13916 18956 13972
rect 19012 13916 19852 13972
rect 19908 13916 19918 13972
rect 25330 13916 25340 13972
rect 25396 13916 28588 13972
rect 28644 13916 29260 13972
rect 29316 13916 29326 13972
rect 19842 13580 19852 13636
rect 19908 13580 22316 13636
rect 22372 13580 22382 13636
rect 22978 13580 22988 13636
rect 23044 13580 23772 13636
rect 23828 13580 23838 13636
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 24882 13132 24892 13188
rect 24948 13132 26236 13188
rect 26292 13132 26302 13188
rect 22306 12908 22316 12964
rect 22372 12908 25228 12964
rect 25284 12908 25294 12964
rect 26338 12796 26348 12852
rect 26404 12796 28140 12852
rect 28196 12796 28206 12852
rect 24322 12684 24332 12740
rect 24388 12684 25228 12740
rect 25284 12684 25452 12740
rect 25508 12684 25518 12740
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 18834 4060 18844 4116
rect 18900 4060 20076 4116
rect 20132 4060 20142 4116
rect 25554 4060 25564 4116
rect 25620 4060 26796 4116
rect 26852 4060 26862 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 26226 3612 26236 3668
rect 26292 3612 29372 3668
rect 29428 3612 29438 3668
rect 24882 3388 24892 3444
rect 24948 3388 26124 3444
rect 26180 3388 26190 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _126_
timestamp 1698175906
transform 1 0 22512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _127_
timestamp 1698175906
transform -1 0 26096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _128_
timestamp 1698175906
transform -1 0 24528 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25424 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 26656 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _131_
timestamp 1698175906
transform 1 0 22288 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _132_
timestamp 1698175906
transform 1 0 23184 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _133_
timestamp 1698175906
transform 1 0 26096 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _134_
timestamp 1698175906
transform 1 0 15904 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _135_
timestamp 1698175906
transform -1 0 17248 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _136_
timestamp 1698175906
transform 1 0 15568 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _137_
timestamp 1698175906
transform 1 0 18144 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _138_
timestamp 1698175906
transform 1 0 19488 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _139_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27776 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _140_
timestamp 1698175906
transform -1 0 30576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _141_
timestamp 1698175906
transform -1 0 24080 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _142_
timestamp 1698175906
transform 1 0 22400 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _143_
timestamp 1698175906
transform 1 0 23184 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _144_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26992 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _145_
timestamp 1698175906
transform 1 0 17808 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _146_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23184 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _147_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22400 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _148_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27776 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _149_
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _150_
timestamp 1698175906
transform 1 0 18592 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _151_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _152_
timestamp 1698175906
transform -1 0 22288 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _153_
timestamp 1698175906
transform -1 0 16128 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _154_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14784 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _155_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17920 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _156_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19040 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _157_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16464 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _158_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15008 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _159_
timestamp 1698175906
transform 1 0 15120 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _160_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16912 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _161_
timestamp 1698175906
transform 1 0 16464 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _162_
timestamp 1698175906
transform -1 0 20608 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _163_
timestamp 1698175906
transform 1 0 20272 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _164_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17024 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _165_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14448 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _166_
timestamp 1698175906
transform 1 0 19040 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _167_
timestamp 1698175906
transform -1 0 21392 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _168_
timestamp 1698175906
transform -1 0 18144 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _169_
timestamp 1698175906
transform 1 0 19488 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _170_
timestamp 1698175906
transform -1 0 21952 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _171_
timestamp 1698175906
transform -1 0 20272 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _172_
timestamp 1698175906
transform 1 0 24080 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _173_
timestamp 1698175906
transform -1 0 24528 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _174_
timestamp 1698175906
transform -1 0 17472 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _175_
timestamp 1698175906
transform 1 0 14448 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _176_
timestamp 1698175906
transform -1 0 13888 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _177_
timestamp 1698175906
transform -1 0 17920 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _178_
timestamp 1698175906
transform -1 0 20720 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _179_
timestamp 1698175906
transform -1 0 17808 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _180_
timestamp 1698175906
transform 1 0 19488 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _181_
timestamp 1698175906
transform 1 0 19040 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _182_
timestamp 1698175906
transform -1 0 18592 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _183_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _184_
timestamp 1698175906
transform 1 0 19488 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _185_
timestamp 1698175906
transform 1 0 16464 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _186_
timestamp 1698175906
transform -1 0 19600 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _187_
timestamp 1698175906
transform 1 0 18928 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _188_
timestamp 1698175906
transform 1 0 18704 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _189_
timestamp 1698175906
transform -1 0 15232 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _190_
timestamp 1698175906
transform -1 0 13776 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _191_
timestamp 1698175906
transform 1 0 21504 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _192_
timestamp 1698175906
transform -1 0 25200 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _193_
timestamp 1698175906
transform -1 0 22848 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _194_
timestamp 1698175906
transform -1 0 22288 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _195_
timestamp 1698175906
transform 1 0 26432 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _196_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 25984 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _197_
timestamp 1698175906
transform -1 0 16688 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _198_
timestamp 1698175906
transform 1 0 18592 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _199_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15792 0 1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _200_
timestamp 1698175906
transform 1 0 14560 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _201_
timestamp 1698175906
transform 1 0 26768 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _202_
timestamp 1698175906
transform 1 0 29904 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _203_
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _204_
timestamp 1698175906
transform 1 0 24752 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _205_
timestamp 1698175906
transform -1 0 29344 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _206_
timestamp 1698175906
transform -1 0 24640 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _207_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23968 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _208_
timestamp 1698175906
transform 1 0 25872 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _209_
timestamp 1698175906
transform -1 0 16240 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _210_
timestamp 1698175906
transform -1 0 16016 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _211_
timestamp 1698175906
transform 1 0 26768 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _212_
timestamp 1698175906
transform -1 0 28224 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _213_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 26768 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _214_
timestamp 1698175906
transform -1 0 19712 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _215_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19040 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _216_
timestamp 1698175906
transform -1 0 17696 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _217_
timestamp 1698175906
transform -1 0 26544 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _218_
timestamp 1698175906
transform -1 0 25648 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _219_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21840 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _220_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23856 0 1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _221_
timestamp 1698175906
transform -1 0 24640 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _222_
timestamp 1698175906
transform -1 0 24080 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _223_
timestamp 1698175906
transform -1 0 21952 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _224_
timestamp 1698175906
transform 1 0 26432 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _225_
timestamp 1698175906
transform -1 0 26768 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _226_
timestamp 1698175906
transform -1 0 21504 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _227_
timestamp 1698175906
transform 1 0 22960 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _228_
timestamp 1698175906
transform -1 0 19488 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _229_
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _230_
timestamp 1698175906
transform 1 0 20720 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _231_
timestamp 1698175906
transform 1 0 21952 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _232_
timestamp 1698175906
transform 1 0 22960 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _233_
timestamp 1698175906
transform -1 0 22400 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _234_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24864 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _235_
timestamp 1698175906
transform -1 0 24864 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _236_
timestamp 1698175906
transform 1 0 23408 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _237_
timestamp 1698175906
transform 1 0 23184 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _238_
timestamp 1698175906
transform -1 0 25648 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _239_
timestamp 1698175906
transform -1 0 28672 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _240_
timestamp 1698175906
transform 1 0 26320 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _241_
timestamp 1698175906
transform -1 0 20384 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _242_
timestamp 1698175906
transform 1 0 17248 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _243_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18816 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _244_
timestamp 1698175906
transform 1 0 18368 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _245_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19152 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _246_
timestamp 1698175906
transform 1 0 19264 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _247_
timestamp 1698175906
transform 1 0 19824 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _248_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _249_
timestamp 1698175906
transform 1 0 26768 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _250_
timestamp 1698175906
transform -1 0 13216 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _251_
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _252_
timestamp 1698175906
transform 1 0 11872 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _253_
timestamp 1698175906
transform 1 0 18816 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _254_
timestamp 1698175906
transform -1 0 27776 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _255_
timestamp 1698175906
transform -1 0 13104 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _256_
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _257_
timestamp 1698175906
transform 1 0 16128 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _258_
timestamp 1698175906
transform -1 0 13104 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _259_
timestamp 1698175906
transform 1 0 25200 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _260_
timestamp 1698175906
transform -1 0 16688 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _261_
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _262_
timestamp 1698175906
transform 1 0 26880 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _263_
timestamp 1698175906
transform -1 0 15344 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _264_
timestamp 1698175906
transform 1 0 25536 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _265_
timestamp 1698175906
transform 1 0 15232 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _266_
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _267_
timestamp 1698175906
transform 1 0 22064 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _268_
timestamp 1698175906
transform 1 0 25424 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _269_
timestamp 1698175906
transform 1 0 19712 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _270_
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _271_
timestamp 1698175906
transform 1 0 22736 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _272_
timestamp 1698175906
transform 1 0 26656 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _273_
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _274_
timestamp 1698175906
transform 1 0 16576 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _275_
timestamp 1698175906
transform -1 0 13104 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _276_
timestamp 1698175906
transform 1 0 25312 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _277_
timestamp 1698175906
transform 1 0 22512 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__A2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18032 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__A2
timestamp 1698175906
transform 1 0 19824 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__A1
timestamp 1698175906
transform 1 0 26992 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__A2
timestamp 1698175906
transform 1 0 24080 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__CLK
timestamp 1698175906
transform 1 0 29568 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__CLK
timestamp 1698175906
transform 1 0 30240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__CLK
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__CLK
timestamp 1698175906
transform 1 0 16800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__CLK
timestamp 1698175906
transform 1 0 15232 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__CLK
timestamp 1698175906
transform 1 0 22288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__CLK
timestamp 1698175906
transform 1 0 27776 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__CLK
timestamp 1698175906
transform 1 0 13104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__CLK
timestamp 1698175906
transform 1 0 16576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__CLK
timestamp 1698175906
transform -1 0 19824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__CLK
timestamp 1698175906
transform 1 0 14000 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__CLK
timestamp 1698175906
transform 1 0 29232 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__CLK
timestamp 1698175906
transform 1 0 16688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__CLK
timestamp 1698175906
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__CLK
timestamp 1698175906
transform 1 0 30800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__CLK
timestamp 1698175906
transform 1 0 16240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__CLK
timestamp 1698175906
transform 1 0 30016 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__CLK
timestamp 1698175906
transform 1 0 18480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__CLK
timestamp 1698175906
transform 1 0 28560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__267__CLK
timestamp 1698175906
transform -1 0 25536 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__CLK
timestamp 1698175906
transform 1 0 28896 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__CLK
timestamp 1698175906
transform 1 0 19488 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__270__CLK
timestamp 1698175906
transform 1 0 24640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__271__CLK
timestamp 1698175906
transform 1 0 26208 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__272__CLK
timestamp 1698175906
transform 1 0 30128 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__273__CLK
timestamp 1698175906
transform -1 0 20944 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__274__CLK
timestamp 1698175906
transform 1 0 20608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 22848 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_206
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_210 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24864 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698175906
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_266
timestamp 1698175906
transform 1 0 31136 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_270
timestamp 1698175906
transform 1 0 31584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698175906
transform 1 0 18144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_154
timestamp 1698175906
transform 1 0 18592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_156
timestamp 1698175906
transform 1 0 18816 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_183 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21840 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_199
timestamp 1698175906
transform 1 0 23632 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_216
timestamp 1698175906
transform 1 0 25536 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_243
timestamp 1698175906
transform 1 0 28560 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_275
timestamp 1698175906
transform 1 0 32144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698175906
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_216
timestamp 1698175906
transform 1 0 25536 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_123
timestamp 1698175906
transform 1 0 15120 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_131
timestamp 1698175906
transform 1 0 16016 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_161
timestamp 1698175906
transform 1 0 19376 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_165
timestamp 1698175906
transform 1 0 19824 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698175906
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_220
timestamp 1698175906
transform 1 0 25984 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_225
timestamp 1698175906
transform 1 0 26544 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_150
timestamp 1698175906
transform 1 0 18144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_152
timestamp 1698175906
transform 1 0 18368 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_155
timestamp 1698175906
transform 1 0 18704 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_185
timestamp 1698175906
transform 1 0 22064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_189
timestamp 1698175906
transform 1 0 22512 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_193
timestamp 1698175906
transform 1 0 22960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698175906
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_241
timestamp 1698175906
transform 1 0 28336 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_245
timestamp 1698175906
transform 1 0 28784 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_277
timestamp 1698175906
transform 1 0 32368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698175906
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_153
timestamp 1698175906
transform 1 0 18480 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_163
timestamp 1698175906
transform 1 0 19600 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_169
timestamp 1698175906
transform 1 0 20272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698175906
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_181
timestamp 1698175906
transform 1 0 21616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_191
timestamp 1698175906
transform 1 0 22736 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_199
timestamp 1698175906
transform 1 0 23632 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_212
timestamp 1698175906
transform 1 0 25088 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_242
timestamp 1698175906
transform 1 0 28448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_251
timestamp 1698175906
transform 1 0 29456 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_163
timestamp 1698175906
transform 1 0 19600 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_184
timestamp 1698175906
transform 1 0 21952 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_200
timestamp 1698175906
transform 1 0 23744 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698175906
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_220
timestamp 1698175906
transform 1 0 25984 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_230
timestamp 1698175906
transform 1 0 27104 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_262
timestamp 1698175906
transform 1 0 30688 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698175906
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_314
timestamp 1698175906
transform 1 0 36512 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_322
timestamp 1698175906
transform 1 0 37408 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_136
timestamp 1698175906
transform 1 0 16576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_140
timestamp 1698175906
transform 1 0 17024 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_156
timestamp 1698175906
transform 1 0 18816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_158
timestamp 1698175906
transform 1 0 19040 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_164
timestamp 1698175906
transform 1 0 19712 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698175906
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_187
timestamp 1698175906
transform 1 0 22288 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_219
timestamp 1698175906
transform 1 0 25872 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_235
timestamp 1698175906
transform 1 0 27664 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_88
timestamp 1698175906
transform 1 0 11200 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_92
timestamp 1698175906
transform 1 0 11648 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_135
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_146
timestamp 1698175906
transform 1 0 17696 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_155
timestamp 1698175906
transform 1 0 18704 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_163
timestamp 1698175906
transform 1 0 19600 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_192
timestamp 1698175906
transform 1 0 22848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_194
timestamp 1698175906
transform 1 0 23072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_201
timestamp 1698175906
transform 1 0 23856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698175906
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_220
timestamp 1698175906
transform 1 0 25984 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_224
timestamp 1698175906
transform 1 0 26432 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_226
timestamp 1698175906
transform 1 0 26656 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_256
timestamp 1698175906
transform 1 0 30016 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_260
timestamp 1698175906
transform 1 0 30464 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_115
timestamp 1698175906
transform 1 0 14224 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_122
timestamp 1698175906
transform 1 0 15008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_126
timestamp 1698175906
transform 1 0 15456 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_133
timestamp 1698175906
transform 1 0 16240 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_135
timestamp 1698175906
transform 1 0 16464 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_148
timestamp 1698175906
transform 1 0 17920 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_156
timestamp 1698175906
transform 1 0 18816 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698175906
transform 1 0 20608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_195
timestamp 1698175906
transform 1 0 23184 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_199
timestamp 1698175906
transform 1 0 23632 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_201
timestamp 1698175906
transform 1 0 23856 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_104
timestamp 1698175906
transform 1 0 12992 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_120
timestamp 1698175906
transform 1 0 14784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_122
timestamp 1698175906
transform 1 0 15008 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_128
timestamp 1698175906
transform 1 0 15680 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_134
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698175906
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_194
timestamp 1698175906
transform 1 0 23072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_203
timestamp 1698175906
transform 1 0 24080 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698175906
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_221
timestamp 1698175906
transform 1 0 26096 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_234
timestamp 1698175906
transform 1 0 27552 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_238
timestamp 1698175906
transform 1 0 28000 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_270
timestamp 1698175906
transform 1 0 31584 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 40320 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_69
timestamp 1698175906
transform 1 0 9072 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_85
timestamp 1698175906
transform 1 0 10864 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_93
timestamp 1698175906
transform 1 0 11760 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_97
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_111
timestamp 1698175906
transform 1 0 13776 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_115
timestamp 1698175906
transform 1 0 14224 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_123
timestamp 1698175906
transform 1 0 15120 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_127
timestamp 1698175906
transform 1 0 15568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_129
timestamp 1698175906
transform 1 0 15792 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_139
timestamp 1698175906
transform 1 0 16912 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_195
timestamp 1698175906
transform 1 0 23184 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_213
timestamp 1698175906
transform 1 0 25200 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_227
timestamp 1698175906
transform 1 0 26768 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_231
timestamp 1698175906
transform 1 0 27216 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_240
timestamp 1698175906
transform 1 0 28224 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_242
timestamp 1698175906
transform 1 0 28448 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_276
timestamp 1698175906
transform 1 0 32256 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_308
timestamp 1698175906
transform 1 0 35840 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698175906
transform 1 0 36288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698175906
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 4480 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 8064 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_76
timestamp 1698175906
transform 1 0 9856 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_112
timestamp 1698175906
transform 1 0 13888 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_120
timestamp 1698175906
transform 1 0 14784 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_124
timestamp 1698175906
transform 1 0 15232 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_132
timestamp 1698175906
transform 1 0 16128 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_134
timestamp 1698175906
transform 1 0 16352 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_168
timestamp 1698175906
transform 1 0 20160 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_191
timestamp 1698175906
transform 1 0 22736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_205
timestamp 1698175906
transform 1 0 24304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_262
timestamp 1698175906
transform 1 0 30688 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698175906
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698175906
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 9072 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 9520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 9744 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_126
timestamp 1698175906
transform 1 0 15456 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_134
timestamp 1698175906
transform 1 0 16352 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_171
timestamp 1698175906
transform 1 0 20496 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_233
timestamp 1698175906
transform 1 0 27440 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698175906
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_260
timestamp 1698175906
transform 1 0 30464 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_292
timestamp 1698175906
transform 1 0 34048 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_308
timestamp 1698175906
transform 1 0 35840 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_312
timestamp 1698175906
transform 1 0 36288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698175906
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 4480 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 8064 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_104
timestamp 1698175906
transform 1 0 12992 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_107
timestamp 1698175906
transform 1 0 13328 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_123
timestamp 1698175906
transform 1 0 15120 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_127
timestamp 1698175906
transform 1 0 15568 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_137
timestamp 1698175906
transform 1 0 16688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698175906
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698175906
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_250
timestamp 1698175906
transform 1 0 29344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_254
timestamp 1698175906
transform 1 0 29792 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_258
timestamp 1698175906
transform 1 0 30240 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_274
timestamp 1698175906
transform 1 0 32032 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 40096 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 40320 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_124
timestamp 1698175906
transform 1 0 15232 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_128
timestamp 1698175906
transform 1 0 15680 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_147
timestamp 1698175906
transform 1 0 17808 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_151
timestamp 1698175906
transform 1 0 18256 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_153
timestamp 1698175906
transform 1 0 18480 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_233
timestamp 1698175906
transform 1 0 27440 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_235
timestamp 1698175906
transform 1 0 27664 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_276
timestamp 1698175906
transform 1 0 32256 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_308
timestamp 1698175906
transform 1 0 35840 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_312
timestamp 1698175906
transform 1 0 36288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698175906
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 4480 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_104
timestamp 1698175906
transform 1 0 12992 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698175906
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_148
timestamp 1698175906
transform 1 0 17920 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_164
timestamp 1698175906
transform 1 0 19712 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_172
timestamp 1698175906
transform 1 0 20608 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_216
timestamp 1698175906
transform 1 0 25536 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_218
timestamp 1698175906
transform 1 0 25760 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_261
timestamp 1698175906
transform 1 0 30576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_265
timestamp 1698175906
transform 1 0 31024 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698175906
transform 1 0 31920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_69
timestamp 1698175906
transform 1 0 9072 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_73
timestamp 1698175906
transform 1 0 9520 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_75
timestamp 1698175906
transform 1 0 9744 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_111
timestamp 1698175906
transform 1 0 13776 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_115
timestamp 1698175906
transform 1 0 14224 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_117
timestamp 1698175906
transform 1 0 14448 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_133
timestamp 1698175906
transform 1 0 16240 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_139
timestamp 1698175906
transform 1 0 16912 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_141
timestamp 1698175906
transform 1 0 17136 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_147
timestamp 1698175906
transform 1 0 17808 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_163
timestamp 1698175906
transform 1 0 19600 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698175906
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_193
timestamp 1698175906
transform 1 0 22960 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_205
timestamp 1698175906
transform 1 0 24304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_217
timestamp 1698175906
transform 1 0 25648 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_221
timestamp 1698175906
transform 1 0 26096 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_231
timestamp 1698175906
transform 1 0 27216 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_88
timestamp 1698175906
transform 1 0 11200 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_125
timestamp 1698175906
transform 1 0 15344 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_131
timestamp 1698175906
transform 1 0 16016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_135
timestamp 1698175906
transform 1 0 16464 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_146
timestamp 1698175906
transform 1 0 17696 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_156
timestamp 1698175906
transform 1 0 18816 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_160
timestamp 1698175906
transform 1 0 19264 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_201
timestamp 1698175906
transform 1 0 23856 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698175906
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_255
timestamp 1698175906
transform 1 0 29904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_259
timestamp 1698175906
transform 1 0 30352 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_275
timestamp 1698175906
transform 1 0 32144 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_123
timestamp 1698175906
transform 1 0 15120 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_131
timestamp 1698175906
transform 1 0 16016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_143
timestamp 1698175906
transform 1 0 17360 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_151
timestamp 1698175906
transform 1 0 18256 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_159
timestamp 1698175906
transform 1 0 19152 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_185
timestamp 1698175906
transform 1 0 22064 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_195
timestamp 1698175906
transform 1 0 23184 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_205
timestamp 1698175906
transform 1 0 24304 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_213
timestamp 1698175906
transform 1 0 25200 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_217
timestamp 1698175906
transform 1 0 25648 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_227
timestamp 1698175906
transform 1 0 26768 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698175906
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698175906
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_147
timestamp 1698175906
transform 1 0 17808 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_151
timestamp 1698175906
transform 1 0 18256 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_170
timestamp 1698175906
transform 1 0 20384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_174
timestamp 1698175906
transform 1 0 20832 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_190
timestamp 1698175906
transform 1 0 22624 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_194
timestamp 1698175906
transform 1 0 23072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_204
timestamp 1698175906
transform 1 0 24192 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_214
timestamp 1698175906
transform 1 0 25312 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_244
timestamp 1698175906
transform 1 0 28672 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_248
timestamp 1698175906
transform 1 0 29120 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698175906
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_185
timestamp 1698175906
transform 1 0 22064 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_189
timestamp 1698175906
transform 1 0 22512 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_220
timestamp 1698175906
transform 1 0 25984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_230
timestamp 1698175906
transform 1 0 27104 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698175906
transform 1 0 28000 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_171
timestamp 1698175906
transform 1 0 20496 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_175
timestamp 1698175906
transform 1 0 20944 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_179
timestamp 1698175906
transform 1 0 21392 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_181
timestamp 1698175906
transform 1 0 21616 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_188
timestamp 1698175906
transform 1 0 22400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_192
timestamp 1698175906
transform 1 0 22848 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_199
timestamp 1698175906
transform 1 0 23632 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698175906
transform 1 0 24528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_206
timestamp 1698175906
transform 1 0 24416 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_210
timestamp 1698175906
transform 1 0 24864 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_242
timestamp 1698175906
transform 1 0 28448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698175906
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_193
timestamp 1698175906
transform 1 0 22960 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_197
timestamp 1698175906
transform 1 0 23408 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_225
timestamp 1698175906
transform 1 0 26544 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_168
timestamp 1698175906
transform 1 0 20160 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_195
timestamp 1698175906
transform 1 0 23184 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698175906
transform 1 0 24080 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 25536 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_243
timestamp 1698175906
transform 1 0 28560 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698175906
transform 1 0 32144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24192 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 20272 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 17472 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform -1 0 20384 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 4480 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform -1 0 4480 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 24976 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 25648 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 37520 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform -1 0 4480 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 23632 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 37520 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 18928 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 4480 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 25648 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 37520 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 20160 41200 20272 42000 0 FreeSans 448 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 41200 20160 42000 20272 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 19488 41200 19600 42000 0 FreeSans 448 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 25536 41200 25648 42000 0 FreeSans 448 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 41200 24864 42000 24976 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 22848 41200 22960 42000 0 FreeSans 448 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 23520 41200 23632 42000 0 FreeSans 448 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 41200 14784 42000 14896 0 FreeSans 448 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 16800 41200 16912 42000 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 41200 16800 42000 16912 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 41200 26880 42000 26992 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 30016 22456 30016 22456 0 _000_
rlabel metal2 27720 17024 27720 17024 0 _001_
rlabel metal3 13048 20328 13048 20328 0 _002_
rlabel metal2 14280 16800 14280 16800 0 _003_
rlabel metal2 14504 17192 14504 17192 0 _004_
rlabel metal2 19768 13888 19768 13888 0 _005_
rlabel metal2 24248 17808 24248 17808 0 _006_
rlabel metal3 12768 19880 12768 19880 0 _007_
rlabel metal2 14280 26264 14280 26264 0 _008_
rlabel metal2 17080 13664 17080 13664 0 _009_
rlabel metal3 12824 23800 12824 23800 0 _010_
rlabel metal2 26152 14728 26152 14728 0 _011_
rlabel metal2 15064 23464 15064 23464 0 _012_
rlabel metal2 29960 19600 29960 19600 0 _013_
rlabel metal3 27104 23016 27104 23016 0 _014_
rlabel metal3 14952 24696 14952 24696 0 _015_
rlabel metal2 25816 20328 25816 20328 0 _016_
rlabel metal3 16800 15176 16800 15176 0 _017_
rlabel metal2 26040 14056 26040 14056 0 _018_
rlabel metal2 23016 13328 23016 13328 0 _019_
rlabel metal2 26488 25704 26488 25704 0 _020_
rlabel metal2 20608 24584 20608 24584 0 _021_
rlabel metal2 22120 28280 22120 28280 0 _022_
rlabel metal2 23688 26712 23688 26712 0 _023_
rlabel metal2 26600 24304 26600 24304 0 _024_
rlabel metal2 18312 27720 18312 27720 0 _025_
rlabel metal3 18816 26936 18816 26936 0 _026_
rlabel metal3 20888 23072 20888 23072 0 _027_
rlabel metal3 21056 14504 21056 14504 0 _028_
rlabel metal2 24584 17304 24584 17304 0 _029_
rlabel metal2 15064 20888 15064 20888 0 _030_
rlabel metal2 14952 20356 14952 20356 0 _031_
rlabel metal2 17920 24696 17920 24696 0 _032_
rlabel metal2 17864 26264 17864 26264 0 _033_
rlabel metal2 16632 25760 16632 25760 0 _034_
rlabel metal2 20440 21224 20440 21224 0 _035_
rlabel metal2 15064 22064 15064 22064 0 _036_
rlabel metal2 21784 22624 21784 22624 0 _037_
rlabel metal2 23352 21840 23352 21840 0 _038_
rlabel metal3 18592 22344 18592 22344 0 _039_
rlabel metal2 18928 14504 18928 14504 0 _040_
rlabel metal2 22232 14896 22232 14896 0 _041_
rlabel metal2 14504 23128 14504 23128 0 _042_
rlabel metal2 24920 18200 24920 18200 0 _043_
rlabel metal3 23800 21616 23800 21616 0 _044_
rlabel metal2 19544 15624 19544 15624 0 _045_
rlabel metal3 22960 15848 22960 15848 0 _046_
rlabel metal2 26264 15288 26264 15288 0 _047_
rlabel metal2 16408 22064 16408 22064 0 _048_
rlabel metal3 17472 20888 17472 20888 0 _049_
rlabel metal2 14840 23184 14840 23184 0 _050_
rlabel metal3 27552 20552 27552 20552 0 _051_
rlabel metal2 29848 20888 29848 20888 0 _052_
rlabel metal3 23632 23912 23632 23912 0 _053_
rlabel metal2 26376 22064 26376 22064 0 _054_
rlabel metal3 24528 23800 24528 23800 0 _055_
rlabel metal2 26040 22512 26040 22512 0 _056_
rlabel metal2 15792 24024 15792 24024 0 _057_
rlabel metal2 26600 20272 26600 20272 0 _058_
rlabel metal3 26992 19096 26992 19096 0 _059_
rlabel metal2 18200 15680 18200 15680 0 _060_
rlabel metal2 17528 15456 17528 15456 0 _061_
rlabel metal3 25592 13160 25592 13160 0 _062_
rlabel metal2 23688 14000 23688 14000 0 _063_
rlabel metal2 23464 14112 23464 14112 0 _064_
rlabel metal2 24136 13776 24136 13776 0 _065_
rlabel metal2 24696 23800 24696 23800 0 _066_
rlabel metal2 26712 26152 26712 26152 0 _067_
rlabel metal2 21784 24304 21784 24304 0 _068_
rlabel metal3 22400 24920 22400 24920 0 _069_
rlabel metal2 19152 26264 19152 26264 0 _070_
rlabel metal3 21672 23128 21672 23128 0 _071_
rlabel metal2 22120 22904 22120 22904 0 _072_
rlabel metal2 22736 27832 22736 27832 0 _073_
rlabel metal2 24584 23464 24584 23464 0 _074_
rlabel metal2 24192 26264 24192 26264 0 _075_
rlabel metal2 23632 24024 23632 24024 0 _076_
rlabel metal3 25928 23688 25928 23688 0 _077_
rlabel metal2 27664 23912 27664 23912 0 _078_
rlabel metal3 19376 26488 19376 26488 0 _079_
rlabel metal2 17752 24080 17752 24080 0 _080_
rlabel metal2 18088 24920 18088 24920 0 _081_
rlabel metal2 18816 27048 18816 27048 0 _082_
rlabel metal2 19880 26964 19880 26964 0 _083_
rlabel metal2 20664 18816 20664 18816 0 _084_
rlabel metal3 21840 23240 21840 23240 0 _085_
rlabel metal2 26432 26936 26432 26936 0 _086_
rlabel metal2 24360 18704 24360 18704 0 _087_
rlabel metal2 17976 19824 17976 19824 0 _088_
rlabel metal2 26712 15064 26712 15064 0 _089_
rlabel metal2 14616 22120 14616 22120 0 _090_
rlabel metal2 18648 20048 18648 20048 0 _091_
rlabel metal2 21448 22344 21448 22344 0 _092_
rlabel metal2 26600 22680 26600 22680 0 _093_
rlabel metal3 16856 18424 16856 18424 0 _094_
rlabel metal2 18200 21504 18200 21504 0 _095_
rlabel metal2 21336 17808 21336 17808 0 _096_
rlabel metal2 26488 18984 26488 18984 0 _097_
rlabel metal2 28504 22736 28504 22736 0 _098_
rlabel metal2 21448 17528 21448 17528 0 _099_
rlabel metal2 22288 19992 22288 19992 0 _100_
rlabel metal2 24528 13832 24528 13832 0 _101_
rlabel metal2 28168 17808 28168 17808 0 _102_
rlabel metal2 21784 17640 21784 17640 0 _103_
rlabel metal2 22064 18984 22064 18984 0 _104_
rlabel metal2 21672 19432 21672 19432 0 _105_
rlabel metal2 13944 20468 13944 20468 0 _106_
rlabel metal2 22456 21000 22456 21000 0 _107_
rlabel metal3 14392 20048 14392 20048 0 _108_
rlabel metal2 19320 18144 19320 18144 0 _109_
rlabel metal2 14840 22176 14840 22176 0 _110_
rlabel metal2 14280 20832 14280 20832 0 _111_
rlabel metal2 18984 19544 18984 19544 0 _112_
rlabel metal2 17752 21448 17752 21448 0 _113_
rlabel metal2 15288 17248 15288 17248 0 _114_
rlabel metal2 15624 18928 15624 18928 0 _115_
rlabel metal2 13832 21224 13832 21224 0 _116_
rlabel metal2 17192 18312 17192 18312 0 _117_
rlabel metal2 20552 21448 20552 21448 0 _118_
rlabel metal2 18984 20328 18984 20328 0 _119_
rlabel metal2 13496 20272 13496 20272 0 _120_
rlabel metal3 19600 14280 19600 14280 0 _121_
rlabel metal2 20888 16184 20888 16184 0 _122_
rlabel metal2 17976 20608 17976 20608 0 _123_
rlabel metal3 2478 28280 2478 28280 0 clk
rlabel metal2 25200 20664 25200 20664 0 clknet_0_clk
rlabel metal2 20776 27720 20776 27720 0 clknet_1_0__leaf_clk
rlabel metal2 22904 27104 22904 27104 0 clknet_1_1__leaf_clk
rlabel metal2 17976 17752 17976 17752 0 dut22.count\[0\]
rlabel metal2 15400 16800 15400 16800 0 dut22.count\[1\]
rlabel metal2 21672 17976 21672 17976 0 dut22.count\[2\]
rlabel metal2 24696 18032 24696 18032 0 dut22.count\[3\]
rlabel metal2 23800 24808 23800 24808 0 net1
rlabel metal2 25144 12880 25144 12880 0 net10
rlabel metal2 29960 22960 29960 22960 0 net11
rlabel metal2 12264 25032 12264 25032 0 net12
rlabel metal2 25816 32200 25816 32200 0 net13
rlabel metal3 33712 24584 33712 24584 0 net14
rlabel metal2 13608 23072 13608 23072 0 net15
rlabel metal2 24528 31920 24528 31920 0 net16
rlabel metal2 23464 28280 23464 28280 0 net17
rlabel metal3 32984 15288 32984 15288 0 net18
rlabel metal2 10024 23800 10024 23800 0 net19
rlabel metal2 20328 29820 20328 29820 0 net2
rlabel metal2 19152 13048 19152 13048 0 net20
rlabel metal3 16912 27160 16912 27160 0 net21
rlabel metal2 10024 20776 10024 20776 0 net22
rlabel metal2 25816 8512 25816 8512 0 net23
rlabel metal2 29848 17192 29848 17192 0 net24
rlabel metal2 26936 26992 26936 26992 0 net25
rlabel metal2 32088 22792 32088 22792 0 net26
rlabel metal2 28616 21112 28616 21112 0 net3
rlabel metal2 17640 5964 17640 5964 0 net4
rlabel metal2 19600 27160 19600 27160 0 net5
rlabel metal3 8456 20776 8456 20776 0 net6
rlabel metal2 28168 12712 28168 12712 0 net7
rlabel metal2 32088 19656 32088 19656 0 net8
rlabel metal2 10136 19936 10136 19936 0 net9
rlabel metal2 22232 39690 22232 39690 0 segm[0]
rlabel metal2 20216 39354 20216 39354 0 segm[10]
rlabel metal2 40040 20552 40040 20552 0 segm[11]
rlabel metal2 18200 2198 18200 2198 0 segm[12]
rlabel metal2 19544 39746 19544 39746 0 segm[13]
rlabel metal3 1414 20216 1414 20216 0 segm[1]
rlabel metal2 26264 2198 26264 2198 0 segm[2]
rlabel metal2 40040 19656 40040 19656 0 segm[3]
rlabel metal3 1358 19544 1358 19544 0 segm[4]
rlabel metal2 24920 2086 24920 2086 0 segm[5]
rlabel metal2 40040 22344 40040 22344 0 segm[6]
rlabel metal3 1358 24920 1358 24920 0 segm[7]
rlabel metal2 25592 39914 25592 39914 0 segm[8]
rlabel metal2 40040 25256 40040 25256 0 segm[9]
rlabel metal3 1358 22904 1358 22904 0 sel[0]
rlabel metal2 22904 39746 22904 39746 0 sel[10]
rlabel metal2 23576 38962 23576 38962 0 sel[11]
rlabel metal2 40040 15008 40040 15008 0 sel[1]
rlabel metal3 1358 23576 1358 23576 0 sel[2]
rlabel metal2 18872 2422 18872 2422 0 sel[3]
rlabel metal2 16856 39354 16856 39354 0 sel[4]
rlabel metal3 1358 20888 1358 20888 0 sel[5]
rlabel metal2 25592 2422 25592 2422 0 sel[6]
rlabel metal2 40040 17304 40040 17304 0 sel[7]
rlabel metal2 40040 27048 40040 27048 0 sel[8]
rlabel metal3 40642 22904 40642 22904 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
